module NV_NVDLA_CMAC_CORE_active(nvdla_core_clk, nvdla_core_rstn, cfg_is_fp16, cfg_is_int16, cfg_is_int8, cfg_reg_en, in_dat_data0, in_dat_data1, in_dat_data10, in_dat_data100, in_dat_data101, in_dat_data102, in_dat_data103, in_dat_data104, in_dat_data105, in_dat_data106, in_dat_data107, in_dat_data108, in_dat_data109, in_dat_data11, in_dat_data110, in_dat_data111, in_dat_data112, in_dat_data113, in_dat_data114, in_dat_data115, in_dat_data116, in_dat_data117, in_dat_data118, in_dat_data119, in_dat_data12, in_dat_data120, in_dat_data121, in_dat_data122, in_dat_data123, in_dat_data124, in_dat_data125, in_dat_data126, in_dat_data127, in_dat_data13, in_dat_data14, in_dat_data15, in_dat_data16, in_dat_data17, in_dat_data18, in_dat_data19, in_dat_data2, in_dat_data20, in_dat_data21, in_dat_data22, in_dat_data23, in_dat_data24, in_dat_data25, in_dat_data26, in_dat_data27, in_dat_data28, in_dat_data29, in_dat_data3, in_dat_data30, in_dat_data31, in_dat_data32, in_dat_data33, in_dat_data34, in_dat_data35, in_dat_data36, in_dat_data37, in_dat_data38, in_dat_data39, in_dat_data4, in_dat_data40, in_dat_data41, in_dat_data42, in_dat_data43, in_dat_data44, in_dat_data45, in_dat_data46, in_dat_data47, in_dat_data48, in_dat_data49, in_dat_data5, in_dat_data50, in_dat_data51, in_dat_data52, in_dat_data53, in_dat_data54, in_dat_data55, in_dat_data56, in_dat_data57, in_dat_data58, in_dat_data59, in_dat_data6, in_dat_data60, in_dat_data61, in_dat_data62, in_dat_data63, in_dat_data64, in_dat_data65, in_dat_data66, in_dat_data67, in_dat_data68, in_dat_data69, in_dat_data7, in_dat_data70, in_dat_data71, in_dat_data72, in_dat_data73, in_dat_data74, in_dat_data75, in_dat_data76, in_dat_data77, in_dat_data78, in_dat_data79, in_dat_data8, in_dat_data80, in_dat_data81, in_dat_data82, in_dat_data83, in_dat_data84, in_dat_data85, in_dat_data86, in_dat_data87, in_dat_data88, in_dat_data89, in_dat_data9, in_dat_data90, in_dat_data91, in_dat_data92, in_dat_data93, in_dat_data94, in_dat_data95, in_dat_data96, in_dat_data97, in_dat_data98, in_dat_data99, in_dat_mask, in_dat_pvld, in_dat_stripe_end, in_dat_stripe_st, in_wt_data0, in_wt_data1, in_wt_data10, in_wt_data100, in_wt_data101, in_wt_data102, in_wt_data103, in_wt_data104, in_wt_data105, in_wt_data106, in_wt_data107, in_wt_data108, in_wt_data109, in_wt_data11, in_wt_data110, in_wt_data111, in_wt_data112, in_wt_data113, in_wt_data114, in_wt_data115, in_wt_data116, in_wt_data117, in_wt_data118, in_wt_data119, in_wt_data12, in_wt_data120, in_wt_data121, in_wt_data122, in_wt_data123, in_wt_data124, in_wt_data125, in_wt_data126, in_wt_data127, in_wt_data13, in_wt_data14, in_wt_data15, in_wt_data16, in_wt_data17, in_wt_data18, in_wt_data19, in_wt_data2, in_wt_data20, in_wt_data21, in_wt_data22, in_wt_data23, in_wt_data24, in_wt_data25, in_wt_data26, in_wt_data27, in_wt_data28, in_wt_data29, in_wt_data3, in_wt_data30, in_wt_data31, in_wt_data32, in_wt_data33, in_wt_data34, in_wt_data35, in_wt_data36, in_wt_data37, in_wt_data38, in_wt_data39, in_wt_data4, in_wt_data40, in_wt_data41, in_wt_data42, in_wt_data43, in_wt_data44, in_wt_data45, in_wt_data46, in_wt_data47, in_wt_data48, in_wt_data49, in_wt_data5, in_wt_data50, in_wt_data51, in_wt_data52, in_wt_data53, in_wt_data54, in_wt_data55, in_wt_data56, in_wt_data57, in_wt_data58, in_wt_data59, in_wt_data6, in_wt_data60, in_wt_data61, in_wt_data62, in_wt_data63, in_wt_data64, in_wt_data65, in_wt_data66, in_wt_data67, in_wt_data68, in_wt_data69, in_wt_data7, in_wt_data70, in_wt_data71, in_wt_data72, in_wt_data73, in_wt_data74, in_wt_data75, in_wt_data76, in_wt_data77, in_wt_data78, in_wt_data79, in_wt_data8, in_wt_data80, in_wt_data81, in_wt_data82, in_wt_data83, in_wt_data84, in_wt_data85, in_wt_data86, in_wt_data87, in_wt_data88, in_wt_data89, in_wt_data9, in_wt_data90, in_wt_data91, in_wt_data92, in_wt_data93, in_wt_data94, in_wt_data95, in_wt_data96, in_wt_data97, in_wt_data98, in_wt_data99, in_wt_mask, in_wt_pvld, in_wt_sel, dat0_actv_data, dat0_actv_nan, dat0_actv_nz, dat0_actv_pvld, dat0_pre_exp, dat0_pre_mask, dat0_pre_pvld, dat0_pre_stripe_end, dat0_pre_stripe_st, dat1_actv_data, dat1_actv_nan, dat1_actv_nz, dat1_actv_pvld, dat1_pre_exp, dat1_pre_mask, dat1_pre_pvld, dat1_pre_stripe_end, dat1_pre_stripe_st, dat2_actv_data, dat2_actv_nan, dat2_actv_nz, dat2_actv_pvld, dat2_pre_exp, dat2_pre_mask, dat2_pre_pvld, dat2_pre_stripe_end, dat2_pre_stripe_st, dat3_actv_data, dat3_actv_nan, dat3_actv_nz, dat3_actv_pvld, dat3_pre_exp, dat3_pre_mask, dat3_pre_pvld, dat3_pre_stripe_end, dat3_pre_stripe_st, dat4_actv_data, dat4_actv_nan, dat4_actv_nz, dat4_actv_pvld, dat4_pre_exp, dat4_pre_mask, dat4_pre_pvld, dat4_pre_stripe_end, dat4_pre_stripe_st, dat5_actv_data, dat5_actv_nan, dat5_actv_nz, dat5_actv_pvld, dat5_pre_exp, dat5_pre_mask, dat5_pre_pvld, dat5_pre_stripe_end, dat5_pre_stripe_st, dat6_actv_data, dat6_actv_nan, dat6_actv_nz, dat6_actv_pvld, dat6_pre_exp, dat6_pre_mask, dat6_pre_pvld, dat6_pre_stripe_end, dat6_pre_stripe_st, dat7_actv_data, dat7_actv_nan, dat7_actv_nz, dat7_actv_pvld, dat7_pre_exp, dat7_pre_mask, dat7_pre_pvld, dat7_pre_stripe_end, dat7_pre_stripe_st, wt0_actv_data, wt0_actv_nan, wt0_actv_nz, wt0_actv_pvld, wt0_sd_exp, wt0_sd_mask, wt0_sd_pvld, wt1_actv_data, wt1_actv_nan, wt1_actv_nz, wt1_actv_pvld, wt1_sd_exp, wt1_sd_mask, wt1_sd_pvld, wt2_actv_data, wt2_actv_nan, wt2_actv_nz, wt2_actv_pvld, wt2_sd_exp, wt2_sd_mask, wt2_sd_pvld, wt3_actv_data, wt3_actv_nan, wt3_actv_nz, wt3_actv_pvld, wt3_sd_exp, wt3_sd_mask, wt3_sd_pvld, wt4_actv_data, wt4_actv_nan, wt4_actv_nz, wt4_actv_pvld, wt4_sd_exp, wt4_sd_mask, wt4_sd_pvld, wt5_actv_data, wt5_actv_nan, wt5_actv_nz, wt5_actv_pvld, wt5_sd_exp, wt5_sd_mask, wt5_sd_pvld, wt6_actv_data, wt6_actv_nan, wt6_actv_nz, wt6_actv_pvld, wt6_sd_exp, wt6_sd_mask, wt6_sd_pvld, wt7_actv_data, wt7_actv_nan, wt7_actv_nz, wt7_actv_pvld, wt7_sd_exp, wt7_sd_mask, wt7_sd_pvld);
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1783" *)
  wire [97:0] _00000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1844" *)
  wire [63:0] _00001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1722" *)
  wire [64:0] _00002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31923" *)
  wire [7:0] _00003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31933" *)
  wire [7:0] _00004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31943" *)
  wire [7:0] _00005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30793" *)
  wire [7:0] _00006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30803" *)
  wire [7:0] _00007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30813" *)
  wire [7:0] _00008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30823" *)
  wire [7:0] _00009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30833" *)
  wire [7:0] _00010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30843" *)
  wire [7:0] _00011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30853" *)
  wire [7:0] _00012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30863" *)
  wire [7:0] _00013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30683" *)
  wire [7:0] _00014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30873" *)
  wire [7:0] _00015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30883" *)
  wire [7:0] _00016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30893" *)
  wire [7:0] _00017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30903" *)
  wire [7:0] _00018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30913" *)
  wire [7:0] _00019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30923" *)
  wire [7:0] _00020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30933" *)
  wire [7:0] _00021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30943" *)
  wire [7:0] _00022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30953" *)
  wire [7:0] _00023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30963" *)
  wire [7:0] _00024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30693" *)
  wire [7:0] _00025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30973" *)
  wire [7:0] _00026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30983" *)
  wire [7:0] _00027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30993" *)
  wire [7:0] _00028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31003" *)
  wire [7:0] _00029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31013" *)
  wire [7:0] _00030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31023" *)
  wire [7:0] _00031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31033" *)
  wire [7:0] _00032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31043" *)
  wire [7:0] _00033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31053" *)
  wire [7:0] _00034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31063" *)
  wire [7:0] _00035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30703" *)
  wire [7:0] _00036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31073" *)
  wire [7:0] _00037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31083" *)
  wire [7:0] _00038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31093" *)
  wire [7:0] _00039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31103" *)
  wire [7:0] _00040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31113" *)
  wire [7:0] _00041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31123" *)
  wire [7:0] _00042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31133" *)
  wire [7:0] _00043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31143" *)
  wire [7:0] _00044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31153" *)
  wire [7:0] _00045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31163" *)
  wire [7:0] _00046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30713" *)
  wire [7:0] _00047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31173" *)
  wire [7:0] _00048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31183" *)
  wire [7:0] _00049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31193" *)
  wire [7:0] _00050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31203" *)
  wire [7:0] _00051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31213" *)
  wire [7:0] _00052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31223" *)
  wire [7:0] _00053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31233" *)
  wire [7:0] _00054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31243" *)
  wire [7:0] _00055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31253" *)
  wire [7:0] _00056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31263" *)
  wire [7:0] _00057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30723" *)
  wire [7:0] _00058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31273" *)
  wire [7:0] _00059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31283" *)
  wire [7:0] _00060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31293" *)
  wire [7:0] _00061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31303" *)
  wire [7:0] _00062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31313" *)
  wire [7:0] _00063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31323" *)
  wire [7:0] _00064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31333" *)
  wire [7:0] _00065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31343" *)
  wire [7:0] _00066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31353" *)
  wire [7:0] _00067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31363" *)
  wire [7:0] _00068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30733" *)
  wire [7:0] _00069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31373" *)
  wire [7:0] _00070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31383" *)
  wire [7:0] _00071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31393" *)
  wire [7:0] _00072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31403" *)
  wire [7:0] _00073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31413" *)
  wire [7:0] _00074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31423" *)
  wire [7:0] _00075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31433" *)
  wire [7:0] _00076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31443" *)
  wire [7:0] _00077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31453" *)
  wire [7:0] _00078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31463" *)
  wire [7:0] _00079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30743" *)
  wire [7:0] _00080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31473" *)
  wire [7:0] _00081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31483" *)
  wire [7:0] _00082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31493" *)
  wire [7:0] _00083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31503" *)
  wire [7:0] _00084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31513" *)
  wire [7:0] _00085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31523" *)
  wire [7:0] _00086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31533" *)
  wire [7:0] _00087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31543" *)
  wire [7:0] _00088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31553" *)
  wire [7:0] _00089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31563" *)
  wire [7:0] _00090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30753" *)
  wire [7:0] _00091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31573" *)
  wire [7:0] _00092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31583" *)
  wire [7:0] _00093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31593" *)
  wire [7:0] _00094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31603" *)
  wire [7:0] _00095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31613" *)
  wire [7:0] _00096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31623" *)
  wire [7:0] _00097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31633" *)
  wire [7:0] _00098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31643" *)
  wire [7:0] _00099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31653" *)
  wire [7:0] _00100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31663" *)
  wire [7:0] _00101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30763" *)
  wire [7:0] _00102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30673" *)
  wire [7:0] _00103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31673" *)
  wire [7:0] _00104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31683" *)
  wire [7:0] _00105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31693" *)
  wire [7:0] _00106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31703" *)
  wire [7:0] _00107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31713" *)
  wire [7:0] _00108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31723" *)
  wire [7:0] _00109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31733" *)
  wire [7:0] _00110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31743" *)
  wire [7:0] _00111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31753" *)
  wire [7:0] _00112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31763" *)
  wire [7:0] _00113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30773" *)
  wire [7:0] _00114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31773" *)
  wire [7:0] _00115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31783" *)
  wire [7:0] _00116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31793" *)
  wire [7:0] _00117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31803" *)
  wire [7:0] _00118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31813" *)
  wire [7:0] _00119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31823" *)
  wire [7:0] _00120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31833" *)
  wire [7:0] _00121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31843" *)
  wire [7:0] _00122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31853" *)
  wire [7:0] _00123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31863" *)
  wire [7:0] _00124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30783" *)
  wire [7:0] _00125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31873" *)
  wire [7:0] _00126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31883" *)
  wire [7:0] _00127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31893" *)
  wire [7:0] _00128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31903" *)
  wire [7:0] _00129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31913" *)
  wire [7:0] _00130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33230" *)
  wire [7:0] _00131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33240" *)
  wire [7:0] _00132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33250" *)
  wire [7:0] _00133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32100" *)
  wire [7:0] _00134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32110" *)
  wire [7:0] _00135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32120" *)
  wire [7:0] _00136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32130" *)
  wire [7:0] _00137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32140" *)
  wire [7:0] _00138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32150" *)
  wire [7:0] _00139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32160" *)
  wire [7:0] _00140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32170" *)
  wire [7:0] _00141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31990" *)
  wire [7:0] _00142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32180" *)
  wire [7:0] _00143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32190" *)
  wire [7:0] _00144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32200" *)
  wire [7:0] _00145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32210" *)
  wire [7:0] _00146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32220" *)
  wire [7:0] _00147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32230" *)
  wire [7:0] _00148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32240" *)
  wire [7:0] _00149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32250" *)
  wire [7:0] _00150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32260" *)
  wire [7:0] _00151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32270" *)
  wire [7:0] _00152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32000" *)
  wire [7:0] _00153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32280" *)
  wire [7:0] _00154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32290" *)
  wire [7:0] _00155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32300" *)
  wire [7:0] _00156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32310" *)
  wire [7:0] _00157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32320" *)
  wire [7:0] _00158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32330" *)
  wire [7:0] _00159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32340" *)
  wire [7:0] _00160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32350" *)
  wire [7:0] _00161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32360" *)
  wire [7:0] _00162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32370" *)
  wire [7:0] _00163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32010" *)
  wire [7:0] _00164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32380" *)
  wire [7:0] _00165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32390" *)
  wire [7:0] _00166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32400" *)
  wire [7:0] _00167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32410" *)
  wire [7:0] _00168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32420" *)
  wire [7:0] _00169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32430" *)
  wire [7:0] _00170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32440" *)
  wire [7:0] _00171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32450" *)
  wire [7:0] _00172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32460" *)
  wire [7:0] _00173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32470" *)
  wire [7:0] _00174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32020" *)
  wire [7:0] _00175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32480" *)
  wire [7:0] _00176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32490" *)
  wire [7:0] _00177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32500" *)
  wire [7:0] _00178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32510" *)
  wire [7:0] _00179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32520" *)
  wire [7:0] _00180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32530" *)
  wire [7:0] _00181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32540" *)
  wire [7:0] _00182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32550" *)
  wire [7:0] _00183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32560" *)
  wire [7:0] _00184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32570" *)
  wire [7:0] _00185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32030" *)
  wire [7:0] _00186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32580" *)
  wire [7:0] _00187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32590" *)
  wire [7:0] _00188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32600" *)
  wire [7:0] _00189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32610" *)
  wire [7:0] _00190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32620" *)
  wire [7:0] _00191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32630" *)
  wire [7:0] _00192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32640" *)
  wire [7:0] _00193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32650" *)
  wire [7:0] _00194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32660" *)
  wire [7:0] _00195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32670" *)
  wire [7:0] _00196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32040" *)
  wire [7:0] _00197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32680" *)
  wire [7:0] _00198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32690" *)
  wire [7:0] _00199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32700" *)
  wire [7:0] _00200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32710" *)
  wire [7:0] _00201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32720" *)
  wire [7:0] _00202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32730" *)
  wire [7:0] _00203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32740" *)
  wire [7:0] _00204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32750" *)
  wire [7:0] _00205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32760" *)
  wire [7:0] _00206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32770" *)
  wire [7:0] _00207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32050" *)
  wire [7:0] _00208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32780" *)
  wire [7:0] _00209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32790" *)
  wire [7:0] _00210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32800" *)
  wire [7:0] _00211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32810" *)
  wire [7:0] _00212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32820" *)
  wire [7:0] _00213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32830" *)
  wire [7:0] _00214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32840" *)
  wire [7:0] _00215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32850" *)
  wire [7:0] _00216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32860" *)
  wire [7:0] _00217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32870" *)
  wire [7:0] _00218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32060" *)
  wire [7:0] _00219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32880" *)
  wire [7:0] _00220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32890" *)
  wire [7:0] _00221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32900" *)
  wire [7:0] _00222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32910" *)
  wire [7:0] _00223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32920" *)
  wire [7:0] _00224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32930" *)
  wire [7:0] _00225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32940" *)
  wire [7:0] _00226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32950" *)
  wire [7:0] _00227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32960" *)
  wire [7:0] _00228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32970" *)
  wire [7:0] _00229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32070" *)
  wire [7:0] _00230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31980" *)
  wire [7:0] _00231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32980" *)
  wire [7:0] _00232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32990" *)
  wire [7:0] _00233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33000" *)
  wire [7:0] _00234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33010" *)
  wire [7:0] _00235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33020" *)
  wire [7:0] _00236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33030" *)
  wire [7:0] _00237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33040" *)
  wire [7:0] _00238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33050" *)
  wire [7:0] _00239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33060" *)
  wire [7:0] _00240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33070" *)
  wire [7:0] _00241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32080" *)
  wire [7:0] _00242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33080" *)
  wire [7:0] _00243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33090" *)
  wire [7:0] _00244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33100" *)
  wire [7:0] _00245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33110" *)
  wire [7:0] _00246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33120" *)
  wire [7:0] _00247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33130" *)
  wire [7:0] _00248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33140" *)
  wire [7:0] _00249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33150" *)
  wire [7:0] _00250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33160" *)
  wire [7:0] _00251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33170" *)
  wire [7:0] _00252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32090" *)
  wire [7:0] _00253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33180" *)
  wire [7:0] _00254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33190" *)
  wire [7:0] _00255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33200" *)
  wire [7:0] _00256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33210" *)
  wire [7:0] _00257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33220" *)
  wire [7:0] _00258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34537" *)
  wire [7:0] _00259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34547" *)
  wire [7:0] _00260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34557" *)
  wire [7:0] _00261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33407" *)
  wire [7:0] _00262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33417" *)
  wire [7:0] _00263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33427" *)
  wire [7:0] _00264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33437" *)
  wire [7:0] _00265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33447" *)
  wire [7:0] _00266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33457" *)
  wire [7:0] _00267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33467" *)
  wire [7:0] _00268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33477" *)
  wire [7:0] _00269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33297" *)
  wire [7:0] _00270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33487" *)
  wire [7:0] _00271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33497" *)
  wire [7:0] _00272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33507" *)
  wire [7:0] _00273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33517" *)
  wire [7:0] _00274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33527" *)
  wire [7:0] _00275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33537" *)
  wire [7:0] _00276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33547" *)
  wire [7:0] _00277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33557" *)
  wire [7:0] _00278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33567" *)
  wire [7:0] _00279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33577" *)
  wire [7:0] _00280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33307" *)
  wire [7:0] _00281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33587" *)
  wire [7:0] _00282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33597" *)
  wire [7:0] _00283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33607" *)
  wire [7:0] _00284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33617" *)
  wire [7:0] _00285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33627" *)
  wire [7:0] _00286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33637" *)
  wire [7:0] _00287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33647" *)
  wire [7:0] _00288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33657" *)
  wire [7:0] _00289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33667" *)
  wire [7:0] _00290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33677" *)
  wire [7:0] _00291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33317" *)
  wire [7:0] _00292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33687" *)
  wire [7:0] _00293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33697" *)
  wire [7:0] _00294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33707" *)
  wire [7:0] _00295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33717" *)
  wire [7:0] _00296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33727" *)
  wire [7:0] _00297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33737" *)
  wire [7:0] _00298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33747" *)
  wire [7:0] _00299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33757" *)
  wire [7:0] _00300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33767" *)
  wire [7:0] _00301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33777" *)
  wire [7:0] _00302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33327" *)
  wire [7:0] _00303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33787" *)
  wire [7:0] _00304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33797" *)
  wire [7:0] _00305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33807" *)
  wire [7:0] _00306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33817" *)
  wire [7:0] _00307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33827" *)
  wire [7:0] _00308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33837" *)
  wire [7:0] _00309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33847" *)
  wire [7:0] _00310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33857" *)
  wire [7:0] _00311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33867" *)
  wire [7:0] _00312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33877" *)
  wire [7:0] _00313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33337" *)
  wire [7:0] _00314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33887" *)
  wire [7:0] _00315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33897" *)
  wire [7:0] _00316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33907" *)
  wire [7:0] _00317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33917" *)
  wire [7:0] _00318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33927" *)
  wire [7:0] _00319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33937" *)
  wire [7:0] _00320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33947" *)
  wire [7:0] _00321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33957" *)
  wire [7:0] _00322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33967" *)
  wire [7:0] _00323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33977" *)
  wire [7:0] _00324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33347" *)
  wire [7:0] _00325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33987" *)
  wire [7:0] _00326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33997" *)
  wire [7:0] _00327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34007" *)
  wire [7:0] _00328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34017" *)
  wire [7:0] _00329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34027" *)
  wire [7:0] _00330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34037" *)
  wire [7:0] _00331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34047" *)
  wire [7:0] _00332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34057" *)
  wire [7:0] _00333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34067" *)
  wire [7:0] _00334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34077" *)
  wire [7:0] _00335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33357" *)
  wire [7:0] _00336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34087" *)
  wire [7:0] _00337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34097" *)
  wire [7:0] _00338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34107" *)
  wire [7:0] _00339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34117" *)
  wire [7:0] _00340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34127" *)
  wire [7:0] _00341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34137" *)
  wire [7:0] _00342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34147" *)
  wire [7:0] _00343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34157" *)
  wire [7:0] _00344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34167" *)
  wire [7:0] _00345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34177" *)
  wire [7:0] _00346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33367" *)
  wire [7:0] _00347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34187" *)
  wire [7:0] _00348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34197" *)
  wire [7:0] _00349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34207" *)
  wire [7:0] _00350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34217" *)
  wire [7:0] _00351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34227" *)
  wire [7:0] _00352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34237" *)
  wire [7:0] _00353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34247" *)
  wire [7:0] _00354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34257" *)
  wire [7:0] _00355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34267" *)
  wire [7:0] _00356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34277" *)
  wire [7:0] _00357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33377" *)
  wire [7:0] _00358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33287" *)
  wire [7:0] _00359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34287" *)
  wire [7:0] _00360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34297" *)
  wire [7:0] _00361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34307" *)
  wire [7:0] _00362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34317" *)
  wire [7:0] _00363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34327" *)
  wire [7:0] _00364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34337" *)
  wire [7:0] _00365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34347" *)
  wire [7:0] _00366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34357" *)
  wire [7:0] _00367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34367" *)
  wire [7:0] _00368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34377" *)
  wire [7:0] _00369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33387" *)
  wire [7:0] _00370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34387" *)
  wire [7:0] _00371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34397" *)
  wire [7:0] _00372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34407" *)
  wire [7:0] _00373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34417" *)
  wire [7:0] _00374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34427" *)
  wire [7:0] _00375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34437" *)
  wire [7:0] _00376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34447" *)
  wire [7:0] _00377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34457" *)
  wire [7:0] _00378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34467" *)
  wire [7:0] _00379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34477" *)
  wire [7:0] _00380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33397" *)
  wire [7:0] _00381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34487" *)
  wire [7:0] _00382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34497" *)
  wire [7:0] _00383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34507" *)
  wire [7:0] _00384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34517" *)
  wire [7:0] _00385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34527" *)
  wire [7:0] _00386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35844" *)
  wire [7:0] _00387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35854" *)
  wire [7:0] _00388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35864" *)
  wire [7:0] _00389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34714" *)
  wire [7:0] _00390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34724" *)
  wire [7:0] _00391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34734" *)
  wire [7:0] _00392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34744" *)
  wire [7:0] _00393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34754" *)
  wire [7:0] _00394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34764" *)
  wire [7:0] _00395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34774" *)
  wire [7:0] _00396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34784" *)
  wire [7:0] _00397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34604" *)
  wire [7:0] _00398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34794" *)
  wire [7:0] _00399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34804" *)
  wire [7:0] _00400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34814" *)
  wire [7:0] _00401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34824" *)
  wire [7:0] _00402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34834" *)
  wire [7:0] _00403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34844" *)
  wire [7:0] _00404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34854" *)
  wire [7:0] _00405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34864" *)
  wire [7:0] _00406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34874" *)
  wire [7:0] _00407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34884" *)
  wire [7:0] _00408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34614" *)
  wire [7:0] _00409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34894" *)
  wire [7:0] _00410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34904" *)
  wire [7:0] _00411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34914" *)
  wire [7:0] _00412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34924" *)
  wire [7:0] _00413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34934" *)
  wire [7:0] _00414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34944" *)
  wire [7:0] _00415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34954" *)
  wire [7:0] _00416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34964" *)
  wire [7:0] _00417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34974" *)
  wire [7:0] _00418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34984" *)
  wire [7:0] _00419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34624" *)
  wire [7:0] _00420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34994" *)
  wire [7:0] _00421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35004" *)
  wire [7:0] _00422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35014" *)
  wire [7:0] _00423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35024" *)
  wire [7:0] _00424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35034" *)
  wire [7:0] _00425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35044" *)
  wire [7:0] _00426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35054" *)
  wire [7:0] _00427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35064" *)
  wire [7:0] _00428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35074" *)
  wire [7:0] _00429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35084" *)
  wire [7:0] _00430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34634" *)
  wire [7:0] _00431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35094" *)
  wire [7:0] _00432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35104" *)
  wire [7:0] _00433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35114" *)
  wire [7:0] _00434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35124" *)
  wire [7:0] _00435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35134" *)
  wire [7:0] _00436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35144" *)
  wire [7:0] _00437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35154" *)
  wire [7:0] _00438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35164" *)
  wire [7:0] _00439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35174" *)
  wire [7:0] _00440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35184" *)
  wire [7:0] _00441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34644" *)
  wire [7:0] _00442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35194" *)
  wire [7:0] _00443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35204" *)
  wire [7:0] _00444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35214" *)
  wire [7:0] _00445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35224" *)
  wire [7:0] _00446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35234" *)
  wire [7:0] _00447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35244" *)
  wire [7:0] _00448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35254" *)
  wire [7:0] _00449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35264" *)
  wire [7:0] _00450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35274" *)
  wire [7:0] _00451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35284" *)
  wire [7:0] _00452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34654" *)
  wire [7:0] _00453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35294" *)
  wire [7:0] _00454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35304" *)
  wire [7:0] _00455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35314" *)
  wire [7:0] _00456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35324" *)
  wire [7:0] _00457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35334" *)
  wire [7:0] _00458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35344" *)
  wire [7:0] _00459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35354" *)
  wire [7:0] _00460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35364" *)
  wire [7:0] _00461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35374" *)
  wire [7:0] _00462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35384" *)
  wire [7:0] _00463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34664" *)
  wire [7:0] _00464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35394" *)
  wire [7:0] _00465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35404" *)
  wire [7:0] _00466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35414" *)
  wire [7:0] _00467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35424" *)
  wire [7:0] _00468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35434" *)
  wire [7:0] _00469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35444" *)
  wire [7:0] _00470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35454" *)
  wire [7:0] _00471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35464" *)
  wire [7:0] _00472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35474" *)
  wire [7:0] _00473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35484" *)
  wire [7:0] _00474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34674" *)
  wire [7:0] _00475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35494" *)
  wire [7:0] _00476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35504" *)
  wire [7:0] _00477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35514" *)
  wire [7:0] _00478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35524" *)
  wire [7:0] _00479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35534" *)
  wire [7:0] _00480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35544" *)
  wire [7:0] _00481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35554" *)
  wire [7:0] _00482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35564" *)
  wire [7:0] _00483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35574" *)
  wire [7:0] _00484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35584" *)
  wire [7:0] _00485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34684" *)
  wire [7:0] _00486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34594" *)
  wire [7:0] _00487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35594" *)
  wire [7:0] _00488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35604" *)
  wire [7:0] _00489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35614" *)
  wire [7:0] _00490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35624" *)
  wire [7:0] _00491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35634" *)
  wire [7:0] _00492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35644" *)
  wire [7:0] _00493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35654" *)
  wire [7:0] _00494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35664" *)
  wire [7:0] _00495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35674" *)
  wire [7:0] _00496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35684" *)
  wire [7:0] _00497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34694" *)
  wire [7:0] _00498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35694" *)
  wire [7:0] _00499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35704" *)
  wire [7:0] _00500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35714" *)
  wire [7:0] _00501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35724" *)
  wire [7:0] _00502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35734" *)
  wire [7:0] _00503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35744" *)
  wire [7:0] _00504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35754" *)
  wire [7:0] _00505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35764" *)
  wire [7:0] _00506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35774" *)
  wire [7:0] _00507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35784" *)
  wire [7:0] _00508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34704" *)
  wire [7:0] _00509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35794" *)
  wire [7:0] _00510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35804" *)
  wire [7:0] _00511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35814" *)
  wire [7:0] _00512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35824" *)
  wire [7:0] _00513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35834" *)
  wire [7:0] _00514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37151" *)
  wire [7:0] _00515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37161" *)
  wire [7:0] _00516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37171" *)
  wire [7:0] _00517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36021" *)
  wire [7:0] _00518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36031" *)
  wire [7:0] _00519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36041" *)
  wire [7:0] _00520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36051" *)
  wire [7:0] _00521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36061" *)
  wire [7:0] _00522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36071" *)
  wire [7:0] _00523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36081" *)
  wire [7:0] _00524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36091" *)
  wire [7:0] _00525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35911" *)
  wire [7:0] _00526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36101" *)
  wire [7:0] _00527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36111" *)
  wire [7:0] _00528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36121" *)
  wire [7:0] _00529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36131" *)
  wire [7:0] _00530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36141" *)
  wire [7:0] _00531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36151" *)
  wire [7:0] _00532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36161" *)
  wire [7:0] _00533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36171" *)
  wire [7:0] _00534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36181" *)
  wire [7:0] _00535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36191" *)
  wire [7:0] _00536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35921" *)
  wire [7:0] _00537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36201" *)
  wire [7:0] _00538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36211" *)
  wire [7:0] _00539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36221" *)
  wire [7:0] _00540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36231" *)
  wire [7:0] _00541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36241" *)
  wire [7:0] _00542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36251" *)
  wire [7:0] _00543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36261" *)
  wire [7:0] _00544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36271" *)
  wire [7:0] _00545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36281" *)
  wire [7:0] _00546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36291" *)
  wire [7:0] _00547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35931" *)
  wire [7:0] _00548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36301" *)
  wire [7:0] _00549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36311" *)
  wire [7:0] _00550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36321" *)
  wire [7:0] _00551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36331" *)
  wire [7:0] _00552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36341" *)
  wire [7:0] _00553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36351" *)
  wire [7:0] _00554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36361" *)
  wire [7:0] _00555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36371" *)
  wire [7:0] _00556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36381" *)
  wire [7:0] _00557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36391" *)
  wire [7:0] _00558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35941" *)
  wire [7:0] _00559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36401" *)
  wire [7:0] _00560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36411" *)
  wire [7:0] _00561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36421" *)
  wire [7:0] _00562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36431" *)
  wire [7:0] _00563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36441" *)
  wire [7:0] _00564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36451" *)
  wire [7:0] _00565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36461" *)
  wire [7:0] _00566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36471" *)
  wire [7:0] _00567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36481" *)
  wire [7:0] _00568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36491" *)
  wire [7:0] _00569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35951" *)
  wire [7:0] _00570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36501" *)
  wire [7:0] _00571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36511" *)
  wire [7:0] _00572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36521" *)
  wire [7:0] _00573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36531" *)
  wire [7:0] _00574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36541" *)
  wire [7:0] _00575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36551" *)
  wire [7:0] _00576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36561" *)
  wire [7:0] _00577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36571" *)
  wire [7:0] _00578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36581" *)
  wire [7:0] _00579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36591" *)
  wire [7:0] _00580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35961" *)
  wire [7:0] _00581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36601" *)
  wire [7:0] _00582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36611" *)
  wire [7:0] _00583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36621" *)
  wire [7:0] _00584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36631" *)
  wire [7:0] _00585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36641" *)
  wire [7:0] _00586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36651" *)
  wire [7:0] _00587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36661" *)
  wire [7:0] _00588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36671" *)
  wire [7:0] _00589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36681" *)
  wire [7:0] _00590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36691" *)
  wire [7:0] _00591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35971" *)
  wire [7:0] _00592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36701" *)
  wire [7:0] _00593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36711" *)
  wire [7:0] _00594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36721" *)
  wire [7:0] _00595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36731" *)
  wire [7:0] _00596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36741" *)
  wire [7:0] _00597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36751" *)
  wire [7:0] _00598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36761" *)
  wire [7:0] _00599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36771" *)
  wire [7:0] _00600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36781" *)
  wire [7:0] _00601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36791" *)
  wire [7:0] _00602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35981" *)
  wire [7:0] _00603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36801" *)
  wire [7:0] _00604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36811" *)
  wire [7:0] _00605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36821" *)
  wire [7:0] _00606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36831" *)
  wire [7:0] _00607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36841" *)
  wire [7:0] _00608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36851" *)
  wire [7:0] _00609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36861" *)
  wire [7:0] _00610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36871" *)
  wire [7:0] _00611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36881" *)
  wire [7:0] _00612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36891" *)
  wire [7:0] _00613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35991" *)
  wire [7:0] _00614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35901" *)
  wire [7:0] _00615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36901" *)
  wire [7:0] _00616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36911" *)
  wire [7:0] _00617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36921" *)
  wire [7:0] _00618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36931" *)
  wire [7:0] _00619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36941" *)
  wire [7:0] _00620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36951" *)
  wire [7:0] _00621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36961" *)
  wire [7:0] _00622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36971" *)
  wire [7:0] _00623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36981" *)
  wire [7:0] _00624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36991" *)
  wire [7:0] _00625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36001" *)
  wire [7:0] _00626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37001" *)
  wire [7:0] _00627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37011" *)
  wire [7:0] _00628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37021" *)
  wire [7:0] _00629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37031" *)
  wire [7:0] _00630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37041" *)
  wire [7:0] _00631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37051" *)
  wire [7:0] _00632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37061" *)
  wire [7:0] _00633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37071" *)
  wire [7:0] _00634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37081" *)
  wire [7:0] _00635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37091" *)
  wire [7:0] _00636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36011" *)
  wire [7:0] _00637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37101" *)
  wire [7:0] _00638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37111" *)
  wire [7:0] _00639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37121" *)
  wire [7:0] _00640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37131" *)
  wire [7:0] _00641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37141" *)
  wire [7:0] _00642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38458" *)
  wire [7:0] _00643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38468" *)
  wire [7:0] _00644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38478" *)
  wire [7:0] _00645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37328" *)
  wire [7:0] _00646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37338" *)
  wire [7:0] _00647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37348" *)
  wire [7:0] _00648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37358" *)
  wire [7:0] _00649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37368" *)
  wire [7:0] _00650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37378" *)
  wire [7:0] _00651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37388" *)
  wire [7:0] _00652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37398" *)
  wire [7:0] _00653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37218" *)
  wire [7:0] _00654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37408" *)
  wire [7:0] _00655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37418" *)
  wire [7:0] _00656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37428" *)
  wire [7:0] _00657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37438" *)
  wire [7:0] _00658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37448" *)
  wire [7:0] _00659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37458" *)
  wire [7:0] _00660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37468" *)
  wire [7:0] _00661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37478" *)
  wire [7:0] _00662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37488" *)
  wire [7:0] _00663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37498" *)
  wire [7:0] _00664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37228" *)
  wire [7:0] _00665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37508" *)
  wire [7:0] _00666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37518" *)
  wire [7:0] _00667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37528" *)
  wire [7:0] _00668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37538" *)
  wire [7:0] _00669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37548" *)
  wire [7:0] _00670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37558" *)
  wire [7:0] _00671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37568" *)
  wire [7:0] _00672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37578" *)
  wire [7:0] _00673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37588" *)
  wire [7:0] _00674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37598" *)
  wire [7:0] _00675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37238" *)
  wire [7:0] _00676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37608" *)
  wire [7:0] _00677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37618" *)
  wire [7:0] _00678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37628" *)
  wire [7:0] _00679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37638" *)
  wire [7:0] _00680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37648" *)
  wire [7:0] _00681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37658" *)
  wire [7:0] _00682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37668" *)
  wire [7:0] _00683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37678" *)
  wire [7:0] _00684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37688" *)
  wire [7:0] _00685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37698" *)
  wire [7:0] _00686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37248" *)
  wire [7:0] _00687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37708" *)
  wire [7:0] _00688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37718" *)
  wire [7:0] _00689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37728" *)
  wire [7:0] _00690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37738" *)
  wire [7:0] _00691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37748" *)
  wire [7:0] _00692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37758" *)
  wire [7:0] _00693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37768" *)
  wire [7:0] _00694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37778" *)
  wire [7:0] _00695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37788" *)
  wire [7:0] _00696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37798" *)
  wire [7:0] _00697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37258" *)
  wire [7:0] _00698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37808" *)
  wire [7:0] _00699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37818" *)
  wire [7:0] _00700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37828" *)
  wire [7:0] _00701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37838" *)
  wire [7:0] _00702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37848" *)
  wire [7:0] _00703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37858" *)
  wire [7:0] _00704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37868" *)
  wire [7:0] _00705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37878" *)
  wire [7:0] _00706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37888" *)
  wire [7:0] _00707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37898" *)
  wire [7:0] _00708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37268" *)
  wire [7:0] _00709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37908" *)
  wire [7:0] _00710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37918" *)
  wire [7:0] _00711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37928" *)
  wire [7:0] _00712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37938" *)
  wire [7:0] _00713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37948" *)
  wire [7:0] _00714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37958" *)
  wire [7:0] _00715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37968" *)
  wire [7:0] _00716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37978" *)
  wire [7:0] _00717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37988" *)
  wire [7:0] _00718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37998" *)
  wire [7:0] _00719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37278" *)
  wire [7:0] _00720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38008" *)
  wire [7:0] _00721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38018" *)
  wire [7:0] _00722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38028" *)
  wire [7:0] _00723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38038" *)
  wire [7:0] _00724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38048" *)
  wire [7:0] _00725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38058" *)
  wire [7:0] _00726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38068" *)
  wire [7:0] _00727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38078" *)
  wire [7:0] _00728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38088" *)
  wire [7:0] _00729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38098" *)
  wire [7:0] _00730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37288" *)
  wire [7:0] _00731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38108" *)
  wire [7:0] _00732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38118" *)
  wire [7:0] _00733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38128" *)
  wire [7:0] _00734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38138" *)
  wire [7:0] _00735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38148" *)
  wire [7:0] _00736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38158" *)
  wire [7:0] _00737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38168" *)
  wire [7:0] _00738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38178" *)
  wire [7:0] _00739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38188" *)
  wire [7:0] _00740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38198" *)
  wire [7:0] _00741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37298" *)
  wire [7:0] _00742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37208" *)
  wire [7:0] _00743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38208" *)
  wire [7:0] _00744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38218" *)
  wire [7:0] _00745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38228" *)
  wire [7:0] _00746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38238" *)
  wire [7:0] _00747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38248" *)
  wire [7:0] _00748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38258" *)
  wire [7:0] _00749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38268" *)
  wire [7:0] _00750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38278" *)
  wire [7:0] _00751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38288" *)
  wire [7:0] _00752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38298" *)
  wire [7:0] _00753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37308" *)
  wire [7:0] _00754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38308" *)
  wire [7:0] _00755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38318" *)
  wire [7:0] _00756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38328" *)
  wire [7:0] _00757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38338" *)
  wire [7:0] _00758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38348" *)
  wire [7:0] _00759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38358" *)
  wire [7:0] _00760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38368" *)
  wire [7:0] _00761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38378" *)
  wire [7:0] _00762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38388" *)
  wire [7:0] _00763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38398" *)
  wire [7:0] _00764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37318" *)
  wire [7:0] _00765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38408" *)
  wire [7:0] _00766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38418" *)
  wire [7:0] _00767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38428" *)
  wire [7:0] _00768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38438" *)
  wire [7:0] _00769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38448" *)
  wire [7:0] _00770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39765" *)
  wire [7:0] _00771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39775" *)
  wire [7:0] _00772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39785" *)
  wire [7:0] _00773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38635" *)
  wire [7:0] _00774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38645" *)
  wire [7:0] _00775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38655" *)
  wire [7:0] _00776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38665" *)
  wire [7:0] _00777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38675" *)
  wire [7:0] _00778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38685" *)
  wire [7:0] _00779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38695" *)
  wire [7:0] _00780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38705" *)
  wire [7:0] _00781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38525" *)
  wire [7:0] _00782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38715" *)
  wire [7:0] _00783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38725" *)
  wire [7:0] _00784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38735" *)
  wire [7:0] _00785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38745" *)
  wire [7:0] _00786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38755" *)
  wire [7:0] _00787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38765" *)
  wire [7:0] _00788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38775" *)
  wire [7:0] _00789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38785" *)
  wire [7:0] _00790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38795" *)
  wire [7:0] _00791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38805" *)
  wire [7:0] _00792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38535" *)
  wire [7:0] _00793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38815" *)
  wire [7:0] _00794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38825" *)
  wire [7:0] _00795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38835" *)
  wire [7:0] _00796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38845" *)
  wire [7:0] _00797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38855" *)
  wire [7:0] _00798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38865" *)
  wire [7:0] _00799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38875" *)
  wire [7:0] _00800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38885" *)
  wire [7:0] _00801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38895" *)
  wire [7:0] _00802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38905" *)
  wire [7:0] _00803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38545" *)
  wire [7:0] _00804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38915" *)
  wire [7:0] _00805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38925" *)
  wire [7:0] _00806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38935" *)
  wire [7:0] _00807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38945" *)
  wire [7:0] _00808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38955" *)
  wire [7:0] _00809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38965" *)
  wire [7:0] _00810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38975" *)
  wire [7:0] _00811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38985" *)
  wire [7:0] _00812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38995" *)
  wire [7:0] _00813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39005" *)
  wire [7:0] _00814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38555" *)
  wire [7:0] _00815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39015" *)
  wire [7:0] _00816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39025" *)
  wire [7:0] _00817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39035" *)
  wire [7:0] _00818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39045" *)
  wire [7:0] _00819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39055" *)
  wire [7:0] _00820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39065" *)
  wire [7:0] _00821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39075" *)
  wire [7:0] _00822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39085" *)
  wire [7:0] _00823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39095" *)
  wire [7:0] _00824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39105" *)
  wire [7:0] _00825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38565" *)
  wire [7:0] _00826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39115" *)
  wire [7:0] _00827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39125" *)
  wire [7:0] _00828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39135" *)
  wire [7:0] _00829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39145" *)
  wire [7:0] _00830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39155" *)
  wire [7:0] _00831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39165" *)
  wire [7:0] _00832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39175" *)
  wire [7:0] _00833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39185" *)
  wire [7:0] _00834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39195" *)
  wire [7:0] _00835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39205" *)
  wire [7:0] _00836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38575" *)
  wire [7:0] _00837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39215" *)
  wire [7:0] _00838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39225" *)
  wire [7:0] _00839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39235" *)
  wire [7:0] _00840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39245" *)
  wire [7:0] _00841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39255" *)
  wire [7:0] _00842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39265" *)
  wire [7:0] _00843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39275" *)
  wire [7:0] _00844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39285" *)
  wire [7:0] _00845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39295" *)
  wire [7:0] _00846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39305" *)
  wire [7:0] _00847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38585" *)
  wire [7:0] _00848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39315" *)
  wire [7:0] _00849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39325" *)
  wire [7:0] _00850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39335" *)
  wire [7:0] _00851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39345" *)
  wire [7:0] _00852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39355" *)
  wire [7:0] _00853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39365" *)
  wire [7:0] _00854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39375" *)
  wire [7:0] _00855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39385" *)
  wire [7:0] _00856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39395" *)
  wire [7:0] _00857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39405" *)
  wire [7:0] _00858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38595" *)
  wire [7:0] _00859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39415" *)
  wire [7:0] _00860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39425" *)
  wire [7:0] _00861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39435" *)
  wire [7:0] _00862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39445" *)
  wire [7:0] _00863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39455" *)
  wire [7:0] _00864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39465" *)
  wire [7:0] _00865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39475" *)
  wire [7:0] _00866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39485" *)
  wire [7:0] _00867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39495" *)
  wire [7:0] _00868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39505" *)
  wire [7:0] _00869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38605" *)
  wire [7:0] _00870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38515" *)
  wire [7:0] _00871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39515" *)
  wire [7:0] _00872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39525" *)
  wire [7:0] _00873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39535" *)
  wire [7:0] _00874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39545" *)
  wire [7:0] _00875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39555" *)
  wire [7:0] _00876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39565" *)
  wire [7:0] _00877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39575" *)
  wire [7:0] _00878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39585" *)
  wire [7:0] _00879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39595" *)
  wire [7:0] _00880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39605" *)
  wire [7:0] _00881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38615" *)
  wire [7:0] _00882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39615" *)
  wire [7:0] _00883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39625" *)
  wire [7:0] _00884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39635" *)
  wire [7:0] _00885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39645" *)
  wire [7:0] _00886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39655" *)
  wire [7:0] _00887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39665" *)
  wire [7:0] _00888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39675" *)
  wire [7:0] _00889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39685" *)
  wire [7:0] _00890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39695" *)
  wire [7:0] _00891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39705" *)
  wire [7:0] _00892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38625" *)
  wire [7:0] _00893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39715" *)
  wire [7:0] _00894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39725" *)
  wire [7:0] _00895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39735" *)
  wire [7:0] _00896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39745" *)
  wire [7:0] _00897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39755" *)
  wire [7:0] _00898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41072" *)
  wire [7:0] _00899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41082" *)
  wire [7:0] _00900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41092" *)
  wire [7:0] _00901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39942" *)
  wire [7:0] _00902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39952" *)
  wire [7:0] _00903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39962" *)
  wire [7:0] _00904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39972" *)
  wire [7:0] _00905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39982" *)
  wire [7:0] _00906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39992" *)
  wire [7:0] _00907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40002" *)
  wire [7:0] _00908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40012" *)
  wire [7:0] _00909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39832" *)
  wire [7:0] _00910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40022" *)
  wire [7:0] _00911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40032" *)
  wire [7:0] _00912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40042" *)
  wire [7:0] _00913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40052" *)
  wire [7:0] _00914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40062" *)
  wire [7:0] _00915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40072" *)
  wire [7:0] _00916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40082" *)
  wire [7:0] _00917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40092" *)
  wire [7:0] _00918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40102" *)
  wire [7:0] _00919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40112" *)
  wire [7:0] _00920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39842" *)
  wire [7:0] _00921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40122" *)
  wire [7:0] _00922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40132" *)
  wire [7:0] _00923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40142" *)
  wire [7:0] _00924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40152" *)
  wire [7:0] _00925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40162" *)
  wire [7:0] _00926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40172" *)
  wire [7:0] _00927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40182" *)
  wire [7:0] _00928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40192" *)
  wire [7:0] _00929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40202" *)
  wire [7:0] _00930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40212" *)
  wire [7:0] _00931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39852" *)
  wire [7:0] _00932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40222" *)
  wire [7:0] _00933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40232" *)
  wire [7:0] _00934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40242" *)
  wire [7:0] _00935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40252" *)
  wire [7:0] _00936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40262" *)
  wire [7:0] _00937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40272" *)
  wire [7:0] _00938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40282" *)
  wire [7:0] _00939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40292" *)
  wire [7:0] _00940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40302" *)
  wire [7:0] _00941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40312" *)
  wire [7:0] _00942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39862" *)
  wire [7:0] _00943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40322" *)
  wire [7:0] _00944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40332" *)
  wire [7:0] _00945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40342" *)
  wire [7:0] _00946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40352" *)
  wire [7:0] _00947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40362" *)
  wire [7:0] _00948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40372" *)
  wire [7:0] _00949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40382" *)
  wire [7:0] _00950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40392" *)
  wire [7:0] _00951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40402" *)
  wire [7:0] _00952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40412" *)
  wire [7:0] _00953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39872" *)
  wire [7:0] _00954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40422" *)
  wire [7:0] _00955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40432" *)
  wire [7:0] _00956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40442" *)
  wire [7:0] _00957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40452" *)
  wire [7:0] _00958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40462" *)
  wire [7:0] _00959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40472" *)
  wire [7:0] _00960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40482" *)
  wire [7:0] _00961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40492" *)
  wire [7:0] _00962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40502" *)
  wire [7:0] _00963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40512" *)
  wire [7:0] _00964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39882" *)
  wire [7:0] _00965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40522" *)
  wire [7:0] _00966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40532" *)
  wire [7:0] _00967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40542" *)
  wire [7:0] _00968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40552" *)
  wire [7:0] _00969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40562" *)
  wire [7:0] _00970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40572" *)
  wire [7:0] _00971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40582" *)
  wire [7:0] _00972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40592" *)
  wire [7:0] _00973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40602" *)
  wire [7:0] _00974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40612" *)
  wire [7:0] _00975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39892" *)
  wire [7:0] _00976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40622" *)
  wire [7:0] _00977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40632" *)
  wire [7:0] _00978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40642" *)
  wire [7:0] _00979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40652" *)
  wire [7:0] _00980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40662" *)
  wire [7:0] _00981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40672" *)
  wire [7:0] _00982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40682" *)
  wire [7:0] _00983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40692" *)
  wire [7:0] _00984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40702" *)
  wire [7:0] _00985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40712" *)
  wire [7:0] _00986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39902" *)
  wire [7:0] _00987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40722" *)
  wire [7:0] _00988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40732" *)
  wire [7:0] _00989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40742" *)
  wire [7:0] _00990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40752" *)
  wire [7:0] _00991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40762" *)
  wire [7:0] _00992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40772" *)
  wire [7:0] _00993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40782" *)
  wire [7:0] _00994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40792" *)
  wire [7:0] _00995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40802" *)
  wire [7:0] _00996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40812" *)
  wire [7:0] _00997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39912" *)
  wire [7:0] _00998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39822" *)
  wire [7:0] _00999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40822" *)
  wire [7:0] _01000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40832" *)
  wire [7:0] _01001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40842" *)
  wire [7:0] _01002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40852" *)
  wire [7:0] _01003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40862" *)
  wire [7:0] _01004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40872" *)
  wire [7:0] _01005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40882" *)
  wire [7:0] _01006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40892" *)
  wire [7:0] _01007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40902" *)
  wire [7:0] _01008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40912" *)
  wire [7:0] _01009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39922" *)
  wire [7:0] _01010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40922" *)
  wire [7:0] _01011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40932" *)
  wire [7:0] _01012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40942" *)
  wire [7:0] _01013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40952" *)
  wire [7:0] _01014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40962" *)
  wire [7:0] _01015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40972" *)
  wire [7:0] _01016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40982" *)
  wire [7:0] _01017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40992" *)
  wire [7:0] _01018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41002" *)
  wire [7:0] _01019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41012" *)
  wire [7:0] _01020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39932" *)
  wire [7:0] _01021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41022" *)
  wire [7:0] _01022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41032" *)
  wire [7:0] _01023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41042" *)
  wire [7:0] _01024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41052" *)
  wire [7:0] _01025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41062" *)
  wire [7:0] _01026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30663" *)
  wire [63:0] _01027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31970" *)
  wire [63:0] _01028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33277" *)
  wire [63:0] _01029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34584" *)
  wire [63:0] _01030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35891" *)
  wire [63:0] _01031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37198" *)
  wire [63:0] _01032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38505" *)
  wire [63:0] _01033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39812" *)
  wire [63:0] _01034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30653" *)
  wire [127:0] _01035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31960" *)
  wire [127:0] _01036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33267" *)
  wire [127:0] _01037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34574" *)
  wire [127:0] _01038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35881" *)
  wire [127:0] _01039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37188" *)
  wire [127:0] _01040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38495" *)
  wire [127:0] _01041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39802" *)
  wire [127:0] _01042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30335" *)
  wire [7:0] _01043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30345" *)
  wire [7:0] _01044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30355" *)
  wire [7:0] _01045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29205" *)
  wire [7:0] _01046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29215" *)
  wire [7:0] _01047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29225" *)
  wire [7:0] _01048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29235" *)
  wire [7:0] _01049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29245" *)
  wire [7:0] _01050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29255" *)
  wire [7:0] _01051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29265" *)
  wire [7:0] _01052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29275" *)
  wire [7:0] _01053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29095" *)
  wire [7:0] _01054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29285" *)
  wire [7:0] _01055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29295" *)
  wire [7:0] _01056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29305" *)
  wire [7:0] _01057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29315" *)
  wire [7:0] _01058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29325" *)
  wire [7:0] _01059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29335" *)
  wire [7:0] _01060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29345" *)
  wire [7:0] _01061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29355" *)
  wire [7:0] _01062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29365" *)
  wire [7:0] _01063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29375" *)
  wire [7:0] _01064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29105" *)
  wire [7:0] _01065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29385" *)
  wire [7:0] _01066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29395" *)
  wire [7:0] _01067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29405" *)
  wire [7:0] _01068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29415" *)
  wire [7:0] _01069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29425" *)
  wire [7:0] _01070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29435" *)
  wire [7:0] _01071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29445" *)
  wire [7:0] _01072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29455" *)
  wire [7:0] _01073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29465" *)
  wire [7:0] _01074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29475" *)
  wire [7:0] _01075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29115" *)
  wire [7:0] _01076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29485" *)
  wire [7:0] _01077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29495" *)
  wire [7:0] _01078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29505" *)
  wire [7:0] _01079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29515" *)
  wire [7:0] _01080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29525" *)
  wire [7:0] _01081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29535" *)
  wire [7:0] _01082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29545" *)
  wire [7:0] _01083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29555" *)
  wire [7:0] _01084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29565" *)
  wire [7:0] _01085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29575" *)
  wire [7:0] _01086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29125" *)
  wire [7:0] _01087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29585" *)
  wire [7:0] _01088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29595" *)
  wire [7:0] _01089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29605" *)
  wire [7:0] _01090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29615" *)
  wire [7:0] _01091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29625" *)
  wire [7:0] _01092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29635" *)
  wire [7:0] _01093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29645" *)
  wire [7:0] _01094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29655" *)
  wire [7:0] _01095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29665" *)
  wire [7:0] _01096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29675" *)
  wire [7:0] _01097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29135" *)
  wire [7:0] _01098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29685" *)
  wire [7:0] _01099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29695" *)
  wire [7:0] _01100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29705" *)
  wire [7:0] _01101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29715" *)
  wire [7:0] _01102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29725" *)
  wire [7:0] _01103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29735" *)
  wire [7:0] _01104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29745" *)
  wire [7:0] _01105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29755" *)
  wire [7:0] _01106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29765" *)
  wire [7:0] _01107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29775" *)
  wire [7:0] _01108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29145" *)
  wire [7:0] _01109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29785" *)
  wire [7:0] _01110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29795" *)
  wire [7:0] _01111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29805" *)
  wire [7:0] _01112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29815" *)
  wire [7:0] _01113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29825" *)
  wire [7:0] _01114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29835" *)
  wire [7:0] _01115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29845" *)
  wire [7:0] _01116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29855" *)
  wire [7:0] _01117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29865" *)
  wire [7:0] _01118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29875" *)
  wire [7:0] _01119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29155" *)
  wire [7:0] _01120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29885" *)
  wire [7:0] _01121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29895" *)
  wire [7:0] _01122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29905" *)
  wire [7:0] _01123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29915" *)
  wire [7:0] _01124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29925" *)
  wire [7:0] _01125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29935" *)
  wire [7:0] _01126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29945" *)
  wire [7:0] _01127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29955" *)
  wire [7:0] _01128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29965" *)
  wire [7:0] _01129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29975" *)
  wire [7:0] _01130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29165" *)
  wire [7:0] _01131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29985" *)
  wire [7:0] _01132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29995" *)
  wire [7:0] _01133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30005" *)
  wire [7:0] _01134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30015" *)
  wire [7:0] _01135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30025" *)
  wire [7:0] _01136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30035" *)
  wire [7:0] _01137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30045" *)
  wire [7:0] _01138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30055" *)
  wire [7:0] _01139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30065" *)
  wire [7:0] _01140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30075" *)
  wire [7:0] _01141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29175" *)
  wire [7:0] _01142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29085" *)
  wire [7:0] _01143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30085" *)
  wire [7:0] _01144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30095" *)
  wire [7:0] _01145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30105" *)
  wire [7:0] _01146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30115" *)
  wire [7:0] _01147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30125" *)
  wire [7:0] _01148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30135" *)
  wire [7:0] _01149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30145" *)
  wire [7:0] _01150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30155" *)
  wire [7:0] _01151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30165" *)
  wire [7:0] _01152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30175" *)
  wire [7:0] _01153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29185" *)
  wire [7:0] _01154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30185" *)
  wire [7:0] _01155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30195" *)
  wire [7:0] _01156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30205" *)
  wire [7:0] _01157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30215" *)
  wire [7:0] _01158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30225" *)
  wire [7:0] _01159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30235" *)
  wire [7:0] _01160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30245" *)
  wire [7:0] _01161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30255" *)
  wire [7:0] _01162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30265" *)
  wire [7:0] _01163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30275" *)
  wire [7:0] _01164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29195" *)
  wire [7:0] _01165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30285" *)
  wire [7:0] _01166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30295" *)
  wire [7:0] _01167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30305" *)
  wire [7:0] _01168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30315" *)
  wire [7:0] _01169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30325" *)
  wire [7:0] _01170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30389" *)
  wire [191:0] _01171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30409" *)
  wire [191:0] _01172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30429" *)
  wire [191:0] _01173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30449" *)
  wire [191:0] _01174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30469" *)
  wire [191:0] _01175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30489" *)
  wire [191:0] _01176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30509" *)
  wire [191:0] _01177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30529" *)
  wire [191:0] _01178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30379" *)
  wire [63:0] _01179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30399" *)
  wire [63:0] _01180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30419" *)
  wire [63:0] _01181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30439" *)
  wire [63:0] _01182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30459" *)
  wire [63:0] _01183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30479" *)
  wire [63:0] _01184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30499" *)
  wire [63:0] _01185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30519" *)
  wire [63:0] _01186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29075" *)
  wire [63:0] _01187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29065" *)
  wire [127:0] _01188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30372" *)
  wire [8:0] _01189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30365" *)
  wire [15:0] _01190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17297" *)
  wire [7:0] _01191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17307" *)
  wire [7:0] _01192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17317" *)
  wire [7:0] _01193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16167" *)
  wire [7:0] _01194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16177" *)
  wire [7:0] _01195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16187" *)
  wire [7:0] _01196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16197" *)
  wire [7:0] _01197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16207" *)
  wire [7:0] _01198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16217" *)
  wire [7:0] _01199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16227" *)
  wire [7:0] _01200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16237" *)
  wire [7:0] _01201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16057" *)
  wire [7:0] _01202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16247" *)
  wire [7:0] _01203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16257" *)
  wire [7:0] _01204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16267" *)
  wire [7:0] _01205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16277" *)
  wire [7:0] _01206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16287" *)
  wire [7:0] _01207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16297" *)
  wire [7:0] _01208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16307" *)
  wire [7:0] _01209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16317" *)
  wire [7:0] _01210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16327" *)
  wire [7:0] _01211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16337" *)
  wire [7:0] _01212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16067" *)
  wire [7:0] _01213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16347" *)
  wire [7:0] _01214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16357" *)
  wire [7:0] _01215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16367" *)
  wire [7:0] _01216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16377" *)
  wire [7:0] _01217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16387" *)
  wire [7:0] _01218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16397" *)
  wire [7:0] _01219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16407" *)
  wire [7:0] _01220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16417" *)
  wire [7:0] _01221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16427" *)
  wire [7:0] _01222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16437" *)
  wire [7:0] _01223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16077" *)
  wire [7:0] _01224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16447" *)
  wire [7:0] _01225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16457" *)
  wire [7:0] _01226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16467" *)
  wire [7:0] _01227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16477" *)
  wire [7:0] _01228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16487" *)
  wire [7:0] _01229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16497" *)
  wire [7:0] _01230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16507" *)
  wire [7:0] _01231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16517" *)
  wire [7:0] _01232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16527" *)
  wire [7:0] _01233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16537" *)
  wire [7:0] _01234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16087" *)
  wire [7:0] _01235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16547" *)
  wire [7:0] _01236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16557" *)
  wire [7:0] _01237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16567" *)
  wire [7:0] _01238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16577" *)
  wire [7:0] _01239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16587" *)
  wire [7:0] _01240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16597" *)
  wire [7:0] _01241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16607" *)
  wire [7:0] _01242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16617" *)
  wire [7:0] _01243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16627" *)
  wire [7:0] _01244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16637" *)
  wire [7:0] _01245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16097" *)
  wire [7:0] _01246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16647" *)
  wire [7:0] _01247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16657" *)
  wire [7:0] _01248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16667" *)
  wire [7:0] _01249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16677" *)
  wire [7:0] _01250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16687" *)
  wire [7:0] _01251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16697" *)
  wire [7:0] _01252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16707" *)
  wire [7:0] _01253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16717" *)
  wire [7:0] _01254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16727" *)
  wire [7:0] _01255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16737" *)
  wire [7:0] _01256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16107" *)
  wire [7:0] _01257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16747" *)
  wire [7:0] _01258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16757" *)
  wire [7:0] _01259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16767" *)
  wire [7:0] _01260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16777" *)
  wire [7:0] _01261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16787" *)
  wire [7:0] _01262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16797" *)
  wire [7:0] _01263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16807" *)
  wire [7:0] _01264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16817" *)
  wire [7:0] _01265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16827" *)
  wire [7:0] _01266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16837" *)
  wire [7:0] _01267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16117" *)
  wire [7:0] _01268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16847" *)
  wire [7:0] _01269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16857" *)
  wire [7:0] _01270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16867" *)
  wire [7:0] _01271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16877" *)
  wire [7:0] _01272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16887" *)
  wire [7:0] _01273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16897" *)
  wire [7:0] _01274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16907" *)
  wire [7:0] _01275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16917" *)
  wire [7:0] _01276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16927" *)
  wire [7:0] _01277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16937" *)
  wire [7:0] _01278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16127" *)
  wire [7:0] _01279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16947" *)
  wire [7:0] _01280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16957" *)
  wire [7:0] _01281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16967" *)
  wire [7:0] _01282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16977" *)
  wire [7:0] _01283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16987" *)
  wire [7:0] _01284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16997" *)
  wire [7:0] _01285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17007" *)
  wire [7:0] _01286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17017" *)
  wire [7:0] _01287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17027" *)
  wire [7:0] _01288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17037" *)
  wire [7:0] _01289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16137" *)
  wire [7:0] _01290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16047" *)
  wire [7:0] _01291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17047" *)
  wire [7:0] _01292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17057" *)
  wire [7:0] _01293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17067" *)
  wire [7:0] _01294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17077" *)
  wire [7:0] _01295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17087" *)
  wire [7:0] _01296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17097" *)
  wire [7:0] _01297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17107" *)
  wire [7:0] _01298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17117" *)
  wire [7:0] _01299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17127" *)
  wire [7:0] _01300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17137" *)
  wire [7:0] _01301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16147" *)
  wire [7:0] _01302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17147" *)
  wire [7:0] _01303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17157" *)
  wire [7:0] _01304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17167" *)
  wire [7:0] _01305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17177" *)
  wire [7:0] _01306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17187" *)
  wire [7:0] _01307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17197" *)
  wire [7:0] _01308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17207" *)
  wire [7:0] _01309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17217" *)
  wire [7:0] _01310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17227" *)
  wire [7:0] _01311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17237" *)
  wire [7:0] _01312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16157" *)
  wire [7:0] _01313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17247" *)
  wire [7:0] _01314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17257" *)
  wire [7:0] _01315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17267" *)
  wire [7:0] _01316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17277" *)
  wire [7:0] _01317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17287" *)
  wire [7:0] _01318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16037" *)
  wire [63:0] _01319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16027" *)
  wire [127:0] _01320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6621" *)
  wire [7:0] _01321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6631" *)
  wire [7:0] _01322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6641" *)
  wire [7:0] _01323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5491" *)
  wire [7:0] _01324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5501" *)
  wire [7:0] _01325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5511" *)
  wire [7:0] _01326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5521" *)
  wire [7:0] _01327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5531" *)
  wire [7:0] _01328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5541" *)
  wire [7:0] _01329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5551" *)
  wire [7:0] _01330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5561" *)
  wire [7:0] _01331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5381" *)
  wire [7:0] _01332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5571" *)
  wire [7:0] _01333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5581" *)
  wire [7:0] _01334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5591" *)
  wire [7:0] _01335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5601" *)
  wire [7:0] _01336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5611" *)
  wire [7:0] _01337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5621" *)
  wire [7:0] _01338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5631" *)
  wire [7:0] _01339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5641" *)
  wire [7:0] _01340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5651" *)
  wire [7:0] _01341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5661" *)
  wire [7:0] _01342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5391" *)
  wire [7:0] _01343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5671" *)
  wire [7:0] _01344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5681" *)
  wire [7:0] _01345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5691" *)
  wire [7:0] _01346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5701" *)
  wire [7:0] _01347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5711" *)
  wire [7:0] _01348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5721" *)
  wire [7:0] _01349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5731" *)
  wire [7:0] _01350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5741" *)
  wire [7:0] _01351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5751" *)
  wire [7:0] _01352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5761" *)
  wire [7:0] _01353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5401" *)
  wire [7:0] _01354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5771" *)
  wire [7:0] _01355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5781" *)
  wire [7:0] _01356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5791" *)
  wire [7:0] _01357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5801" *)
  wire [7:0] _01358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5811" *)
  wire [7:0] _01359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5821" *)
  wire [7:0] _01360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5831" *)
  wire [7:0] _01361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5841" *)
  wire [7:0] _01362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5851" *)
  wire [7:0] _01363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5861" *)
  wire [7:0] _01364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5411" *)
  wire [7:0] _01365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5871" *)
  wire [7:0] _01366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5881" *)
  wire [7:0] _01367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5891" *)
  wire [7:0] _01368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5901" *)
  wire [7:0] _01369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5911" *)
  wire [7:0] _01370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5921" *)
  wire [7:0] _01371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5931" *)
  wire [7:0] _01372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5941" *)
  wire [7:0] _01373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5951" *)
  wire [7:0] _01374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5961" *)
  wire [7:0] _01375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5421" *)
  wire [7:0] _01376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5971" *)
  wire [7:0] _01377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5981" *)
  wire [7:0] _01378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5991" *)
  wire [7:0] _01379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6001" *)
  wire [7:0] _01380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6011" *)
  wire [7:0] _01381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6021" *)
  wire [7:0] _01382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6031" *)
  wire [7:0] _01383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6041" *)
  wire [7:0] _01384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6051" *)
  wire [7:0] _01385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6061" *)
  wire [7:0] _01386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5431" *)
  wire [7:0] _01387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6071" *)
  wire [7:0] _01388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6081" *)
  wire [7:0] _01389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6091" *)
  wire [7:0] _01390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6101" *)
  wire [7:0] _01391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6111" *)
  wire [7:0] _01392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6121" *)
  wire [7:0] _01393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6131" *)
  wire [7:0] _01394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6141" *)
  wire [7:0] _01395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6151" *)
  wire [7:0] _01396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6161" *)
  wire [7:0] _01397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5441" *)
  wire [7:0] _01398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6171" *)
  wire [7:0] _01399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6181" *)
  wire [7:0] _01400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6191" *)
  wire [7:0] _01401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6201" *)
  wire [7:0] _01402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6211" *)
  wire [7:0] _01403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6221" *)
  wire [7:0] _01404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6231" *)
  wire [7:0] _01405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6241" *)
  wire [7:0] _01406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6251" *)
  wire [7:0] _01407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6261" *)
  wire [7:0] _01408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5451" *)
  wire [7:0] _01409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6271" *)
  wire [7:0] _01410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6281" *)
  wire [7:0] _01411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6291" *)
  wire [7:0] _01412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6301" *)
  wire [7:0] _01413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6311" *)
  wire [7:0] _01414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6321" *)
  wire [7:0] _01415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6331" *)
  wire [7:0] _01416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6341" *)
  wire [7:0] _01417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6351" *)
  wire [7:0] _01418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6361" *)
  wire [7:0] _01419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5461" *)
  wire [7:0] _01420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5371" *)
  wire [7:0] _01421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6371" *)
  wire [7:0] _01422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6381" *)
  wire [7:0] _01423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6391" *)
  wire [7:0] _01424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6401" *)
  wire [7:0] _01425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6411" *)
  wire [7:0] _01426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6421" *)
  wire [7:0] _01427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6431" *)
  wire [7:0] _01428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6441" *)
  wire [7:0] _01429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6451" *)
  wire [7:0] _01430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6461" *)
  wire [7:0] _01431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5471" *)
  wire [7:0] _01432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6471" *)
  wire [7:0] _01433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6481" *)
  wire [7:0] _01434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6491" *)
  wire [7:0] _01435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6501" *)
  wire [7:0] _01436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6511" *)
  wire [7:0] _01437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6521" *)
  wire [7:0] _01438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6531" *)
  wire [7:0] _01439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6541" *)
  wire [7:0] _01440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6551" *)
  wire [7:0] _01441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6561" *)
  wire [7:0] _01442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5481" *)
  wire [7:0] _01443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6571" *)
  wire [7:0] _01444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6581" *)
  wire [7:0] _01445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6591" *)
  wire [7:0] _01446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6601" *)
  wire [7:0] _01447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6611" *)
  wire [7:0] _01448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5351" *)
  wire [191:0] _01449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5341" *)
  wire [63:0] _01450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5361" *)
  wire [63:0] _01451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5331" *)
  wire [127:0] _01452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18621" *)
  wire [7:0] _01453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18631" *)
  wire [7:0] _01454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18641" *)
  wire [7:0] _01455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17491" *)
  wire [7:0] _01456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17501" *)
  wire [7:0] _01457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17511" *)
  wire [7:0] _01458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17521" *)
  wire [7:0] _01459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17531" *)
  wire [7:0] _01460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17541" *)
  wire [7:0] _01461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17551" *)
  wire [7:0] _01462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17561" *)
  wire [7:0] _01463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17381" *)
  wire [7:0] _01464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17571" *)
  wire [7:0] _01465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17581" *)
  wire [7:0] _01466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17591" *)
  wire [7:0] _01467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17601" *)
  wire [7:0] _01468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17611" *)
  wire [7:0] _01469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17621" *)
  wire [7:0] _01470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17631" *)
  wire [7:0] _01471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17641" *)
  wire [7:0] _01472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17651" *)
  wire [7:0] _01473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17661" *)
  wire [7:0] _01474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17391" *)
  wire [7:0] _01475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17671" *)
  wire [7:0] _01476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17681" *)
  wire [7:0] _01477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17691" *)
  wire [7:0] _01478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17701" *)
  wire [7:0] _01479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17711" *)
  wire [7:0] _01480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17721" *)
  wire [7:0] _01481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17731" *)
  wire [7:0] _01482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17741" *)
  wire [7:0] _01483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17751" *)
  wire [7:0] _01484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17761" *)
  wire [7:0] _01485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17401" *)
  wire [7:0] _01486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17771" *)
  wire [7:0] _01487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17781" *)
  wire [7:0] _01488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17791" *)
  wire [7:0] _01489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17801" *)
  wire [7:0] _01490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17811" *)
  wire [7:0] _01491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17821" *)
  wire [7:0] _01492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17831" *)
  wire [7:0] _01493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17841" *)
  wire [7:0] _01494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17851" *)
  wire [7:0] _01495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17861" *)
  wire [7:0] _01496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17411" *)
  wire [7:0] _01497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17871" *)
  wire [7:0] _01498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17881" *)
  wire [7:0] _01499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17891" *)
  wire [7:0] _01500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17901" *)
  wire [7:0] _01501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17911" *)
  wire [7:0] _01502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17921" *)
  wire [7:0] _01503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17931" *)
  wire [7:0] _01504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17941" *)
  wire [7:0] _01505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17951" *)
  wire [7:0] _01506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17961" *)
  wire [7:0] _01507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17421" *)
  wire [7:0] _01508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17971" *)
  wire [7:0] _01509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17981" *)
  wire [7:0] _01510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17991" *)
  wire [7:0] _01511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18001" *)
  wire [7:0] _01512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18011" *)
  wire [7:0] _01513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18021" *)
  wire [7:0] _01514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18031" *)
  wire [7:0] _01515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18041" *)
  wire [7:0] _01516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18051" *)
  wire [7:0] _01517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18061" *)
  wire [7:0] _01518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17431" *)
  wire [7:0] _01519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18071" *)
  wire [7:0] _01520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18081" *)
  wire [7:0] _01521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18091" *)
  wire [7:0] _01522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18101" *)
  wire [7:0] _01523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18111" *)
  wire [7:0] _01524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18121" *)
  wire [7:0] _01525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18131" *)
  wire [7:0] _01526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18141" *)
  wire [7:0] _01527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18151" *)
  wire [7:0] _01528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18161" *)
  wire [7:0] _01529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17441" *)
  wire [7:0] _01530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18171" *)
  wire [7:0] _01531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18181" *)
  wire [7:0] _01532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18191" *)
  wire [7:0] _01533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18201" *)
  wire [7:0] _01534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18211" *)
  wire [7:0] _01535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18221" *)
  wire [7:0] _01536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18231" *)
  wire [7:0] _01537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18241" *)
  wire [7:0] _01538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18251" *)
  wire [7:0] _01539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18261" *)
  wire [7:0] _01540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17451" *)
  wire [7:0] _01541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18271" *)
  wire [7:0] _01542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18281" *)
  wire [7:0] _01543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18291" *)
  wire [7:0] _01544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18301" *)
  wire [7:0] _01545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18311" *)
  wire [7:0] _01546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18321" *)
  wire [7:0] _01547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18331" *)
  wire [7:0] _01548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18341" *)
  wire [7:0] _01549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18351" *)
  wire [7:0] _01550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18361" *)
  wire [7:0] _01551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17461" *)
  wire [7:0] _01552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17371" *)
  wire [7:0] _01553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18371" *)
  wire [7:0] _01554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18381" *)
  wire [7:0] _01555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18391" *)
  wire [7:0] _01556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18401" *)
  wire [7:0] _01557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18411" *)
  wire [7:0] _01558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18421" *)
  wire [7:0] _01559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18431" *)
  wire [7:0] _01560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18441" *)
  wire [7:0] _01561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18451" *)
  wire [7:0] _01562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18461" *)
  wire [7:0] _01563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17471" *)
  wire [7:0] _01564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18471" *)
  wire [7:0] _01565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18481" *)
  wire [7:0] _01566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18491" *)
  wire [7:0] _01567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18501" *)
  wire [7:0] _01568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18511" *)
  wire [7:0] _01569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18521" *)
  wire [7:0] _01570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18531" *)
  wire [7:0] _01571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18541" *)
  wire [7:0] _01572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18551" *)
  wire [7:0] _01573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18561" *)
  wire [7:0] _01574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17481" *)
  wire [7:0] _01575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18571" *)
  wire [7:0] _01576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18581" *)
  wire [7:0] _01577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18591" *)
  wire [7:0] _01578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18601" *)
  wire [7:0] _01579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18611" *)
  wire [7:0] _01580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17361" *)
  wire [63:0] _01581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17351" *)
  wire [127:0] _01582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7957" *)
  wire [7:0] _01583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7967" *)
  wire [7:0] _01584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7977" *)
  wire [7:0] _01585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6827" *)
  wire [7:0] _01586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6837" *)
  wire [7:0] _01587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6847" *)
  wire [7:0] _01588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6857" *)
  wire [7:0] _01589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6867" *)
  wire [7:0] _01590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6877" *)
  wire [7:0] _01591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6887" *)
  wire [7:0] _01592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6897" *)
  wire [7:0] _01593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6717" *)
  wire [7:0] _01594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6907" *)
  wire [7:0] _01595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6917" *)
  wire [7:0] _01596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6927" *)
  wire [7:0] _01597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6937" *)
  wire [7:0] _01598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6947" *)
  wire [7:0] _01599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6957" *)
  wire [7:0] _01600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6967" *)
  wire [7:0] _01601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6977" *)
  wire [7:0] _01602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6987" *)
  wire [7:0] _01603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6997" *)
  wire [7:0] _01604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6727" *)
  wire [7:0] _01605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7007" *)
  wire [7:0] _01606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7017" *)
  wire [7:0] _01607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7027" *)
  wire [7:0] _01608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7037" *)
  wire [7:0] _01609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7047" *)
  wire [7:0] _01610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7057" *)
  wire [7:0] _01611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7067" *)
  wire [7:0] _01612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7077" *)
  wire [7:0] _01613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7087" *)
  wire [7:0] _01614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7097" *)
  wire [7:0] _01615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6737" *)
  wire [7:0] _01616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7107" *)
  wire [7:0] _01617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7117" *)
  wire [7:0] _01618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7127" *)
  wire [7:0] _01619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7137" *)
  wire [7:0] _01620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7147" *)
  wire [7:0] _01621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7157" *)
  wire [7:0] _01622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7167" *)
  wire [7:0] _01623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7177" *)
  wire [7:0] _01624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7187" *)
  wire [7:0] _01625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7197" *)
  wire [7:0] _01626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6747" *)
  wire [7:0] _01627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7207" *)
  wire [7:0] _01628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7217" *)
  wire [7:0] _01629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7227" *)
  wire [7:0] _01630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7237" *)
  wire [7:0] _01631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7247" *)
  wire [7:0] _01632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7257" *)
  wire [7:0] _01633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7267" *)
  wire [7:0] _01634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7277" *)
  wire [7:0] _01635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7287" *)
  wire [7:0] _01636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7297" *)
  wire [7:0] _01637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6757" *)
  wire [7:0] _01638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7307" *)
  wire [7:0] _01639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7317" *)
  wire [7:0] _01640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7327" *)
  wire [7:0] _01641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7337" *)
  wire [7:0] _01642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7347" *)
  wire [7:0] _01643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7357" *)
  wire [7:0] _01644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7367" *)
  wire [7:0] _01645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7377" *)
  wire [7:0] _01646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7387" *)
  wire [7:0] _01647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7397" *)
  wire [7:0] _01648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6767" *)
  wire [7:0] _01649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7407" *)
  wire [7:0] _01650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7417" *)
  wire [7:0] _01651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7427" *)
  wire [7:0] _01652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7437" *)
  wire [7:0] _01653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7447" *)
  wire [7:0] _01654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7457" *)
  wire [7:0] _01655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7467" *)
  wire [7:0] _01656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7477" *)
  wire [7:0] _01657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7487" *)
  wire [7:0] _01658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7497" *)
  wire [7:0] _01659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6777" *)
  wire [7:0] _01660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7507" *)
  wire [7:0] _01661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7517" *)
  wire [7:0] _01662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7527" *)
  wire [7:0] _01663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7537" *)
  wire [7:0] _01664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7547" *)
  wire [7:0] _01665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7557" *)
  wire [7:0] _01666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7567" *)
  wire [7:0] _01667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7577" *)
  wire [7:0] _01668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7587" *)
  wire [7:0] _01669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7597" *)
  wire [7:0] _01670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6787" *)
  wire [7:0] _01671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7607" *)
  wire [7:0] _01672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7617" *)
  wire [7:0] _01673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7627" *)
  wire [7:0] _01674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7637" *)
  wire [7:0] _01675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7647" *)
  wire [7:0] _01676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7657" *)
  wire [7:0] _01677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7667" *)
  wire [7:0] _01678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7677" *)
  wire [7:0] _01679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7687" *)
  wire [7:0] _01680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7697" *)
  wire [7:0] _01681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6797" *)
  wire [7:0] _01682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6707" *)
  wire [7:0] _01683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7707" *)
  wire [7:0] _01684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7717" *)
  wire [7:0] _01685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7727" *)
  wire [7:0] _01686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7737" *)
  wire [7:0] _01687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7747" *)
  wire [7:0] _01688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7757" *)
  wire [7:0] _01689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7767" *)
  wire [7:0] _01690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7777" *)
  wire [7:0] _01691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7787" *)
  wire [7:0] _01692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7797" *)
  wire [7:0] _01693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6807" *)
  wire [7:0] _01694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7807" *)
  wire [7:0] _01695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7817" *)
  wire [7:0] _01696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7827" *)
  wire [7:0] _01697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7837" *)
  wire [7:0] _01698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7847" *)
  wire [7:0] _01699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7857" *)
  wire [7:0] _01700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7867" *)
  wire [7:0] _01701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7877" *)
  wire [7:0] _01702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7887" *)
  wire [7:0] _01703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7897" *)
  wire [7:0] _01704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6817" *)
  wire [7:0] _01705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7907" *)
  wire [7:0] _01706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7917" *)
  wire [7:0] _01707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7927" *)
  wire [7:0] _01708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7937" *)
  wire [7:0] _01709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7947" *)
  wire [7:0] _01710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6687" *)
  wire [191:0] _01711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6677" *)
  wire [63:0] _01712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6697" *)
  wire [63:0] _01713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6667" *)
  wire [127:0] _01714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19945" *)
  wire [7:0] _01715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19955" *)
  wire [7:0] _01716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19965" *)
  wire [7:0] _01717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18815" *)
  wire [7:0] _01718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18825" *)
  wire [7:0] _01719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18835" *)
  wire [7:0] _01720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18845" *)
  wire [7:0] _01721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18855" *)
  wire [7:0] _01722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18865" *)
  wire [7:0] _01723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18875" *)
  wire [7:0] _01724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18885" *)
  wire [7:0] _01725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18705" *)
  wire [7:0] _01726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18895" *)
  wire [7:0] _01727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18905" *)
  wire [7:0] _01728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18915" *)
  wire [7:0] _01729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18925" *)
  wire [7:0] _01730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18935" *)
  wire [7:0] _01731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18945" *)
  wire [7:0] _01732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18955" *)
  wire [7:0] _01733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18965" *)
  wire [7:0] _01734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18975" *)
  wire [7:0] _01735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18985" *)
  wire [7:0] _01736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18715" *)
  wire [7:0] _01737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18995" *)
  wire [7:0] _01738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19005" *)
  wire [7:0] _01739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19015" *)
  wire [7:0] _01740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19025" *)
  wire [7:0] _01741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19035" *)
  wire [7:0] _01742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19045" *)
  wire [7:0] _01743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19055" *)
  wire [7:0] _01744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19065" *)
  wire [7:0] _01745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19075" *)
  wire [7:0] _01746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19085" *)
  wire [7:0] _01747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18725" *)
  wire [7:0] _01748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19095" *)
  wire [7:0] _01749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19105" *)
  wire [7:0] _01750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19115" *)
  wire [7:0] _01751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19125" *)
  wire [7:0] _01752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19135" *)
  wire [7:0] _01753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19145" *)
  wire [7:0] _01754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19155" *)
  wire [7:0] _01755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19165" *)
  wire [7:0] _01756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19175" *)
  wire [7:0] _01757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19185" *)
  wire [7:0] _01758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18735" *)
  wire [7:0] _01759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19195" *)
  wire [7:0] _01760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19205" *)
  wire [7:0] _01761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19215" *)
  wire [7:0] _01762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19225" *)
  wire [7:0] _01763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19235" *)
  wire [7:0] _01764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19245" *)
  wire [7:0] _01765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19255" *)
  wire [7:0] _01766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19265" *)
  wire [7:0] _01767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19275" *)
  wire [7:0] _01768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19285" *)
  wire [7:0] _01769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18745" *)
  wire [7:0] _01770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19295" *)
  wire [7:0] _01771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19305" *)
  wire [7:0] _01772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19315" *)
  wire [7:0] _01773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19325" *)
  wire [7:0] _01774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19335" *)
  wire [7:0] _01775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19345" *)
  wire [7:0] _01776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19355" *)
  wire [7:0] _01777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19365" *)
  wire [7:0] _01778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19375" *)
  wire [7:0] _01779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19385" *)
  wire [7:0] _01780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18755" *)
  wire [7:0] _01781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19395" *)
  wire [7:0] _01782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19405" *)
  wire [7:0] _01783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19415" *)
  wire [7:0] _01784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19425" *)
  wire [7:0] _01785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19435" *)
  wire [7:0] _01786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19445" *)
  wire [7:0] _01787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19455" *)
  wire [7:0] _01788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19465" *)
  wire [7:0] _01789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19475" *)
  wire [7:0] _01790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19485" *)
  wire [7:0] _01791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18765" *)
  wire [7:0] _01792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19495" *)
  wire [7:0] _01793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19505" *)
  wire [7:0] _01794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19515" *)
  wire [7:0] _01795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19525" *)
  wire [7:0] _01796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19535" *)
  wire [7:0] _01797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19545" *)
  wire [7:0] _01798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19555" *)
  wire [7:0] _01799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19565" *)
  wire [7:0] _01800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19575" *)
  wire [7:0] _01801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19585" *)
  wire [7:0] _01802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18775" *)
  wire [7:0] _01803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19595" *)
  wire [7:0] _01804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19605" *)
  wire [7:0] _01805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19615" *)
  wire [7:0] _01806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19625" *)
  wire [7:0] _01807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19635" *)
  wire [7:0] _01808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19645" *)
  wire [7:0] _01809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19655" *)
  wire [7:0] _01810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19665" *)
  wire [7:0] _01811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19675" *)
  wire [7:0] _01812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19685" *)
  wire [7:0] _01813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18785" *)
  wire [7:0] _01814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18695" *)
  wire [7:0] _01815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19695" *)
  wire [7:0] _01816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19705" *)
  wire [7:0] _01817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19715" *)
  wire [7:0] _01818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19725" *)
  wire [7:0] _01819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19735" *)
  wire [7:0] _01820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19745" *)
  wire [7:0] _01821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19755" *)
  wire [7:0] _01822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19765" *)
  wire [7:0] _01823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19775" *)
  wire [7:0] _01824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19785" *)
  wire [7:0] _01825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18795" *)
  wire [7:0] _01826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19795" *)
  wire [7:0] _01827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19805" *)
  wire [7:0] _01828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19815" *)
  wire [7:0] _01829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19825" *)
  wire [7:0] _01830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19835" *)
  wire [7:0] _01831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19845" *)
  wire [7:0] _01832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19855" *)
  wire [7:0] _01833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19865" *)
  wire [7:0] _01834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19875" *)
  wire [7:0] _01835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19885" *)
  wire [7:0] _01836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18805" *)
  wire [7:0] _01837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19895" *)
  wire [7:0] _01838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19905" *)
  wire [7:0] _01839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19915" *)
  wire [7:0] _01840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19925" *)
  wire [7:0] _01841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19935" *)
  wire [7:0] _01842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18685" *)
  wire [63:0] _01843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18675" *)
  wire [127:0] _01844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9293" *)
  wire [7:0] _01845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9303" *)
  wire [7:0] _01846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9313" *)
  wire [7:0] _01847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8163" *)
  wire [7:0] _01848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8173" *)
  wire [7:0] _01849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8183" *)
  wire [7:0] _01850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8193" *)
  wire [7:0] _01851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8203" *)
  wire [7:0] _01852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8213" *)
  wire [7:0] _01853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8223" *)
  wire [7:0] _01854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8233" *)
  wire [7:0] _01855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8053" *)
  wire [7:0] _01856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8243" *)
  wire [7:0] _01857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8253" *)
  wire [7:0] _01858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8263" *)
  wire [7:0] _01859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8273" *)
  wire [7:0] _01860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8283" *)
  wire [7:0] _01861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8293" *)
  wire [7:0] _01862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8303" *)
  wire [7:0] _01863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8313" *)
  wire [7:0] _01864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8323" *)
  wire [7:0] _01865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8333" *)
  wire [7:0] _01866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8063" *)
  wire [7:0] _01867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8343" *)
  wire [7:0] _01868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8353" *)
  wire [7:0] _01869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8363" *)
  wire [7:0] _01870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8373" *)
  wire [7:0] _01871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8383" *)
  wire [7:0] _01872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8393" *)
  wire [7:0] _01873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8403" *)
  wire [7:0] _01874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8413" *)
  wire [7:0] _01875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8423" *)
  wire [7:0] _01876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8433" *)
  wire [7:0] _01877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8073" *)
  wire [7:0] _01878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8443" *)
  wire [7:0] _01879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8453" *)
  wire [7:0] _01880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8463" *)
  wire [7:0] _01881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8473" *)
  wire [7:0] _01882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8483" *)
  wire [7:0] _01883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8493" *)
  wire [7:0] _01884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8503" *)
  wire [7:0] _01885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8513" *)
  wire [7:0] _01886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8523" *)
  wire [7:0] _01887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8533" *)
  wire [7:0] _01888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8083" *)
  wire [7:0] _01889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8543" *)
  wire [7:0] _01890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8553" *)
  wire [7:0] _01891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8563" *)
  wire [7:0] _01892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8573" *)
  wire [7:0] _01893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8583" *)
  wire [7:0] _01894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8593" *)
  wire [7:0] _01895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8603" *)
  wire [7:0] _01896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8613" *)
  wire [7:0] _01897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8623" *)
  wire [7:0] _01898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8633" *)
  wire [7:0] _01899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8093" *)
  wire [7:0] _01900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8643" *)
  wire [7:0] _01901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8653" *)
  wire [7:0] _01902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8663" *)
  wire [7:0] _01903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8673" *)
  wire [7:0] _01904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8683" *)
  wire [7:0] _01905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8693" *)
  wire [7:0] _01906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8703" *)
  wire [7:0] _01907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8713" *)
  wire [7:0] _01908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8723" *)
  wire [7:0] _01909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8733" *)
  wire [7:0] _01910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8103" *)
  wire [7:0] _01911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8743" *)
  wire [7:0] _01912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8753" *)
  wire [7:0] _01913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8763" *)
  wire [7:0] _01914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8773" *)
  wire [7:0] _01915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8783" *)
  wire [7:0] _01916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8793" *)
  wire [7:0] _01917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8803" *)
  wire [7:0] _01918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8813" *)
  wire [7:0] _01919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8823" *)
  wire [7:0] _01920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8833" *)
  wire [7:0] _01921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8113" *)
  wire [7:0] _01922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8843" *)
  wire [7:0] _01923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8853" *)
  wire [7:0] _01924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8863" *)
  wire [7:0] _01925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8873" *)
  wire [7:0] _01926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8883" *)
  wire [7:0] _01927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8893" *)
  wire [7:0] _01928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8903" *)
  wire [7:0] _01929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8913" *)
  wire [7:0] _01930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8923" *)
  wire [7:0] _01931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8933" *)
  wire [7:0] _01932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8123" *)
  wire [7:0] _01933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8943" *)
  wire [7:0] _01934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8953" *)
  wire [7:0] _01935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8963" *)
  wire [7:0] _01936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8973" *)
  wire [7:0] _01937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8983" *)
  wire [7:0] _01938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8993" *)
  wire [7:0] _01939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9003" *)
  wire [7:0] _01940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9013" *)
  wire [7:0] _01941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9023" *)
  wire [7:0] _01942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9033" *)
  wire [7:0] _01943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8133" *)
  wire [7:0] _01944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8043" *)
  wire [7:0] _01945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9043" *)
  wire [7:0] _01946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9053" *)
  wire [7:0] _01947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9063" *)
  wire [7:0] _01948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9073" *)
  wire [7:0] _01949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9083" *)
  wire [7:0] _01950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9093" *)
  wire [7:0] _01951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9103" *)
  wire [7:0] _01952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9113" *)
  wire [7:0] _01953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9123" *)
  wire [7:0] _01954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9133" *)
  wire [7:0] _01955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8143" *)
  wire [7:0] _01956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9143" *)
  wire [7:0] _01957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9153" *)
  wire [7:0] _01958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9163" *)
  wire [7:0] _01959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9173" *)
  wire [7:0] _01960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9183" *)
  wire [7:0] _01961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9193" *)
  wire [7:0] _01962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9203" *)
  wire [7:0] _01963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9213" *)
  wire [7:0] _01964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9223" *)
  wire [7:0] _01965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9233" *)
  wire [7:0] _01966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8153" *)
  wire [7:0] _01967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9243" *)
  wire [7:0] _01968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9253" *)
  wire [7:0] _01969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9263" *)
  wire [7:0] _01970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9273" *)
  wire [7:0] _01971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9283" *)
  wire [7:0] _01972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8023" *)
  wire [191:0] _01973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8013" *)
  wire [63:0] _01974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8033" *)
  wire [63:0] _01975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8003" *)
  wire [127:0] _01976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21269" *)
  wire [7:0] _01977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21279" *)
  wire [7:0] _01978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21289" *)
  wire [7:0] _01979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20139" *)
  wire [7:0] _01980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20149" *)
  wire [7:0] _01981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20159" *)
  wire [7:0] _01982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20169" *)
  wire [7:0] _01983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20179" *)
  wire [7:0] _01984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20189" *)
  wire [7:0] _01985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20199" *)
  wire [7:0] _01986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20209" *)
  wire [7:0] _01987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20029" *)
  wire [7:0] _01988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20219" *)
  wire [7:0] _01989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20229" *)
  wire [7:0] _01990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20239" *)
  wire [7:0] _01991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20249" *)
  wire [7:0] _01992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20259" *)
  wire [7:0] _01993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20269" *)
  wire [7:0] _01994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20279" *)
  wire [7:0] _01995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20289" *)
  wire [7:0] _01996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20299" *)
  wire [7:0] _01997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20309" *)
  wire [7:0] _01998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20039" *)
  wire [7:0] _01999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20319" *)
  wire [7:0] _02000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20329" *)
  wire [7:0] _02001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20339" *)
  wire [7:0] _02002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20349" *)
  wire [7:0] _02003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20359" *)
  wire [7:0] _02004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20369" *)
  wire [7:0] _02005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20379" *)
  wire [7:0] _02006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20389" *)
  wire [7:0] _02007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20399" *)
  wire [7:0] _02008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20409" *)
  wire [7:0] _02009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20049" *)
  wire [7:0] _02010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20419" *)
  wire [7:0] _02011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20429" *)
  wire [7:0] _02012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20439" *)
  wire [7:0] _02013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20449" *)
  wire [7:0] _02014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20459" *)
  wire [7:0] _02015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20469" *)
  wire [7:0] _02016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20479" *)
  wire [7:0] _02017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20489" *)
  wire [7:0] _02018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20499" *)
  wire [7:0] _02019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20509" *)
  wire [7:0] _02020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20059" *)
  wire [7:0] _02021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20519" *)
  wire [7:0] _02022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20529" *)
  wire [7:0] _02023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20539" *)
  wire [7:0] _02024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20549" *)
  wire [7:0] _02025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20559" *)
  wire [7:0] _02026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20569" *)
  wire [7:0] _02027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20579" *)
  wire [7:0] _02028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20589" *)
  wire [7:0] _02029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20599" *)
  wire [7:0] _02030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20609" *)
  wire [7:0] _02031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20069" *)
  wire [7:0] _02032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20619" *)
  wire [7:0] _02033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20629" *)
  wire [7:0] _02034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20639" *)
  wire [7:0] _02035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20649" *)
  wire [7:0] _02036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20659" *)
  wire [7:0] _02037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20669" *)
  wire [7:0] _02038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20679" *)
  wire [7:0] _02039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20689" *)
  wire [7:0] _02040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20699" *)
  wire [7:0] _02041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20709" *)
  wire [7:0] _02042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20079" *)
  wire [7:0] _02043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20719" *)
  wire [7:0] _02044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20729" *)
  wire [7:0] _02045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20739" *)
  wire [7:0] _02046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20749" *)
  wire [7:0] _02047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20759" *)
  wire [7:0] _02048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20769" *)
  wire [7:0] _02049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20779" *)
  wire [7:0] _02050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20789" *)
  wire [7:0] _02051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20799" *)
  wire [7:0] _02052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20809" *)
  wire [7:0] _02053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20089" *)
  wire [7:0] _02054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20819" *)
  wire [7:0] _02055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20829" *)
  wire [7:0] _02056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20839" *)
  wire [7:0] _02057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20849" *)
  wire [7:0] _02058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20859" *)
  wire [7:0] _02059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20869" *)
  wire [7:0] _02060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20879" *)
  wire [7:0] _02061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20889" *)
  wire [7:0] _02062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20899" *)
  wire [7:0] _02063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20909" *)
  wire [7:0] _02064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20099" *)
  wire [7:0] _02065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20919" *)
  wire [7:0] _02066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20929" *)
  wire [7:0] _02067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20939" *)
  wire [7:0] _02068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20949" *)
  wire [7:0] _02069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20959" *)
  wire [7:0] _02070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20969" *)
  wire [7:0] _02071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20979" *)
  wire [7:0] _02072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20989" *)
  wire [7:0] _02073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20999" *)
  wire [7:0] _02074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21009" *)
  wire [7:0] _02075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20109" *)
  wire [7:0] _02076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20019" *)
  wire [7:0] _02077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21019" *)
  wire [7:0] _02078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21029" *)
  wire [7:0] _02079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21039" *)
  wire [7:0] _02080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21049" *)
  wire [7:0] _02081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21059" *)
  wire [7:0] _02082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21069" *)
  wire [7:0] _02083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21079" *)
  wire [7:0] _02084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21089" *)
  wire [7:0] _02085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21099" *)
  wire [7:0] _02086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21109" *)
  wire [7:0] _02087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20119" *)
  wire [7:0] _02088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21119" *)
  wire [7:0] _02089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21129" *)
  wire [7:0] _02090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21139" *)
  wire [7:0] _02091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21149" *)
  wire [7:0] _02092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21159" *)
  wire [7:0] _02093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21169" *)
  wire [7:0] _02094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21179" *)
  wire [7:0] _02095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21189" *)
  wire [7:0] _02096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21199" *)
  wire [7:0] _02097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21209" *)
  wire [7:0] _02098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20129" *)
  wire [7:0] _02099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21219" *)
  wire [7:0] _02100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21229" *)
  wire [7:0] _02101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21239" *)
  wire [7:0] _02102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21249" *)
  wire [7:0] _02103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21259" *)
  wire [7:0] _02104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20009" *)
  wire [63:0] _02105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19999" *)
  wire [127:0] _02106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10629" *)
  wire [7:0] _02107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10639" *)
  wire [7:0] _02108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10649" *)
  wire [7:0] _02109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9499" *)
  wire [7:0] _02110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9509" *)
  wire [7:0] _02111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9519" *)
  wire [7:0] _02112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9529" *)
  wire [7:0] _02113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9539" *)
  wire [7:0] _02114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9549" *)
  wire [7:0] _02115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9559" *)
  wire [7:0] _02116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9569" *)
  wire [7:0] _02117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9389" *)
  wire [7:0] _02118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9579" *)
  wire [7:0] _02119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9589" *)
  wire [7:0] _02120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9599" *)
  wire [7:0] _02121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9609" *)
  wire [7:0] _02122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9619" *)
  wire [7:0] _02123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9629" *)
  wire [7:0] _02124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9639" *)
  wire [7:0] _02125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9649" *)
  wire [7:0] _02126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9659" *)
  wire [7:0] _02127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9669" *)
  wire [7:0] _02128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9399" *)
  wire [7:0] _02129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9679" *)
  wire [7:0] _02130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9689" *)
  wire [7:0] _02131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9699" *)
  wire [7:0] _02132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9709" *)
  wire [7:0] _02133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9719" *)
  wire [7:0] _02134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9729" *)
  wire [7:0] _02135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9739" *)
  wire [7:0] _02136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9749" *)
  wire [7:0] _02137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9759" *)
  wire [7:0] _02138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9769" *)
  wire [7:0] _02139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9409" *)
  wire [7:0] _02140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9779" *)
  wire [7:0] _02141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9789" *)
  wire [7:0] _02142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9799" *)
  wire [7:0] _02143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9809" *)
  wire [7:0] _02144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9819" *)
  wire [7:0] _02145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9829" *)
  wire [7:0] _02146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9839" *)
  wire [7:0] _02147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9849" *)
  wire [7:0] _02148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9859" *)
  wire [7:0] _02149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9869" *)
  wire [7:0] _02150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9419" *)
  wire [7:0] _02151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9879" *)
  wire [7:0] _02152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9889" *)
  wire [7:0] _02153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9899" *)
  wire [7:0] _02154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9909" *)
  wire [7:0] _02155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9919" *)
  wire [7:0] _02156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9929" *)
  wire [7:0] _02157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9939" *)
  wire [7:0] _02158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9949" *)
  wire [7:0] _02159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9959" *)
  wire [7:0] _02160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9969" *)
  wire [7:0] _02161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9429" *)
  wire [7:0] _02162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9979" *)
  wire [7:0] _02163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9989" *)
  wire [7:0] _02164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9999" *)
  wire [7:0] _02165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10009" *)
  wire [7:0] _02166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10019" *)
  wire [7:0] _02167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10029" *)
  wire [7:0] _02168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10039" *)
  wire [7:0] _02169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10049" *)
  wire [7:0] _02170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10059" *)
  wire [7:0] _02171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10069" *)
  wire [7:0] _02172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9439" *)
  wire [7:0] _02173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10079" *)
  wire [7:0] _02174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10089" *)
  wire [7:0] _02175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10099" *)
  wire [7:0] _02176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10109" *)
  wire [7:0] _02177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10119" *)
  wire [7:0] _02178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10129" *)
  wire [7:0] _02179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10139" *)
  wire [7:0] _02180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10149" *)
  wire [7:0] _02181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10159" *)
  wire [7:0] _02182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10169" *)
  wire [7:0] _02183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9449" *)
  wire [7:0] _02184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10179" *)
  wire [7:0] _02185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10189" *)
  wire [7:0] _02186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10199" *)
  wire [7:0] _02187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10209" *)
  wire [7:0] _02188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10219" *)
  wire [7:0] _02189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10229" *)
  wire [7:0] _02190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10239" *)
  wire [7:0] _02191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10249" *)
  wire [7:0] _02192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10259" *)
  wire [7:0] _02193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10269" *)
  wire [7:0] _02194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9459" *)
  wire [7:0] _02195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10279" *)
  wire [7:0] _02196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10289" *)
  wire [7:0] _02197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10299" *)
  wire [7:0] _02198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10309" *)
  wire [7:0] _02199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10319" *)
  wire [7:0] _02200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10329" *)
  wire [7:0] _02201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10339" *)
  wire [7:0] _02202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10349" *)
  wire [7:0] _02203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10359" *)
  wire [7:0] _02204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10369" *)
  wire [7:0] _02205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9469" *)
  wire [7:0] _02206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9379" *)
  wire [7:0] _02207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10379" *)
  wire [7:0] _02208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10389" *)
  wire [7:0] _02209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10399" *)
  wire [7:0] _02210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10409" *)
  wire [7:0] _02211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10419" *)
  wire [7:0] _02212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10429" *)
  wire [7:0] _02213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10439" *)
  wire [7:0] _02214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10449" *)
  wire [7:0] _02215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10459" *)
  wire [7:0] _02216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10469" *)
  wire [7:0] _02217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9479" *)
  wire [7:0] _02218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10479" *)
  wire [7:0] _02219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10489" *)
  wire [7:0] _02220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10499" *)
  wire [7:0] _02221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10509" *)
  wire [7:0] _02222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10519" *)
  wire [7:0] _02223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10529" *)
  wire [7:0] _02224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10539" *)
  wire [7:0] _02225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10549" *)
  wire [7:0] _02226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10559" *)
  wire [7:0] _02227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10569" *)
  wire [7:0] _02228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9489" *)
  wire [7:0] _02229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10579" *)
  wire [7:0] _02230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10589" *)
  wire [7:0] _02231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10599" *)
  wire [7:0] _02232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10609" *)
  wire [7:0] _02233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10619" *)
  wire [7:0] _02234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9359" *)
  wire [191:0] _02235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9349" *)
  wire [63:0] _02236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9369" *)
  wire [63:0] _02237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9339" *)
  wire [127:0] _02238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22593" *)
  wire [7:0] _02239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22603" *)
  wire [7:0] _02240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22613" *)
  wire [7:0] _02241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21463" *)
  wire [7:0] _02242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21473" *)
  wire [7:0] _02243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21483" *)
  wire [7:0] _02244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21493" *)
  wire [7:0] _02245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21503" *)
  wire [7:0] _02246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21513" *)
  wire [7:0] _02247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21523" *)
  wire [7:0] _02248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21533" *)
  wire [7:0] _02249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21353" *)
  wire [7:0] _02250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21543" *)
  wire [7:0] _02251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21553" *)
  wire [7:0] _02252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21563" *)
  wire [7:0] _02253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21573" *)
  wire [7:0] _02254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21583" *)
  wire [7:0] _02255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21593" *)
  wire [7:0] _02256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21603" *)
  wire [7:0] _02257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21613" *)
  wire [7:0] _02258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21623" *)
  wire [7:0] _02259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21633" *)
  wire [7:0] _02260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21363" *)
  wire [7:0] _02261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21643" *)
  wire [7:0] _02262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21653" *)
  wire [7:0] _02263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21663" *)
  wire [7:0] _02264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21673" *)
  wire [7:0] _02265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21683" *)
  wire [7:0] _02266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21693" *)
  wire [7:0] _02267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21703" *)
  wire [7:0] _02268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21713" *)
  wire [7:0] _02269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21723" *)
  wire [7:0] _02270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21733" *)
  wire [7:0] _02271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21373" *)
  wire [7:0] _02272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21743" *)
  wire [7:0] _02273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21753" *)
  wire [7:0] _02274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21763" *)
  wire [7:0] _02275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21773" *)
  wire [7:0] _02276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21783" *)
  wire [7:0] _02277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21793" *)
  wire [7:0] _02278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21803" *)
  wire [7:0] _02279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21813" *)
  wire [7:0] _02280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21823" *)
  wire [7:0] _02281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21833" *)
  wire [7:0] _02282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21383" *)
  wire [7:0] _02283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21843" *)
  wire [7:0] _02284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21853" *)
  wire [7:0] _02285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21863" *)
  wire [7:0] _02286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21873" *)
  wire [7:0] _02287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21883" *)
  wire [7:0] _02288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21893" *)
  wire [7:0] _02289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21903" *)
  wire [7:0] _02290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21913" *)
  wire [7:0] _02291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21923" *)
  wire [7:0] _02292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21933" *)
  wire [7:0] _02293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21393" *)
  wire [7:0] _02294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21943" *)
  wire [7:0] _02295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21953" *)
  wire [7:0] _02296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21963" *)
  wire [7:0] _02297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21973" *)
  wire [7:0] _02298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21983" *)
  wire [7:0] _02299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21993" *)
  wire [7:0] _02300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22003" *)
  wire [7:0] _02301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22013" *)
  wire [7:0] _02302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22023" *)
  wire [7:0] _02303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22033" *)
  wire [7:0] _02304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21403" *)
  wire [7:0] _02305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22043" *)
  wire [7:0] _02306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22053" *)
  wire [7:0] _02307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22063" *)
  wire [7:0] _02308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22073" *)
  wire [7:0] _02309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22083" *)
  wire [7:0] _02310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22093" *)
  wire [7:0] _02311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22103" *)
  wire [7:0] _02312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22113" *)
  wire [7:0] _02313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22123" *)
  wire [7:0] _02314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22133" *)
  wire [7:0] _02315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21413" *)
  wire [7:0] _02316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22143" *)
  wire [7:0] _02317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22153" *)
  wire [7:0] _02318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22163" *)
  wire [7:0] _02319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22173" *)
  wire [7:0] _02320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22183" *)
  wire [7:0] _02321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22193" *)
  wire [7:0] _02322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22203" *)
  wire [7:0] _02323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22213" *)
  wire [7:0] _02324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22223" *)
  wire [7:0] _02325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22233" *)
  wire [7:0] _02326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21423" *)
  wire [7:0] _02327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22243" *)
  wire [7:0] _02328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22253" *)
  wire [7:0] _02329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22263" *)
  wire [7:0] _02330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22273" *)
  wire [7:0] _02331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22283" *)
  wire [7:0] _02332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22293" *)
  wire [7:0] _02333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22303" *)
  wire [7:0] _02334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22313" *)
  wire [7:0] _02335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22323" *)
  wire [7:0] _02336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22333" *)
  wire [7:0] _02337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21433" *)
  wire [7:0] _02338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21343" *)
  wire [7:0] _02339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22343" *)
  wire [7:0] _02340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22353" *)
  wire [7:0] _02341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22363" *)
  wire [7:0] _02342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22373" *)
  wire [7:0] _02343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22383" *)
  wire [7:0] _02344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22393" *)
  wire [7:0] _02345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22403" *)
  wire [7:0] _02346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22413" *)
  wire [7:0] _02347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22423" *)
  wire [7:0] _02348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22433" *)
  wire [7:0] _02349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21443" *)
  wire [7:0] _02350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22443" *)
  wire [7:0] _02351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22453" *)
  wire [7:0] _02352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22463" *)
  wire [7:0] _02353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22473" *)
  wire [7:0] _02354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22483" *)
  wire [7:0] _02355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22493" *)
  wire [7:0] _02356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22503" *)
  wire [7:0] _02357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22513" *)
  wire [7:0] _02358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22523" *)
  wire [7:0] _02359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22533" *)
  wire [7:0] _02360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21453" *)
  wire [7:0] _02361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22543" *)
  wire [7:0] _02362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22553" *)
  wire [7:0] _02363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22563" *)
  wire [7:0] _02364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22573" *)
  wire [7:0] _02365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22583" *)
  wire [7:0] _02366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21333" *)
  wire [63:0] _02367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21323" *)
  wire [127:0] _02368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11965" *)
  wire [7:0] _02369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11975" *)
  wire [7:0] _02370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11985" *)
  wire [7:0] _02371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10835" *)
  wire [7:0] _02372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10845" *)
  wire [7:0] _02373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10855" *)
  wire [7:0] _02374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10865" *)
  wire [7:0] _02375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10875" *)
  wire [7:0] _02376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10885" *)
  wire [7:0] _02377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10895" *)
  wire [7:0] _02378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10905" *)
  wire [7:0] _02379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10725" *)
  wire [7:0] _02380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10915" *)
  wire [7:0] _02381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10925" *)
  wire [7:0] _02382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10935" *)
  wire [7:0] _02383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10945" *)
  wire [7:0] _02384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10955" *)
  wire [7:0] _02385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10965" *)
  wire [7:0] _02386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10975" *)
  wire [7:0] _02387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10985" *)
  wire [7:0] _02388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10995" *)
  wire [7:0] _02389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11005" *)
  wire [7:0] _02390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10735" *)
  wire [7:0] _02391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11015" *)
  wire [7:0] _02392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11025" *)
  wire [7:0] _02393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11035" *)
  wire [7:0] _02394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11045" *)
  wire [7:0] _02395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11055" *)
  wire [7:0] _02396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11065" *)
  wire [7:0] _02397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11075" *)
  wire [7:0] _02398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11085" *)
  wire [7:0] _02399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11095" *)
  wire [7:0] _02400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11105" *)
  wire [7:0] _02401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10745" *)
  wire [7:0] _02402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11115" *)
  wire [7:0] _02403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11125" *)
  wire [7:0] _02404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11135" *)
  wire [7:0] _02405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11145" *)
  wire [7:0] _02406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11155" *)
  wire [7:0] _02407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11165" *)
  wire [7:0] _02408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11175" *)
  wire [7:0] _02409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11185" *)
  wire [7:0] _02410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11195" *)
  wire [7:0] _02411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11205" *)
  wire [7:0] _02412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10755" *)
  wire [7:0] _02413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11215" *)
  wire [7:0] _02414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11225" *)
  wire [7:0] _02415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11235" *)
  wire [7:0] _02416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11245" *)
  wire [7:0] _02417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11255" *)
  wire [7:0] _02418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11265" *)
  wire [7:0] _02419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11275" *)
  wire [7:0] _02420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11285" *)
  wire [7:0] _02421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11295" *)
  wire [7:0] _02422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11305" *)
  wire [7:0] _02423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10765" *)
  wire [7:0] _02424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11315" *)
  wire [7:0] _02425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11325" *)
  wire [7:0] _02426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11335" *)
  wire [7:0] _02427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11345" *)
  wire [7:0] _02428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11355" *)
  wire [7:0] _02429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11365" *)
  wire [7:0] _02430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11375" *)
  wire [7:0] _02431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11385" *)
  wire [7:0] _02432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11395" *)
  wire [7:0] _02433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11405" *)
  wire [7:0] _02434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10775" *)
  wire [7:0] _02435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11415" *)
  wire [7:0] _02436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11425" *)
  wire [7:0] _02437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11435" *)
  wire [7:0] _02438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11445" *)
  wire [7:0] _02439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11455" *)
  wire [7:0] _02440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11465" *)
  wire [7:0] _02441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11475" *)
  wire [7:0] _02442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11485" *)
  wire [7:0] _02443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11495" *)
  wire [7:0] _02444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11505" *)
  wire [7:0] _02445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10785" *)
  wire [7:0] _02446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11515" *)
  wire [7:0] _02447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11525" *)
  wire [7:0] _02448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11535" *)
  wire [7:0] _02449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11545" *)
  wire [7:0] _02450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11555" *)
  wire [7:0] _02451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11565" *)
  wire [7:0] _02452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11575" *)
  wire [7:0] _02453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11585" *)
  wire [7:0] _02454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11595" *)
  wire [7:0] _02455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11605" *)
  wire [7:0] _02456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10795" *)
  wire [7:0] _02457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11615" *)
  wire [7:0] _02458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11625" *)
  wire [7:0] _02459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11635" *)
  wire [7:0] _02460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11645" *)
  wire [7:0] _02461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11655" *)
  wire [7:0] _02462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11665" *)
  wire [7:0] _02463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11675" *)
  wire [7:0] _02464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11685" *)
  wire [7:0] _02465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11695" *)
  wire [7:0] _02466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11705" *)
  wire [7:0] _02467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10805" *)
  wire [7:0] _02468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10715" *)
  wire [7:0] _02469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11715" *)
  wire [7:0] _02470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11725" *)
  wire [7:0] _02471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11735" *)
  wire [7:0] _02472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11745" *)
  wire [7:0] _02473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11755" *)
  wire [7:0] _02474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11765" *)
  wire [7:0] _02475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11775" *)
  wire [7:0] _02476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11785" *)
  wire [7:0] _02477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11795" *)
  wire [7:0] _02478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11805" *)
  wire [7:0] _02479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10815" *)
  wire [7:0] _02480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11815" *)
  wire [7:0] _02481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11825" *)
  wire [7:0] _02482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11835" *)
  wire [7:0] _02483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11845" *)
  wire [7:0] _02484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11855" *)
  wire [7:0] _02485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11865" *)
  wire [7:0] _02486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11875" *)
  wire [7:0] _02487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11885" *)
  wire [7:0] _02488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11895" *)
  wire [7:0] _02489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11905" *)
  wire [7:0] _02490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10825" *)
  wire [7:0] _02491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11915" *)
  wire [7:0] _02492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11925" *)
  wire [7:0] _02493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11935" *)
  wire [7:0] _02494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11945" *)
  wire [7:0] _02495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11955" *)
  wire [7:0] _02496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10695" *)
  wire [191:0] _02497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10685" *)
  wire [63:0] _02498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10705" *)
  wire [63:0] _02499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10675" *)
  wire [127:0] _02500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23917" *)
  wire [7:0] _02501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23927" *)
  wire [7:0] _02502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23937" *)
  wire [7:0] _02503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22787" *)
  wire [7:0] _02504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22797" *)
  wire [7:0] _02505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22807" *)
  wire [7:0] _02506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22817" *)
  wire [7:0] _02507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22827" *)
  wire [7:0] _02508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22837" *)
  wire [7:0] _02509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22847" *)
  wire [7:0] _02510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22857" *)
  wire [7:0] _02511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22677" *)
  wire [7:0] _02512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22867" *)
  wire [7:0] _02513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22877" *)
  wire [7:0] _02514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22887" *)
  wire [7:0] _02515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22897" *)
  wire [7:0] _02516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22907" *)
  wire [7:0] _02517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22917" *)
  wire [7:0] _02518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22927" *)
  wire [7:0] _02519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22937" *)
  wire [7:0] _02520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22947" *)
  wire [7:0] _02521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22957" *)
  wire [7:0] _02522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22687" *)
  wire [7:0] _02523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22967" *)
  wire [7:0] _02524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22977" *)
  wire [7:0] _02525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22987" *)
  wire [7:0] _02526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22997" *)
  wire [7:0] _02527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23007" *)
  wire [7:0] _02528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23017" *)
  wire [7:0] _02529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23027" *)
  wire [7:0] _02530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23037" *)
  wire [7:0] _02531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23047" *)
  wire [7:0] _02532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23057" *)
  wire [7:0] _02533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22697" *)
  wire [7:0] _02534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23067" *)
  wire [7:0] _02535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23077" *)
  wire [7:0] _02536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23087" *)
  wire [7:0] _02537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23097" *)
  wire [7:0] _02538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23107" *)
  wire [7:0] _02539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23117" *)
  wire [7:0] _02540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23127" *)
  wire [7:0] _02541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23137" *)
  wire [7:0] _02542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23147" *)
  wire [7:0] _02543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23157" *)
  wire [7:0] _02544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22707" *)
  wire [7:0] _02545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23167" *)
  wire [7:0] _02546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23177" *)
  wire [7:0] _02547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23187" *)
  wire [7:0] _02548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23197" *)
  wire [7:0] _02549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23207" *)
  wire [7:0] _02550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23217" *)
  wire [7:0] _02551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23227" *)
  wire [7:0] _02552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23237" *)
  wire [7:0] _02553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23247" *)
  wire [7:0] _02554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23257" *)
  wire [7:0] _02555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22717" *)
  wire [7:0] _02556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23267" *)
  wire [7:0] _02557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23277" *)
  wire [7:0] _02558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23287" *)
  wire [7:0] _02559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23297" *)
  wire [7:0] _02560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23307" *)
  wire [7:0] _02561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23317" *)
  wire [7:0] _02562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23327" *)
  wire [7:0] _02563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23337" *)
  wire [7:0] _02564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23347" *)
  wire [7:0] _02565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23357" *)
  wire [7:0] _02566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22727" *)
  wire [7:0] _02567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23367" *)
  wire [7:0] _02568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23377" *)
  wire [7:0] _02569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23387" *)
  wire [7:0] _02570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23397" *)
  wire [7:0] _02571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23407" *)
  wire [7:0] _02572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23417" *)
  wire [7:0] _02573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23427" *)
  wire [7:0] _02574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23437" *)
  wire [7:0] _02575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23447" *)
  wire [7:0] _02576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23457" *)
  wire [7:0] _02577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22737" *)
  wire [7:0] _02578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23467" *)
  wire [7:0] _02579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23477" *)
  wire [7:0] _02580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23487" *)
  wire [7:0] _02581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23497" *)
  wire [7:0] _02582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23507" *)
  wire [7:0] _02583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23517" *)
  wire [7:0] _02584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23527" *)
  wire [7:0] _02585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23537" *)
  wire [7:0] _02586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23547" *)
  wire [7:0] _02587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23557" *)
  wire [7:0] _02588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22747" *)
  wire [7:0] _02589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23567" *)
  wire [7:0] _02590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23577" *)
  wire [7:0] _02591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23587" *)
  wire [7:0] _02592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23597" *)
  wire [7:0] _02593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23607" *)
  wire [7:0] _02594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23617" *)
  wire [7:0] _02595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23627" *)
  wire [7:0] _02596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23637" *)
  wire [7:0] _02597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23647" *)
  wire [7:0] _02598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23657" *)
  wire [7:0] _02599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22757" *)
  wire [7:0] _02600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22667" *)
  wire [7:0] _02601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23667" *)
  wire [7:0] _02602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23677" *)
  wire [7:0] _02603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23687" *)
  wire [7:0] _02604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23697" *)
  wire [7:0] _02605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23707" *)
  wire [7:0] _02606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23717" *)
  wire [7:0] _02607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23727" *)
  wire [7:0] _02608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23737" *)
  wire [7:0] _02609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23747" *)
  wire [7:0] _02610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23757" *)
  wire [7:0] _02611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22767" *)
  wire [7:0] _02612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23767" *)
  wire [7:0] _02613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23777" *)
  wire [7:0] _02614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23787" *)
  wire [7:0] _02615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23797" *)
  wire [7:0] _02616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23807" *)
  wire [7:0] _02617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23817" *)
  wire [7:0] _02618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23827" *)
  wire [7:0] _02619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23837" *)
  wire [7:0] _02620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23847" *)
  wire [7:0] _02621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23857" *)
  wire [7:0] _02622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22777" *)
  wire [7:0] _02623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23867" *)
  wire [7:0] _02624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23877" *)
  wire [7:0] _02625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23887" *)
  wire [7:0] _02626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23897" *)
  wire [7:0] _02627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23907" *)
  wire [7:0] _02628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22657" *)
  wire [63:0] _02629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22647" *)
  wire [127:0] _02630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13301" *)
  wire [7:0] _02631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13311" *)
  wire [7:0] _02632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13321" *)
  wire [7:0] _02633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12171" *)
  wire [7:0] _02634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12181" *)
  wire [7:0] _02635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12191" *)
  wire [7:0] _02636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12201" *)
  wire [7:0] _02637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12211" *)
  wire [7:0] _02638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12221" *)
  wire [7:0] _02639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12231" *)
  wire [7:0] _02640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12241" *)
  wire [7:0] _02641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12061" *)
  wire [7:0] _02642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12251" *)
  wire [7:0] _02643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12261" *)
  wire [7:0] _02644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12271" *)
  wire [7:0] _02645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12281" *)
  wire [7:0] _02646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12291" *)
  wire [7:0] _02647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12301" *)
  wire [7:0] _02648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12311" *)
  wire [7:0] _02649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12321" *)
  wire [7:0] _02650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12331" *)
  wire [7:0] _02651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12341" *)
  wire [7:0] _02652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12071" *)
  wire [7:0] _02653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12351" *)
  wire [7:0] _02654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12361" *)
  wire [7:0] _02655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12371" *)
  wire [7:0] _02656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12381" *)
  wire [7:0] _02657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12391" *)
  wire [7:0] _02658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12401" *)
  wire [7:0] _02659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12411" *)
  wire [7:0] _02660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12421" *)
  wire [7:0] _02661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12431" *)
  wire [7:0] _02662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12441" *)
  wire [7:0] _02663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12081" *)
  wire [7:0] _02664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12451" *)
  wire [7:0] _02665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12461" *)
  wire [7:0] _02666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12471" *)
  wire [7:0] _02667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12481" *)
  wire [7:0] _02668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12491" *)
  wire [7:0] _02669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12501" *)
  wire [7:0] _02670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12511" *)
  wire [7:0] _02671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12521" *)
  wire [7:0] _02672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12531" *)
  wire [7:0] _02673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12541" *)
  wire [7:0] _02674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12091" *)
  wire [7:0] _02675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12551" *)
  wire [7:0] _02676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12561" *)
  wire [7:0] _02677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12571" *)
  wire [7:0] _02678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12581" *)
  wire [7:0] _02679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12591" *)
  wire [7:0] _02680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12601" *)
  wire [7:0] _02681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12611" *)
  wire [7:0] _02682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12621" *)
  wire [7:0] _02683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12631" *)
  wire [7:0] _02684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12641" *)
  wire [7:0] _02685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12101" *)
  wire [7:0] _02686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12651" *)
  wire [7:0] _02687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12661" *)
  wire [7:0] _02688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12671" *)
  wire [7:0] _02689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12681" *)
  wire [7:0] _02690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12691" *)
  wire [7:0] _02691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12701" *)
  wire [7:0] _02692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12711" *)
  wire [7:0] _02693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12721" *)
  wire [7:0] _02694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12731" *)
  wire [7:0] _02695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12741" *)
  wire [7:0] _02696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12111" *)
  wire [7:0] _02697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12751" *)
  wire [7:0] _02698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12761" *)
  wire [7:0] _02699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12771" *)
  wire [7:0] _02700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12781" *)
  wire [7:0] _02701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12791" *)
  wire [7:0] _02702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12801" *)
  wire [7:0] _02703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12811" *)
  wire [7:0] _02704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12821" *)
  wire [7:0] _02705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12831" *)
  wire [7:0] _02706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12841" *)
  wire [7:0] _02707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12121" *)
  wire [7:0] _02708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12851" *)
  wire [7:0] _02709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12861" *)
  wire [7:0] _02710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12871" *)
  wire [7:0] _02711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12881" *)
  wire [7:0] _02712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12891" *)
  wire [7:0] _02713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12901" *)
  wire [7:0] _02714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12911" *)
  wire [7:0] _02715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12921" *)
  wire [7:0] _02716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12931" *)
  wire [7:0] _02717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12941" *)
  wire [7:0] _02718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12131" *)
  wire [7:0] _02719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12951" *)
  wire [7:0] _02720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12961" *)
  wire [7:0] _02721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12971" *)
  wire [7:0] _02722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12981" *)
  wire [7:0] _02723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12991" *)
  wire [7:0] _02724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13001" *)
  wire [7:0] _02725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13011" *)
  wire [7:0] _02726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13021" *)
  wire [7:0] _02727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13031" *)
  wire [7:0] _02728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13041" *)
  wire [7:0] _02729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12141" *)
  wire [7:0] _02730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12051" *)
  wire [7:0] _02731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13051" *)
  wire [7:0] _02732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13061" *)
  wire [7:0] _02733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13071" *)
  wire [7:0] _02734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13081" *)
  wire [7:0] _02735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13091" *)
  wire [7:0] _02736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13101" *)
  wire [7:0] _02737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13111" *)
  wire [7:0] _02738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13121" *)
  wire [7:0] _02739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13131" *)
  wire [7:0] _02740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13141" *)
  wire [7:0] _02741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12151" *)
  wire [7:0] _02742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13151" *)
  wire [7:0] _02743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13161" *)
  wire [7:0] _02744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13171" *)
  wire [7:0] _02745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13181" *)
  wire [7:0] _02746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13191" *)
  wire [7:0] _02747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13201" *)
  wire [7:0] _02748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13211" *)
  wire [7:0] _02749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13221" *)
  wire [7:0] _02750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13231" *)
  wire [7:0] _02751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13241" *)
  wire [7:0] _02752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12161" *)
  wire [7:0] _02753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13251" *)
  wire [7:0] _02754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13261" *)
  wire [7:0] _02755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13271" *)
  wire [7:0] _02756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13281" *)
  wire [7:0] _02757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13291" *)
  wire [7:0] _02758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12031" *)
  wire [191:0] _02759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12021" *)
  wire [63:0] _02760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12041" *)
  wire [63:0] _02761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12011" *)
  wire [127:0] _02762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25241" *)
  wire [7:0] _02763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25251" *)
  wire [7:0] _02764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25261" *)
  wire [7:0] _02765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24111" *)
  wire [7:0] _02766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24121" *)
  wire [7:0] _02767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24131" *)
  wire [7:0] _02768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24141" *)
  wire [7:0] _02769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24151" *)
  wire [7:0] _02770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24161" *)
  wire [7:0] _02771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24171" *)
  wire [7:0] _02772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24181" *)
  wire [7:0] _02773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24001" *)
  wire [7:0] _02774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24191" *)
  wire [7:0] _02775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24201" *)
  wire [7:0] _02776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24211" *)
  wire [7:0] _02777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24221" *)
  wire [7:0] _02778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24231" *)
  wire [7:0] _02779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24241" *)
  wire [7:0] _02780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24251" *)
  wire [7:0] _02781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24261" *)
  wire [7:0] _02782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24271" *)
  wire [7:0] _02783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24281" *)
  wire [7:0] _02784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24011" *)
  wire [7:0] _02785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24291" *)
  wire [7:0] _02786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24301" *)
  wire [7:0] _02787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24311" *)
  wire [7:0] _02788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24321" *)
  wire [7:0] _02789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24331" *)
  wire [7:0] _02790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24341" *)
  wire [7:0] _02791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24351" *)
  wire [7:0] _02792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24361" *)
  wire [7:0] _02793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24371" *)
  wire [7:0] _02794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24381" *)
  wire [7:0] _02795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24021" *)
  wire [7:0] _02796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24391" *)
  wire [7:0] _02797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24401" *)
  wire [7:0] _02798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24411" *)
  wire [7:0] _02799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24421" *)
  wire [7:0] _02800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24431" *)
  wire [7:0] _02801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24441" *)
  wire [7:0] _02802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24451" *)
  wire [7:0] _02803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24461" *)
  wire [7:0] _02804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24471" *)
  wire [7:0] _02805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24481" *)
  wire [7:0] _02806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24031" *)
  wire [7:0] _02807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24491" *)
  wire [7:0] _02808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24501" *)
  wire [7:0] _02809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24511" *)
  wire [7:0] _02810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24521" *)
  wire [7:0] _02811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24531" *)
  wire [7:0] _02812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24541" *)
  wire [7:0] _02813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24551" *)
  wire [7:0] _02814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24561" *)
  wire [7:0] _02815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24571" *)
  wire [7:0] _02816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24581" *)
  wire [7:0] _02817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24041" *)
  wire [7:0] _02818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24591" *)
  wire [7:0] _02819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24601" *)
  wire [7:0] _02820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24611" *)
  wire [7:0] _02821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24621" *)
  wire [7:0] _02822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24631" *)
  wire [7:0] _02823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24641" *)
  wire [7:0] _02824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24651" *)
  wire [7:0] _02825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24661" *)
  wire [7:0] _02826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24671" *)
  wire [7:0] _02827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24681" *)
  wire [7:0] _02828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24051" *)
  wire [7:0] _02829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24691" *)
  wire [7:0] _02830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24701" *)
  wire [7:0] _02831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24711" *)
  wire [7:0] _02832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24721" *)
  wire [7:0] _02833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24731" *)
  wire [7:0] _02834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24741" *)
  wire [7:0] _02835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24751" *)
  wire [7:0] _02836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24761" *)
  wire [7:0] _02837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24771" *)
  wire [7:0] _02838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24781" *)
  wire [7:0] _02839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24061" *)
  wire [7:0] _02840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24791" *)
  wire [7:0] _02841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24801" *)
  wire [7:0] _02842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24811" *)
  wire [7:0] _02843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24821" *)
  wire [7:0] _02844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24831" *)
  wire [7:0] _02845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24841" *)
  wire [7:0] _02846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24851" *)
  wire [7:0] _02847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24861" *)
  wire [7:0] _02848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24871" *)
  wire [7:0] _02849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24881" *)
  wire [7:0] _02850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24071" *)
  wire [7:0] _02851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24891" *)
  wire [7:0] _02852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24901" *)
  wire [7:0] _02853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24911" *)
  wire [7:0] _02854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24921" *)
  wire [7:0] _02855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24931" *)
  wire [7:0] _02856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24941" *)
  wire [7:0] _02857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24951" *)
  wire [7:0] _02858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24961" *)
  wire [7:0] _02859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24971" *)
  wire [7:0] _02860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24981" *)
  wire [7:0] _02861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24081" *)
  wire [7:0] _02862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23991" *)
  wire [7:0] _02863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24991" *)
  wire [7:0] _02864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25001" *)
  wire [7:0] _02865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25011" *)
  wire [7:0] _02866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25021" *)
  wire [7:0] _02867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25031" *)
  wire [7:0] _02868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25041" *)
  wire [7:0] _02869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25051" *)
  wire [7:0] _02870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25061" *)
  wire [7:0] _02871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25071" *)
  wire [7:0] _02872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25081" *)
  wire [7:0] _02873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24091" *)
  wire [7:0] _02874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25091" *)
  wire [7:0] _02875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25101" *)
  wire [7:0] _02876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25111" *)
  wire [7:0] _02877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25121" *)
  wire [7:0] _02878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25131" *)
  wire [7:0] _02879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25141" *)
  wire [7:0] _02880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25151" *)
  wire [7:0] _02881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25161" *)
  wire [7:0] _02882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25171" *)
  wire [7:0] _02883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25181" *)
  wire [7:0] _02884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24101" *)
  wire [7:0] _02885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25191" *)
  wire [7:0] _02886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25201" *)
  wire [7:0] _02887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25211" *)
  wire [7:0] _02888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25221" *)
  wire [7:0] _02889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25231" *)
  wire [7:0] _02890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23981" *)
  wire [63:0] _02891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23971" *)
  wire [127:0] _02892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14637" *)
  wire [7:0] _02893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14647" *)
  wire [7:0] _02894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14657" *)
  wire [7:0] _02895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13507" *)
  wire [7:0] _02896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13517" *)
  wire [7:0] _02897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13527" *)
  wire [7:0] _02898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13537" *)
  wire [7:0] _02899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13547" *)
  wire [7:0] _02900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13557" *)
  wire [7:0] _02901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13567" *)
  wire [7:0] _02902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13577" *)
  wire [7:0] _02903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13397" *)
  wire [7:0] _02904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13587" *)
  wire [7:0] _02905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13597" *)
  wire [7:0] _02906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13607" *)
  wire [7:0] _02907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13617" *)
  wire [7:0] _02908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13627" *)
  wire [7:0] _02909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13637" *)
  wire [7:0] _02910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13647" *)
  wire [7:0] _02911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13657" *)
  wire [7:0] _02912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13667" *)
  wire [7:0] _02913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13677" *)
  wire [7:0] _02914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13407" *)
  wire [7:0] _02915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13687" *)
  wire [7:0] _02916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13697" *)
  wire [7:0] _02917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13707" *)
  wire [7:0] _02918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13717" *)
  wire [7:0] _02919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13727" *)
  wire [7:0] _02920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13737" *)
  wire [7:0] _02921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13747" *)
  wire [7:0] _02922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13757" *)
  wire [7:0] _02923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13767" *)
  wire [7:0] _02924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13777" *)
  wire [7:0] _02925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13417" *)
  wire [7:0] _02926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13787" *)
  wire [7:0] _02927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13797" *)
  wire [7:0] _02928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13807" *)
  wire [7:0] _02929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13817" *)
  wire [7:0] _02930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13827" *)
  wire [7:0] _02931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13837" *)
  wire [7:0] _02932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13847" *)
  wire [7:0] _02933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13857" *)
  wire [7:0] _02934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13867" *)
  wire [7:0] _02935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13877" *)
  wire [7:0] _02936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13427" *)
  wire [7:0] _02937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13887" *)
  wire [7:0] _02938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13897" *)
  wire [7:0] _02939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13907" *)
  wire [7:0] _02940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13917" *)
  wire [7:0] _02941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13927" *)
  wire [7:0] _02942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13937" *)
  wire [7:0] _02943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13947" *)
  wire [7:0] _02944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13957" *)
  wire [7:0] _02945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13967" *)
  wire [7:0] _02946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13977" *)
  wire [7:0] _02947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13437" *)
  wire [7:0] _02948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13987" *)
  wire [7:0] _02949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13997" *)
  wire [7:0] _02950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14007" *)
  wire [7:0] _02951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14017" *)
  wire [7:0] _02952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14027" *)
  wire [7:0] _02953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14037" *)
  wire [7:0] _02954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14047" *)
  wire [7:0] _02955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14057" *)
  wire [7:0] _02956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14067" *)
  wire [7:0] _02957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14077" *)
  wire [7:0] _02958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13447" *)
  wire [7:0] _02959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14087" *)
  wire [7:0] _02960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14097" *)
  wire [7:0] _02961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14107" *)
  wire [7:0] _02962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14117" *)
  wire [7:0] _02963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14127" *)
  wire [7:0] _02964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14137" *)
  wire [7:0] _02965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14147" *)
  wire [7:0] _02966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14157" *)
  wire [7:0] _02967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14167" *)
  wire [7:0] _02968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14177" *)
  wire [7:0] _02969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13457" *)
  wire [7:0] _02970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14187" *)
  wire [7:0] _02971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14197" *)
  wire [7:0] _02972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14207" *)
  wire [7:0] _02973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14217" *)
  wire [7:0] _02974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14227" *)
  wire [7:0] _02975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14237" *)
  wire [7:0] _02976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14247" *)
  wire [7:0] _02977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14257" *)
  wire [7:0] _02978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14267" *)
  wire [7:0] _02979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14277" *)
  wire [7:0] _02980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13467" *)
  wire [7:0] _02981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14287" *)
  wire [7:0] _02982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14297" *)
  wire [7:0] _02983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14307" *)
  wire [7:0] _02984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14317" *)
  wire [7:0] _02985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14327" *)
  wire [7:0] _02986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14337" *)
  wire [7:0] _02987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14347" *)
  wire [7:0] _02988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14357" *)
  wire [7:0] _02989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14367" *)
  wire [7:0] _02990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14377" *)
  wire [7:0] _02991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13477" *)
  wire [7:0] _02992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13387" *)
  wire [7:0] _02993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14387" *)
  wire [7:0] _02994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14397" *)
  wire [7:0] _02995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14407" *)
  wire [7:0] _02996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14417" *)
  wire [7:0] _02997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14427" *)
  wire [7:0] _02998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14437" *)
  wire [7:0] _02999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14447" *)
  wire [7:0] _03000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14457" *)
  wire [7:0] _03001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14467" *)
  wire [7:0] _03002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14477" *)
  wire [7:0] _03003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13487" *)
  wire [7:0] _03004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14487" *)
  wire [7:0] _03005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14497" *)
  wire [7:0] _03006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14507" *)
  wire [7:0] _03007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14517" *)
  wire [7:0] _03008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14527" *)
  wire [7:0] _03009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14537" *)
  wire [7:0] _03010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14547" *)
  wire [7:0] _03011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14557" *)
  wire [7:0] _03012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14567" *)
  wire [7:0] _03013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14577" *)
  wire [7:0] _03014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13497" *)
  wire [7:0] _03015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14587" *)
  wire [7:0] _03016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14597" *)
  wire [7:0] _03017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14607" *)
  wire [7:0] _03018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14617" *)
  wire [7:0] _03019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14627" *)
  wire [7:0] _03020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13367" *)
  wire [191:0] _03021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13357" *)
  wire [63:0] _03022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13377" *)
  wire [63:0] _03023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13347" *)
  wire [127:0] _03024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26565" *)
  wire [7:0] _03025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26575" *)
  wire [7:0] _03026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26585" *)
  wire [7:0] _03027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25435" *)
  wire [7:0] _03028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25445" *)
  wire [7:0] _03029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25455" *)
  wire [7:0] _03030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25465" *)
  wire [7:0] _03031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25475" *)
  wire [7:0] _03032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25485" *)
  wire [7:0] _03033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25495" *)
  wire [7:0] _03034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25505" *)
  wire [7:0] _03035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25325" *)
  wire [7:0] _03036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25515" *)
  wire [7:0] _03037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25525" *)
  wire [7:0] _03038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25535" *)
  wire [7:0] _03039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25545" *)
  wire [7:0] _03040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25555" *)
  wire [7:0] _03041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25565" *)
  wire [7:0] _03042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25575" *)
  wire [7:0] _03043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25585" *)
  wire [7:0] _03044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25595" *)
  wire [7:0] _03045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25605" *)
  wire [7:0] _03046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25335" *)
  wire [7:0] _03047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25615" *)
  wire [7:0] _03048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25625" *)
  wire [7:0] _03049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25635" *)
  wire [7:0] _03050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25645" *)
  wire [7:0] _03051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25655" *)
  wire [7:0] _03052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25665" *)
  wire [7:0] _03053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25675" *)
  wire [7:0] _03054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25685" *)
  wire [7:0] _03055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25695" *)
  wire [7:0] _03056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25705" *)
  wire [7:0] _03057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25345" *)
  wire [7:0] _03058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25715" *)
  wire [7:0] _03059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25725" *)
  wire [7:0] _03060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25735" *)
  wire [7:0] _03061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25745" *)
  wire [7:0] _03062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25755" *)
  wire [7:0] _03063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25765" *)
  wire [7:0] _03064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25775" *)
  wire [7:0] _03065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25785" *)
  wire [7:0] _03066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25795" *)
  wire [7:0] _03067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25805" *)
  wire [7:0] _03068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25355" *)
  wire [7:0] _03069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25815" *)
  wire [7:0] _03070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25825" *)
  wire [7:0] _03071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25835" *)
  wire [7:0] _03072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25845" *)
  wire [7:0] _03073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25855" *)
  wire [7:0] _03074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25865" *)
  wire [7:0] _03075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25875" *)
  wire [7:0] _03076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25885" *)
  wire [7:0] _03077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25895" *)
  wire [7:0] _03078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25905" *)
  wire [7:0] _03079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25365" *)
  wire [7:0] _03080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25915" *)
  wire [7:0] _03081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25925" *)
  wire [7:0] _03082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25935" *)
  wire [7:0] _03083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25945" *)
  wire [7:0] _03084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25955" *)
  wire [7:0] _03085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25965" *)
  wire [7:0] _03086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25975" *)
  wire [7:0] _03087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25985" *)
  wire [7:0] _03088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25995" *)
  wire [7:0] _03089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26005" *)
  wire [7:0] _03090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25375" *)
  wire [7:0] _03091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26015" *)
  wire [7:0] _03092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26025" *)
  wire [7:0] _03093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26035" *)
  wire [7:0] _03094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26045" *)
  wire [7:0] _03095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26055" *)
  wire [7:0] _03096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26065" *)
  wire [7:0] _03097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26075" *)
  wire [7:0] _03098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26085" *)
  wire [7:0] _03099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26095" *)
  wire [7:0] _03100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26105" *)
  wire [7:0] _03101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25385" *)
  wire [7:0] _03102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26115" *)
  wire [7:0] _03103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26125" *)
  wire [7:0] _03104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26135" *)
  wire [7:0] _03105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26145" *)
  wire [7:0] _03106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26155" *)
  wire [7:0] _03107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26165" *)
  wire [7:0] _03108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26175" *)
  wire [7:0] _03109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26185" *)
  wire [7:0] _03110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26195" *)
  wire [7:0] _03111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26205" *)
  wire [7:0] _03112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25395" *)
  wire [7:0] _03113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26215" *)
  wire [7:0] _03114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26225" *)
  wire [7:0] _03115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26235" *)
  wire [7:0] _03116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26245" *)
  wire [7:0] _03117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26255" *)
  wire [7:0] _03118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26265" *)
  wire [7:0] _03119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26275" *)
  wire [7:0] _03120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26285" *)
  wire [7:0] _03121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26295" *)
  wire [7:0] _03122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26305" *)
  wire [7:0] _03123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25405" *)
  wire [7:0] _03124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25315" *)
  wire [7:0] _03125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26315" *)
  wire [7:0] _03126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26325" *)
  wire [7:0] _03127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26335" *)
  wire [7:0] _03128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26345" *)
  wire [7:0] _03129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26355" *)
  wire [7:0] _03130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26365" *)
  wire [7:0] _03131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26375" *)
  wire [7:0] _03132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26385" *)
  wire [7:0] _03133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26395" *)
  wire [7:0] _03134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26405" *)
  wire [7:0] _03135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25415" *)
  wire [7:0] _03136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26415" *)
  wire [7:0] _03137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26425" *)
  wire [7:0] _03138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26435" *)
  wire [7:0] _03139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26445" *)
  wire [7:0] _03140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26455" *)
  wire [7:0] _03141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26465" *)
  wire [7:0] _03142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26475" *)
  wire [7:0] _03143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26485" *)
  wire [7:0] _03144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26495" *)
  wire [7:0] _03145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26505" *)
  wire [7:0] _03146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25425" *)
  wire [7:0] _03147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26515" *)
  wire [7:0] _03148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26525" *)
  wire [7:0] _03149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26535" *)
  wire [7:0] _03150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26545" *)
  wire [7:0] _03151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26555" *)
  wire [7:0] _03152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25305" *)
  wire [63:0] _03153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25295" *)
  wire [127:0] _03154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15973" *)
  wire [7:0] _03155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15983" *)
  wire [7:0] _03156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15993" *)
  wire [7:0] _03157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14843" *)
  wire [7:0] _03158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14853" *)
  wire [7:0] _03159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14863" *)
  wire [7:0] _03160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14873" *)
  wire [7:0] _03161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14883" *)
  wire [7:0] _03162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14893" *)
  wire [7:0] _03163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14903" *)
  wire [7:0] _03164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14913" *)
  wire [7:0] _03165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14733" *)
  wire [7:0] _03166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14923" *)
  wire [7:0] _03167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14933" *)
  wire [7:0] _03168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14943" *)
  wire [7:0] _03169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14953" *)
  wire [7:0] _03170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14963" *)
  wire [7:0] _03171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14973" *)
  wire [7:0] _03172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14983" *)
  wire [7:0] _03173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14993" *)
  wire [7:0] _03174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15003" *)
  wire [7:0] _03175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15013" *)
  wire [7:0] _03176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14743" *)
  wire [7:0] _03177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15023" *)
  wire [7:0] _03178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15033" *)
  wire [7:0] _03179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15043" *)
  wire [7:0] _03180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15053" *)
  wire [7:0] _03181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15063" *)
  wire [7:0] _03182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15073" *)
  wire [7:0] _03183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15083" *)
  wire [7:0] _03184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15093" *)
  wire [7:0] _03185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15103" *)
  wire [7:0] _03186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15113" *)
  wire [7:0] _03187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14753" *)
  wire [7:0] _03188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15123" *)
  wire [7:0] _03189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15133" *)
  wire [7:0] _03190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15143" *)
  wire [7:0] _03191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15153" *)
  wire [7:0] _03192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15163" *)
  wire [7:0] _03193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15173" *)
  wire [7:0] _03194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15183" *)
  wire [7:0] _03195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15193" *)
  wire [7:0] _03196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15203" *)
  wire [7:0] _03197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15213" *)
  wire [7:0] _03198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14763" *)
  wire [7:0] _03199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15223" *)
  wire [7:0] _03200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15233" *)
  wire [7:0] _03201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15243" *)
  wire [7:0] _03202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15253" *)
  wire [7:0] _03203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15263" *)
  wire [7:0] _03204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15273" *)
  wire [7:0] _03205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15283" *)
  wire [7:0] _03206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15293" *)
  wire [7:0] _03207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15303" *)
  wire [7:0] _03208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15313" *)
  wire [7:0] _03209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14773" *)
  wire [7:0] _03210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15323" *)
  wire [7:0] _03211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15333" *)
  wire [7:0] _03212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15343" *)
  wire [7:0] _03213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15353" *)
  wire [7:0] _03214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15363" *)
  wire [7:0] _03215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15373" *)
  wire [7:0] _03216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15383" *)
  wire [7:0] _03217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15393" *)
  wire [7:0] _03218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15403" *)
  wire [7:0] _03219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15413" *)
  wire [7:0] _03220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14783" *)
  wire [7:0] _03221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15423" *)
  wire [7:0] _03222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15433" *)
  wire [7:0] _03223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15443" *)
  wire [7:0] _03224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15453" *)
  wire [7:0] _03225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15463" *)
  wire [7:0] _03226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15473" *)
  wire [7:0] _03227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15483" *)
  wire [7:0] _03228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15493" *)
  wire [7:0] _03229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15503" *)
  wire [7:0] _03230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15513" *)
  wire [7:0] _03231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14793" *)
  wire [7:0] _03232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15523" *)
  wire [7:0] _03233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15533" *)
  wire [7:0] _03234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15543" *)
  wire [7:0] _03235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15553" *)
  wire [7:0] _03236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15563" *)
  wire [7:0] _03237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15573" *)
  wire [7:0] _03238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15583" *)
  wire [7:0] _03239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15593" *)
  wire [7:0] _03240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15603" *)
  wire [7:0] _03241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15613" *)
  wire [7:0] _03242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14803" *)
  wire [7:0] _03243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15623" *)
  wire [7:0] _03244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15633" *)
  wire [7:0] _03245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15643" *)
  wire [7:0] _03246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15653" *)
  wire [7:0] _03247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15663" *)
  wire [7:0] _03248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15673" *)
  wire [7:0] _03249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15683" *)
  wire [7:0] _03250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15693" *)
  wire [7:0] _03251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15703" *)
  wire [7:0] _03252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15713" *)
  wire [7:0] _03253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14813" *)
  wire [7:0] _03254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14723" *)
  wire [7:0] _03255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15723" *)
  wire [7:0] _03256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15733" *)
  wire [7:0] _03257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15743" *)
  wire [7:0] _03258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15753" *)
  wire [7:0] _03259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15763" *)
  wire [7:0] _03260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15773" *)
  wire [7:0] _03261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15783" *)
  wire [7:0] _03262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15793" *)
  wire [7:0] _03263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15803" *)
  wire [7:0] _03264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15813" *)
  wire [7:0] _03265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14823" *)
  wire [7:0] _03266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15823" *)
  wire [7:0] _03267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15833" *)
  wire [7:0] _03268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15843" *)
  wire [7:0] _03269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15853" *)
  wire [7:0] _03270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15863" *)
  wire [7:0] _03271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15873" *)
  wire [7:0] _03272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15883" *)
  wire [7:0] _03273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15893" *)
  wire [7:0] _03274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15903" *)
  wire [7:0] _03275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15913" *)
  wire [7:0] _03276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14833" *)
  wire [7:0] _03277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15923" *)
  wire [7:0] _03278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15933" *)
  wire [7:0] _03279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15943" *)
  wire [7:0] _03280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15953" *)
  wire [7:0] _03281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15963" *)
  wire [7:0] _03282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14703" *)
  wire [191:0] _03283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14693" *)
  wire [63:0] _03284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14713" *)
  wire [63:0] _03285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14683" *)
  wire [127:0] _03286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5282" *)
  wire [7:0] _03287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5292" *)
  wire [7:0] _03288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5302" *)
  wire [7:0] _03289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4152" *)
  wire [7:0] _03290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4162" *)
  wire [7:0] _03291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4172" *)
  wire [7:0] _03292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4182" *)
  wire [7:0] _03293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4192" *)
  wire [7:0] _03294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4202" *)
  wire [7:0] _03295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4212" *)
  wire [7:0] _03296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4222" *)
  wire [7:0] _03297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4042" *)
  wire [7:0] _03298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4232" *)
  wire [7:0] _03299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4242" *)
  wire [7:0] _03300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4252" *)
  wire [7:0] _03301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4262" *)
  wire [7:0] _03302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4272" *)
  wire [7:0] _03303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4282" *)
  wire [7:0] _03304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4292" *)
  wire [7:0] _03305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4302" *)
  wire [7:0] _03306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4312" *)
  wire [7:0] _03307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4322" *)
  wire [7:0] _03308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4052" *)
  wire [7:0] _03309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4332" *)
  wire [7:0] _03310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4342" *)
  wire [7:0] _03311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4352" *)
  wire [7:0] _03312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4362" *)
  wire [7:0] _03313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4372" *)
  wire [7:0] _03314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4382" *)
  wire [7:0] _03315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4392" *)
  wire [7:0] _03316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4402" *)
  wire [7:0] _03317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4412" *)
  wire [7:0] _03318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4422" *)
  wire [7:0] _03319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4062" *)
  wire [7:0] _03320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4432" *)
  wire [7:0] _03321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4442" *)
  wire [7:0] _03322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4452" *)
  wire [7:0] _03323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4462" *)
  wire [7:0] _03324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4472" *)
  wire [7:0] _03325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4482" *)
  wire [7:0] _03326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4492" *)
  wire [7:0] _03327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4502" *)
  wire [7:0] _03328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4512" *)
  wire [7:0] _03329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4522" *)
  wire [7:0] _03330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4072" *)
  wire [7:0] _03331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4532" *)
  wire [7:0] _03332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4542" *)
  wire [7:0] _03333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4552" *)
  wire [7:0] _03334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4562" *)
  wire [7:0] _03335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4572" *)
  wire [7:0] _03336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4582" *)
  wire [7:0] _03337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4592" *)
  wire [7:0] _03338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4602" *)
  wire [7:0] _03339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4612" *)
  wire [7:0] _03340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4622" *)
  wire [7:0] _03341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4082" *)
  wire [7:0] _03342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4632" *)
  wire [7:0] _03343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4642" *)
  wire [7:0] _03344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4652" *)
  wire [7:0] _03345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4662" *)
  wire [7:0] _03346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4672" *)
  wire [7:0] _03347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4682" *)
  wire [7:0] _03348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4692" *)
  wire [7:0] _03349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4702" *)
  wire [7:0] _03350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4712" *)
  wire [7:0] _03351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4722" *)
  wire [7:0] _03352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4092" *)
  wire [7:0] _03353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4732" *)
  wire [7:0] _03354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4742" *)
  wire [7:0] _03355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4752" *)
  wire [7:0] _03356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4762" *)
  wire [7:0] _03357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4772" *)
  wire [7:0] _03358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4782" *)
  wire [7:0] _03359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4792" *)
  wire [7:0] _03360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4802" *)
  wire [7:0] _03361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4812" *)
  wire [7:0] _03362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4822" *)
  wire [7:0] _03363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4102" *)
  wire [7:0] _03364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4832" *)
  wire [7:0] _03365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4842" *)
  wire [7:0] _03366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4852" *)
  wire [7:0] _03367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4862" *)
  wire [7:0] _03368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4872" *)
  wire [7:0] _03369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4882" *)
  wire [7:0] _03370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4892" *)
  wire [7:0] _03371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4902" *)
  wire [7:0] _03372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4912" *)
  wire [7:0] _03373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4922" *)
  wire [7:0] _03374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4112" *)
  wire [7:0] _03375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4932" *)
  wire [7:0] _03376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4942" *)
  wire [7:0] _03377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4952" *)
  wire [7:0] _03378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4962" *)
  wire [7:0] _03379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4972" *)
  wire [7:0] _03380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4982" *)
  wire [7:0] _03381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4992" *)
  wire [7:0] _03382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5002" *)
  wire [7:0] _03383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5012" *)
  wire [7:0] _03384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5022" *)
  wire [7:0] _03385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4122" *)
  wire [7:0] _03386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4032" *)
  wire [7:0] _03387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5032" *)
  wire [7:0] _03388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5042" *)
  wire [7:0] _03389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5052" *)
  wire [7:0] _03390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5062" *)
  wire [7:0] _03391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5072" *)
  wire [7:0] _03392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5082" *)
  wire [7:0] _03393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5092" *)
  wire [7:0] _03394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5102" *)
  wire [7:0] _03395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5112" *)
  wire [7:0] _03396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5122" *)
  wire [7:0] _03397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4132" *)
  wire [7:0] _03398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5132" *)
  wire [7:0] _03399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5142" *)
  wire [7:0] _03400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5152" *)
  wire [7:0] _03401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5162" *)
  wire [7:0] _03402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5172" *)
  wire [7:0] _03403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5182" *)
  wire [7:0] _03404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5192" *)
  wire [7:0] _03405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5202" *)
  wire [7:0] _03406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5212" *)
  wire [7:0] _03407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5222" *)
  wire [7:0] _03408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4142" *)
  wire [7:0] _03409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5232" *)
  wire [7:0] _03410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5242" *)
  wire [7:0] _03411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5252" *)
  wire [7:0] _03412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5262" *)
  wire [7:0] _03413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5272" *)
  wire [7:0] _03414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4012" *)
  wire [191:0] _03415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4002" *)
  wire [63:0] _03416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4022" *)
  wire [63:0] _03417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3992" *)
  wire [127:0] _03418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10000" *)
  wire _03419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10010" *)
  wire _03420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10020" *)
  wire _03421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10030" *)
  wire _03422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10040" *)
  wire _03423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10050" *)
  wire _03424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10060" *)
  wire _03425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10070" *)
  wire _03426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10080" *)
  wire _03427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10090" *)
  wire _03428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10100" *)
  wire _03429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10110" *)
  wire _03430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10120" *)
  wire _03431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10130" *)
  wire _03432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10140" *)
  wire _03433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10150" *)
  wire _03434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10160" *)
  wire _03435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10170" *)
  wire _03436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10180" *)
  wire _03437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10190" *)
  wire _03438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10200" *)
  wire _03439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10210" *)
  wire _03440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10220" *)
  wire _03441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10230" *)
  wire _03442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10240" *)
  wire _03443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10250" *)
  wire _03444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10260" *)
  wire _03445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10270" *)
  wire _03446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10280" *)
  wire _03447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10290" *)
  wire _03448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10300" *)
  wire _03449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10310" *)
  wire _03450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10320" *)
  wire _03451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10330" *)
  wire _03452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10340" *)
  wire _03453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10350" *)
  wire _03454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10360" *)
  wire _03455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10370" *)
  wire _03456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10380" *)
  wire _03457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10390" *)
  wire _03458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10400" *)
  wire _03459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10410" *)
  wire _03460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10420" *)
  wire _03461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10430" *)
  wire _03462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10440" *)
  wire _03463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10450" *)
  wire _03464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10460" *)
  wire _03465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10470" *)
  wire _03466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10480" *)
  wire _03467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10490" *)
  wire _03468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10500" *)
  wire _03469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10510" *)
  wire _03470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10520" *)
  wire _03471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10530" *)
  wire _03472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10540" *)
  wire _03473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10550" *)
  wire _03474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10560" *)
  wire _03475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10570" *)
  wire _03476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10580" *)
  wire _03477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10590" *)
  wire _03478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10600" *)
  wire _03479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10610" *)
  wire _03480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10620" *)
  wire _03481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10630" *)
  wire _03482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10640" *)
  wire _03483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10650" *)
  wire _03484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10686" *)
  wire _03485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10716" *)
  wire _03486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10726" *)
  wire _03487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10736" *)
  wire _03488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10746" *)
  wire _03489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10756" *)
  wire _03490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10766" *)
  wire _03491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10776" *)
  wire _03492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10786" *)
  wire _03493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10796" *)
  wire _03494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10806" *)
  wire _03495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10816" *)
  wire _03496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10826" *)
  wire _03497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10836" *)
  wire _03498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10846" *)
  wire _03499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10856" *)
  wire _03500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10866" *)
  wire _03501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10876" *)
  wire _03502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10886" *)
  wire _03503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10896" *)
  wire _03504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10906" *)
  wire _03505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10916" *)
  wire _03506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10926" *)
  wire _03507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10936" *)
  wire _03508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10946" *)
  wire _03509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10956" *)
  wire _03510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10966" *)
  wire _03511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10976" *)
  wire _03512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10986" *)
  wire _03513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10996" *)
  wire _03514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11006" *)
  wire _03515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11016" *)
  wire _03516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11026" *)
  wire _03517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11036" *)
  wire _03518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11046" *)
  wire _03519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11056" *)
  wire _03520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11066" *)
  wire _03521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11076" *)
  wire _03522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11086" *)
  wire _03523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11096" *)
  wire _03524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11106" *)
  wire _03525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11116" *)
  wire _03526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11126" *)
  wire _03527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11136" *)
  wire _03528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11146" *)
  wire _03529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11156" *)
  wire _03530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11166" *)
  wire _03531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11176" *)
  wire _03532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11186" *)
  wire _03533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11196" *)
  wire _03534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11206" *)
  wire _03535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11216" *)
  wire _03536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11226" *)
  wire _03537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11236" *)
  wire _03538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11246" *)
  wire _03539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11256" *)
  wire _03540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11266" *)
  wire _03541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11276" *)
  wire _03542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11286" *)
  wire _03543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11296" *)
  wire _03544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11306" *)
  wire _03545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11316" *)
  wire _03546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11326" *)
  wire _03547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11336" *)
  wire _03548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11346" *)
  wire _03549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11356" *)
  wire _03550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11366" *)
  wire _03551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11376" *)
  wire _03552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11386" *)
  wire _03553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11396" *)
  wire _03554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11406" *)
  wire _03555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11416" *)
  wire _03556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11426" *)
  wire _03557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11436" *)
  wire _03558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11446" *)
  wire _03559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11456" *)
  wire _03560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11466" *)
  wire _03561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11476" *)
  wire _03562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11486" *)
  wire _03563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11496" *)
  wire _03564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11506" *)
  wire _03565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11516" *)
  wire _03566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11526" *)
  wire _03567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11536" *)
  wire _03568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11546" *)
  wire _03569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11556" *)
  wire _03570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11566" *)
  wire _03571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11576" *)
  wire _03572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11586" *)
  wire _03573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11596" *)
  wire _03574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11606" *)
  wire _03575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11616" *)
  wire _03576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11626" *)
  wire _03577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11636" *)
  wire _03578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11646" *)
  wire _03579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11656" *)
  wire _03580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11666" *)
  wire _03581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11676" *)
  wire _03582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11686" *)
  wire _03583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11696" *)
  wire _03584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11706" *)
  wire _03585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11716" *)
  wire _03586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11726" *)
  wire _03587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11736" *)
  wire _03588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11746" *)
  wire _03589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11756" *)
  wire _03590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11766" *)
  wire _03591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11776" *)
  wire _03592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11786" *)
  wire _03593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11796" *)
  wire _03594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11806" *)
  wire _03595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11816" *)
  wire _03596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11826" *)
  wire _03597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11836" *)
  wire _03598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11846" *)
  wire _03599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11856" *)
  wire _03600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11866" *)
  wire _03601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11876" *)
  wire _03602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11886" *)
  wire _03603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11896" *)
  wire _03604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11906" *)
  wire _03605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11916" *)
  wire _03606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11926" *)
  wire _03607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11936" *)
  wire _03608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11946" *)
  wire _03609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11956" *)
  wire _03610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11966" *)
  wire _03611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11976" *)
  wire _03612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11986" *)
  wire _03613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12022" *)
  wire _03614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12052" *)
  wire _03615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12062" *)
  wire _03616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12072" *)
  wire _03617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12082" *)
  wire _03618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12092" *)
  wire _03619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12102" *)
  wire _03620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12112" *)
  wire _03621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12122" *)
  wire _03622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12132" *)
  wire _03623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12142" *)
  wire _03624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12152" *)
  wire _03625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12162" *)
  wire _03626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12172" *)
  wire _03627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12182" *)
  wire _03628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12192" *)
  wire _03629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12202" *)
  wire _03630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12212" *)
  wire _03631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12222" *)
  wire _03632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12232" *)
  wire _03633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12242" *)
  wire _03634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12252" *)
  wire _03635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12262" *)
  wire _03636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12272" *)
  wire _03637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12282" *)
  wire _03638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12292" *)
  wire _03639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12302" *)
  wire _03640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12312" *)
  wire _03641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12322" *)
  wire _03642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12332" *)
  wire _03643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12342" *)
  wire _03644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12352" *)
  wire _03645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12362" *)
  wire _03646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12372" *)
  wire _03647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12382" *)
  wire _03648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12392" *)
  wire _03649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12402" *)
  wire _03650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12412" *)
  wire _03651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12422" *)
  wire _03652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12432" *)
  wire _03653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12442" *)
  wire _03654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12452" *)
  wire _03655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12462" *)
  wire _03656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12472" *)
  wire _03657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12482" *)
  wire _03658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12492" *)
  wire _03659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12502" *)
  wire _03660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12512" *)
  wire _03661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12522" *)
  wire _03662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12532" *)
  wire _03663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12542" *)
  wire _03664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12552" *)
  wire _03665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12562" *)
  wire _03666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12572" *)
  wire _03667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12582" *)
  wire _03668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12592" *)
  wire _03669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12602" *)
  wire _03670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12612" *)
  wire _03671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12622" *)
  wire _03672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12632" *)
  wire _03673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12642" *)
  wire _03674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12652" *)
  wire _03675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12662" *)
  wire _03676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12672" *)
  wire _03677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12682" *)
  wire _03678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12692" *)
  wire _03679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12702" *)
  wire _03680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12712" *)
  wire _03681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12722" *)
  wire _03682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12732" *)
  wire _03683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12742" *)
  wire _03684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12752" *)
  wire _03685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12762" *)
  wire _03686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12772" *)
  wire _03687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12782" *)
  wire _03688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12792" *)
  wire _03689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12802" *)
  wire _03690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12812" *)
  wire _03691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12822" *)
  wire _03692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12832" *)
  wire _03693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12842" *)
  wire _03694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12852" *)
  wire _03695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12862" *)
  wire _03696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12872" *)
  wire _03697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12882" *)
  wire _03698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12892" *)
  wire _03699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12902" *)
  wire _03700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12912" *)
  wire _03701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12922" *)
  wire _03702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12932" *)
  wire _03703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12942" *)
  wire _03704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12952" *)
  wire _03705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12962" *)
  wire _03706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12972" *)
  wire _03707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12982" *)
  wire _03708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12992" *)
  wire _03709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13002" *)
  wire _03710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13012" *)
  wire _03711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13022" *)
  wire _03712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13032" *)
  wire _03713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13042" *)
  wire _03714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13052" *)
  wire _03715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13062" *)
  wire _03716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13072" *)
  wire _03717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13082" *)
  wire _03718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13092" *)
  wire _03719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13102" *)
  wire _03720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13112" *)
  wire _03721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13122" *)
  wire _03722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13132" *)
  wire _03723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13142" *)
  wire _03724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13152" *)
  wire _03725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13162" *)
  wire _03726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13172" *)
  wire _03727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13182" *)
  wire _03728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13192" *)
  wire _03729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13202" *)
  wire _03730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13212" *)
  wire _03731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13222" *)
  wire _03732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13232" *)
  wire _03733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13242" *)
  wire _03734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13252" *)
  wire _03735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13262" *)
  wire _03736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13272" *)
  wire _03737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13282" *)
  wire _03738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13292" *)
  wire _03739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13302" *)
  wire _03740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13312" *)
  wire _03741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13322" *)
  wire _03742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13358" *)
  wire _03743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13388" *)
  wire _03744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13398" *)
  wire _03745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13408" *)
  wire _03746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13418" *)
  wire _03747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13428" *)
  wire _03748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13438" *)
  wire _03749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13448" *)
  wire _03750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13458" *)
  wire _03751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13468" *)
  wire _03752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13478" *)
  wire _03753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13488" *)
  wire _03754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13498" *)
  wire _03755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13508" *)
  wire _03756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13518" *)
  wire _03757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13528" *)
  wire _03758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13538" *)
  wire _03759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13548" *)
  wire _03760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13558" *)
  wire _03761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13568" *)
  wire _03762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13578" *)
  wire _03763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13588" *)
  wire _03764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13598" *)
  wire _03765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13608" *)
  wire _03766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13618" *)
  wire _03767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13628" *)
  wire _03768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13638" *)
  wire _03769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13648" *)
  wire _03770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13658" *)
  wire _03771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13668" *)
  wire _03772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13678" *)
  wire _03773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13688" *)
  wire _03774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13698" *)
  wire _03775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13708" *)
  wire _03776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13718" *)
  wire _03777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13728" *)
  wire _03778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13738" *)
  wire _03779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13748" *)
  wire _03780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13758" *)
  wire _03781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13768" *)
  wire _03782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13778" *)
  wire _03783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13788" *)
  wire _03784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13798" *)
  wire _03785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13808" *)
  wire _03786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13818" *)
  wire _03787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13828" *)
  wire _03788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13838" *)
  wire _03789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13848" *)
  wire _03790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13858" *)
  wire _03791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13868" *)
  wire _03792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13878" *)
  wire _03793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13888" *)
  wire _03794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13898" *)
  wire _03795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13908" *)
  wire _03796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13918" *)
  wire _03797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13928" *)
  wire _03798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13938" *)
  wire _03799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13948" *)
  wire _03800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13958" *)
  wire _03801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13968" *)
  wire _03802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13978" *)
  wire _03803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13988" *)
  wire _03804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13998" *)
  wire _03805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14008" *)
  wire _03806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14018" *)
  wire _03807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14028" *)
  wire _03808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14038" *)
  wire _03809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14048" *)
  wire _03810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14058" *)
  wire _03811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14068" *)
  wire _03812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14078" *)
  wire _03813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14088" *)
  wire _03814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14098" *)
  wire _03815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14108" *)
  wire _03816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14118" *)
  wire _03817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14128" *)
  wire _03818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14138" *)
  wire _03819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14148" *)
  wire _03820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14158" *)
  wire _03821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14168" *)
  wire _03822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14178" *)
  wire _03823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14188" *)
  wire _03824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14198" *)
  wire _03825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14208" *)
  wire _03826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14218" *)
  wire _03827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14228" *)
  wire _03828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14238" *)
  wire _03829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14248" *)
  wire _03830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14258" *)
  wire _03831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14268" *)
  wire _03832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14278" *)
  wire _03833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14288" *)
  wire _03834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14298" *)
  wire _03835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14308" *)
  wire _03836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14318" *)
  wire _03837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14328" *)
  wire _03838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14338" *)
  wire _03839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14348" *)
  wire _03840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14358" *)
  wire _03841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14368" *)
  wire _03842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14378" *)
  wire _03843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14388" *)
  wire _03844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14398" *)
  wire _03845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14408" *)
  wire _03846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14418" *)
  wire _03847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14428" *)
  wire _03848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14438" *)
  wire _03849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14448" *)
  wire _03850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14458" *)
  wire _03851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14468" *)
  wire _03852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14478" *)
  wire _03853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14488" *)
  wire _03854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14498" *)
  wire _03855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14508" *)
  wire _03856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14518" *)
  wire _03857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14528" *)
  wire _03858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14538" *)
  wire _03859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14548" *)
  wire _03860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14558" *)
  wire _03861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14568" *)
  wire _03862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14578" *)
  wire _03863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14588" *)
  wire _03864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14598" *)
  wire _03865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14608" *)
  wire _03866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14618" *)
  wire _03867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14628" *)
  wire _03868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14638" *)
  wire _03869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14648" *)
  wire _03870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14658" *)
  wire _03871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14694" *)
  wire _03872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14724" *)
  wire _03873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14734" *)
  wire _03874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14744" *)
  wire _03875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14754" *)
  wire _03876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14764" *)
  wire _03877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14774" *)
  wire _03878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14784" *)
  wire _03879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14794" *)
  wire _03880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14804" *)
  wire _03881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14814" *)
  wire _03882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14824" *)
  wire _03883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14834" *)
  wire _03884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14844" *)
  wire _03885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14854" *)
  wire _03886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14864" *)
  wire _03887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14874" *)
  wire _03888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14884" *)
  wire _03889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14894" *)
  wire _03890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14904" *)
  wire _03891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14914" *)
  wire _03892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14924" *)
  wire _03893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14934" *)
  wire _03894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14944" *)
  wire _03895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14954" *)
  wire _03896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14964" *)
  wire _03897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14974" *)
  wire _03898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14984" *)
  wire _03899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14994" *)
  wire _03900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15004" *)
  wire _03901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15014" *)
  wire _03902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15024" *)
  wire _03903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15034" *)
  wire _03904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15044" *)
  wire _03905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15054" *)
  wire _03906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15064" *)
  wire _03907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15074" *)
  wire _03908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15084" *)
  wire _03909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15094" *)
  wire _03910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15104" *)
  wire _03911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15114" *)
  wire _03912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15124" *)
  wire _03913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15134" *)
  wire _03914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15144" *)
  wire _03915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15154" *)
  wire _03916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15164" *)
  wire _03917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15174" *)
  wire _03918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15184" *)
  wire _03919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15194" *)
  wire _03920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15204" *)
  wire _03921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15214" *)
  wire _03922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15224" *)
  wire _03923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15234" *)
  wire _03924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15244" *)
  wire _03925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15254" *)
  wire _03926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15264" *)
  wire _03927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15274" *)
  wire _03928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15284" *)
  wire _03929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15294" *)
  wire _03930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15304" *)
  wire _03931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15314" *)
  wire _03932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15324" *)
  wire _03933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15334" *)
  wire _03934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15344" *)
  wire _03935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15354" *)
  wire _03936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15364" *)
  wire _03937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15374" *)
  wire _03938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15384" *)
  wire _03939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15394" *)
  wire _03940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15404" *)
  wire _03941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15414" *)
  wire _03942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15424" *)
  wire _03943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15434" *)
  wire _03944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15444" *)
  wire _03945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15454" *)
  wire _03946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15464" *)
  wire _03947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15474" *)
  wire _03948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15484" *)
  wire _03949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15494" *)
  wire _03950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15504" *)
  wire _03951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15514" *)
  wire _03952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15524" *)
  wire _03953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15534" *)
  wire _03954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15544" *)
  wire _03955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15554" *)
  wire _03956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15564" *)
  wire _03957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15574" *)
  wire _03958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15584" *)
  wire _03959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15594" *)
  wire _03960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15604" *)
  wire _03961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15614" *)
  wire _03962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15624" *)
  wire _03963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15634" *)
  wire _03964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15644" *)
  wire _03965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15654" *)
  wire _03966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15664" *)
  wire _03967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15674" *)
  wire _03968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15684" *)
  wire _03969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15694" *)
  wire _03970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15704" *)
  wire _03971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15714" *)
  wire _03972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15724" *)
  wire _03973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15734" *)
  wire _03974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15744" *)
  wire _03975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15754" *)
  wire _03976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15764" *)
  wire _03977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15774" *)
  wire _03978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15784" *)
  wire _03979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15794" *)
  wire _03980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15804" *)
  wire _03981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15814" *)
  wire _03982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15824" *)
  wire _03983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15834" *)
  wire _03984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15844" *)
  wire _03985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15854" *)
  wire _03986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15864" *)
  wire _03987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15874" *)
  wire _03988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15884" *)
  wire _03989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15894" *)
  wire _03990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15904" *)
  wire _03991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15914" *)
  wire _03992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15924" *)
  wire _03993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15934" *)
  wire _03994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15944" *)
  wire _03995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15954" *)
  wire _03996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15964" *)
  wire _03997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15974" *)
  wire _03998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15984" *)
  wire _03999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15994" *)
  wire _04000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16028" *)
  wire _04001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16038" *)
  wire _04002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16049" *)
  wire [7:0] _04003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16059" *)
  wire [7:0] _04004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16069" *)
  wire [7:0] _04005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16079" *)
  wire [7:0] _04006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16089" *)
  wire [7:0] _04007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16099" *)
  wire [7:0] _04008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16109" *)
  wire [7:0] _04009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16119" *)
  wire [7:0] _04010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16129" *)
  wire [7:0] _04011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16139" *)
  wire [7:0] _04012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16149" *)
  wire [7:0] _04013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16159" *)
  wire [7:0] _04014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16169" *)
  wire [7:0] _04015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16179" *)
  wire [7:0] _04016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16189" *)
  wire [7:0] _04017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16199" *)
  wire [7:0] _04018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16209" *)
  wire [7:0] _04019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16219" *)
  wire [7:0] _04020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16229" *)
  wire [7:0] _04021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16239" *)
  wire [7:0] _04022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16249" *)
  wire [7:0] _04023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16259" *)
  wire [7:0] _04024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16269" *)
  wire [7:0] _04025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16279" *)
  wire [7:0] _04026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16289" *)
  wire [7:0] _04027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16299" *)
  wire [7:0] _04028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16309" *)
  wire [7:0] _04029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16319" *)
  wire [7:0] _04030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16329" *)
  wire [7:0] _04031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16339" *)
  wire [7:0] _04032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16349" *)
  wire [7:0] _04033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16359" *)
  wire [7:0] _04034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16369" *)
  wire [7:0] _04035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16379" *)
  wire [7:0] _04036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16389" *)
  wire [7:0] _04037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16399" *)
  wire [7:0] _04038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16409" *)
  wire [7:0] _04039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16419" *)
  wire [7:0] _04040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16429" *)
  wire [7:0] _04041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16439" *)
  wire [7:0] _04042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16449" *)
  wire [7:0] _04043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16459" *)
  wire [7:0] _04044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16469" *)
  wire [7:0] _04045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16479" *)
  wire [7:0] _04046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16489" *)
  wire [7:0] _04047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16499" *)
  wire [7:0] _04048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16509" *)
  wire [7:0] _04049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16519" *)
  wire [7:0] _04050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16529" *)
  wire [7:0] _04051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16539" *)
  wire [7:0] _04052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16549" *)
  wire [7:0] _04053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16559" *)
  wire [7:0] _04054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16569" *)
  wire [7:0] _04055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16579" *)
  wire [7:0] _04056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16589" *)
  wire [7:0] _04057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16599" *)
  wire [7:0] _04058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16609" *)
  wire [7:0] _04059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16619" *)
  wire [7:0] _04060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16629" *)
  wire [7:0] _04061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16639" *)
  wire [7:0] _04062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16649" *)
  wire [7:0] _04063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16659" *)
  wire [7:0] _04064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16669" *)
  wire [7:0] _04065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16679" *)
  wire [7:0] _04066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16689" *)
  wire [7:0] _04067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16699" *)
  wire [7:0] _04068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16709" *)
  wire [7:0] _04069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16719" *)
  wire [7:0] _04070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16729" *)
  wire [7:0] _04071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16739" *)
  wire [7:0] _04072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16749" *)
  wire [7:0] _04073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16759" *)
  wire [7:0] _04074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16769" *)
  wire [7:0] _04075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16779" *)
  wire [7:0] _04076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16789" *)
  wire [7:0] _04077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16799" *)
  wire [7:0] _04078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16809" *)
  wire [7:0] _04079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16819" *)
  wire [7:0] _04080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16829" *)
  wire [7:0] _04081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16839" *)
  wire [7:0] _04082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16849" *)
  wire [7:0] _04083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16859" *)
  wire [7:0] _04084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16869" *)
  wire [7:0] _04085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16879" *)
  wire [7:0] _04086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16889" *)
  wire [7:0] _04087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16899" *)
  wire [7:0] _04088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16909" *)
  wire [7:0] _04089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16919" *)
  wire [7:0] _04090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16929" *)
  wire [7:0] _04091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16939" *)
  wire [7:0] _04092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16949" *)
  wire [7:0] _04093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16959" *)
  wire [7:0] _04094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16969" *)
  wire [7:0] _04095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16979" *)
  wire [7:0] _04096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16989" *)
  wire [7:0] _04097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16999" *)
  wire [7:0] _04098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17009" *)
  wire [7:0] _04099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17019" *)
  wire [7:0] _04100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17029" *)
  wire [7:0] _04101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17039" *)
  wire [7:0] _04102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17049" *)
  wire [7:0] _04103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17059" *)
  wire [7:0] _04104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17069" *)
  wire [7:0] _04105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17079" *)
  wire [7:0] _04106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17089" *)
  wire [7:0] _04107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17099" *)
  wire [7:0] _04108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17109" *)
  wire [7:0] _04109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17119" *)
  wire [7:0] _04110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17129" *)
  wire [7:0] _04111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17139" *)
  wire [7:0] _04112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17149" *)
  wire [7:0] _04113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17159" *)
  wire [7:0] _04114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17169" *)
  wire [7:0] _04115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17179" *)
  wire [7:0] _04116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17189" *)
  wire [7:0] _04117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17199" *)
  wire [7:0] _04118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17209" *)
  wire [7:0] _04119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17219" *)
  wire [7:0] _04120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17229" *)
  wire [7:0] _04121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17239" *)
  wire [7:0] _04122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17249" *)
  wire [7:0] _04123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17259" *)
  wire [7:0] _04124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17269" *)
  wire [7:0] _04125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17279" *)
  wire [7:0] _04126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17289" *)
  wire [7:0] _04127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17299" *)
  wire [7:0] _04128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17309" *)
  wire [7:0] _04129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17319" *)
  wire [7:0] _04130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17352" *)
  wire _04131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17362" *)
  wire _04132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17373" *)
  wire [7:0] _04133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17383" *)
  wire [7:0] _04134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17393" *)
  wire [7:0] _04135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17403" *)
  wire [7:0] _04136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17413" *)
  wire [7:0] _04137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17423" *)
  wire [7:0] _04138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17433" *)
  wire [7:0] _04139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17443" *)
  wire [7:0] _04140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17453" *)
  wire [7:0] _04141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17463" *)
  wire [7:0] _04142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17473" *)
  wire [7:0] _04143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17483" *)
  wire [7:0] _04144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17493" *)
  wire [7:0] _04145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17503" *)
  wire [7:0] _04146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17513" *)
  wire [7:0] _04147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17523" *)
  wire [7:0] _04148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17533" *)
  wire [7:0] _04149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17543" *)
  wire [7:0] _04150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17553" *)
  wire [7:0] _04151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17563" *)
  wire [7:0] _04152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17573" *)
  wire [7:0] _04153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17583" *)
  wire [7:0] _04154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17593" *)
  wire [7:0] _04155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17603" *)
  wire [7:0] _04156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17613" *)
  wire [7:0] _04157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17623" *)
  wire [7:0] _04158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17633" *)
  wire [7:0] _04159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17643" *)
  wire [7:0] _04160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17653" *)
  wire [7:0] _04161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17663" *)
  wire [7:0] _04162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17673" *)
  wire [7:0] _04163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17683" *)
  wire [7:0] _04164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17693" *)
  wire [7:0] _04165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17703" *)
  wire [7:0] _04166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17713" *)
  wire [7:0] _04167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17723" *)
  wire [7:0] _04168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17733" *)
  wire [7:0] _04169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17743" *)
  wire [7:0] _04170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17753" *)
  wire [7:0] _04171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17763" *)
  wire [7:0] _04172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17773" *)
  wire [7:0] _04173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17783" *)
  wire [7:0] _04174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17793" *)
  wire [7:0] _04175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17803" *)
  wire [7:0] _04176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17813" *)
  wire [7:0] _04177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17823" *)
  wire [7:0] _04178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17833" *)
  wire [7:0] _04179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17843" *)
  wire [7:0] _04180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17853" *)
  wire [7:0] _04181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17863" *)
  wire [7:0] _04182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17873" *)
  wire [7:0] _04183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17883" *)
  wire [7:0] _04184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17893" *)
  wire [7:0] _04185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17903" *)
  wire [7:0] _04186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17913" *)
  wire [7:0] _04187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17923" *)
  wire [7:0] _04188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17933" *)
  wire [7:0] _04189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17943" *)
  wire [7:0] _04190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17953" *)
  wire [7:0] _04191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17963" *)
  wire [7:0] _04192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17973" *)
  wire [7:0] _04193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17983" *)
  wire [7:0] _04194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17993" *)
  wire [7:0] _04195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18003" *)
  wire [7:0] _04196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18013" *)
  wire [7:0] _04197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18023" *)
  wire [7:0] _04198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18033" *)
  wire [7:0] _04199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18043" *)
  wire [7:0] _04200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18053" *)
  wire [7:0] _04201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18063" *)
  wire [7:0] _04202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18073" *)
  wire [7:0] _04203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18083" *)
  wire [7:0] _04204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18093" *)
  wire [7:0] _04205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18103" *)
  wire [7:0] _04206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18113" *)
  wire [7:0] _04207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18123" *)
  wire [7:0] _04208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18133" *)
  wire [7:0] _04209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18143" *)
  wire [7:0] _04210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18153" *)
  wire [7:0] _04211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18163" *)
  wire [7:0] _04212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18173" *)
  wire [7:0] _04213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18183" *)
  wire [7:0] _04214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18193" *)
  wire [7:0] _04215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18203" *)
  wire [7:0] _04216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18213" *)
  wire [7:0] _04217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18223" *)
  wire [7:0] _04218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18233" *)
  wire [7:0] _04219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18243" *)
  wire [7:0] _04220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18253" *)
  wire [7:0] _04221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18263" *)
  wire [7:0] _04222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18273" *)
  wire [7:0] _04223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18283" *)
  wire [7:0] _04224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18293" *)
  wire [7:0] _04225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18303" *)
  wire [7:0] _04226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18313" *)
  wire [7:0] _04227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18323" *)
  wire [7:0] _04228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18333" *)
  wire [7:0] _04229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18343" *)
  wire [7:0] _04230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18353" *)
  wire [7:0] _04231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18363" *)
  wire [7:0] _04232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18373" *)
  wire [7:0] _04233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18383" *)
  wire [7:0] _04234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18393" *)
  wire [7:0] _04235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18403" *)
  wire [7:0] _04236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18413" *)
  wire [7:0] _04237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18423" *)
  wire [7:0] _04238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18433" *)
  wire [7:0] _04239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18443" *)
  wire [7:0] _04240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18453" *)
  wire [7:0] _04241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18463" *)
  wire [7:0] _04242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18473" *)
  wire [7:0] _04243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18483" *)
  wire [7:0] _04244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18493" *)
  wire [7:0] _04245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18503" *)
  wire [7:0] _04246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18513" *)
  wire [7:0] _04247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18523" *)
  wire [7:0] _04248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18533" *)
  wire [7:0] _04249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18543" *)
  wire [7:0] _04250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18553" *)
  wire [7:0] _04251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18563" *)
  wire [7:0] _04252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18573" *)
  wire [7:0] _04253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18583" *)
  wire [7:0] _04254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18593" *)
  wire [7:0] _04255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18603" *)
  wire [7:0] _04256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18613" *)
  wire [7:0] _04257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18623" *)
  wire [7:0] _04258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18633" *)
  wire [7:0] _04259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18643" *)
  wire [7:0] _04260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18676" *)
  wire _04261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18686" *)
  wire _04262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18697" *)
  wire [7:0] _04263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18707" *)
  wire [7:0] _04264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18717" *)
  wire [7:0] _04265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18727" *)
  wire [7:0] _04266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18737" *)
  wire [7:0] _04267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18747" *)
  wire [7:0] _04268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18757" *)
  wire [7:0] _04269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18767" *)
  wire [7:0] _04270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18777" *)
  wire [7:0] _04271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18787" *)
  wire [7:0] _04272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18797" *)
  wire [7:0] _04273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18807" *)
  wire [7:0] _04274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18817" *)
  wire [7:0] _04275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18827" *)
  wire [7:0] _04276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18837" *)
  wire [7:0] _04277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18847" *)
  wire [7:0] _04278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18857" *)
  wire [7:0] _04279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18867" *)
  wire [7:0] _04280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18877" *)
  wire [7:0] _04281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18887" *)
  wire [7:0] _04282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18897" *)
  wire [7:0] _04283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18907" *)
  wire [7:0] _04284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18917" *)
  wire [7:0] _04285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18927" *)
  wire [7:0] _04286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18937" *)
  wire [7:0] _04287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18947" *)
  wire [7:0] _04288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18957" *)
  wire [7:0] _04289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18967" *)
  wire [7:0] _04290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18977" *)
  wire [7:0] _04291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18987" *)
  wire [7:0] _04292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18997" *)
  wire [7:0] _04293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19007" *)
  wire [7:0] _04294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19017" *)
  wire [7:0] _04295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19027" *)
  wire [7:0] _04296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19037" *)
  wire [7:0] _04297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19047" *)
  wire [7:0] _04298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19057" *)
  wire [7:0] _04299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19067" *)
  wire [7:0] _04300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19077" *)
  wire [7:0] _04301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19087" *)
  wire [7:0] _04302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19097" *)
  wire [7:0] _04303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19107" *)
  wire [7:0] _04304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19117" *)
  wire [7:0] _04305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19127" *)
  wire [7:0] _04306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19137" *)
  wire [7:0] _04307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19147" *)
  wire [7:0] _04308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19157" *)
  wire [7:0] _04309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19167" *)
  wire [7:0] _04310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19177" *)
  wire [7:0] _04311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19187" *)
  wire [7:0] _04312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19197" *)
  wire [7:0] _04313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19207" *)
  wire [7:0] _04314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19217" *)
  wire [7:0] _04315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19227" *)
  wire [7:0] _04316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19237" *)
  wire [7:0] _04317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19247" *)
  wire [7:0] _04318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19257" *)
  wire [7:0] _04319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19267" *)
  wire [7:0] _04320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19277" *)
  wire [7:0] _04321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19287" *)
  wire [7:0] _04322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19297" *)
  wire [7:0] _04323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19307" *)
  wire [7:0] _04324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19317" *)
  wire [7:0] _04325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19327" *)
  wire [7:0] _04326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19337" *)
  wire [7:0] _04327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19347" *)
  wire [7:0] _04328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19357" *)
  wire [7:0] _04329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19367" *)
  wire [7:0] _04330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19377" *)
  wire [7:0] _04331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19387" *)
  wire [7:0] _04332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19397" *)
  wire [7:0] _04333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19407" *)
  wire [7:0] _04334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19417" *)
  wire [7:0] _04335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19427" *)
  wire [7:0] _04336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19437" *)
  wire [7:0] _04337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19447" *)
  wire [7:0] _04338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19457" *)
  wire [7:0] _04339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19467" *)
  wire [7:0] _04340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19477" *)
  wire [7:0] _04341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19487" *)
  wire [7:0] _04342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19497" *)
  wire [7:0] _04343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19507" *)
  wire [7:0] _04344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19517" *)
  wire [7:0] _04345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19527" *)
  wire [7:0] _04346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19537" *)
  wire [7:0] _04347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19547" *)
  wire [7:0] _04348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19557" *)
  wire [7:0] _04349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19567" *)
  wire [7:0] _04350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19577" *)
  wire [7:0] _04351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19587" *)
  wire [7:0] _04352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19597" *)
  wire [7:0] _04353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19607" *)
  wire [7:0] _04354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19617" *)
  wire [7:0] _04355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19627" *)
  wire [7:0] _04356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19637" *)
  wire [7:0] _04357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19647" *)
  wire [7:0] _04358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19657" *)
  wire [7:0] _04359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19667" *)
  wire [7:0] _04360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19677" *)
  wire [7:0] _04361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19687" *)
  wire [7:0] _04362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19697" *)
  wire [7:0] _04363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19707" *)
  wire [7:0] _04364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19717" *)
  wire [7:0] _04365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19727" *)
  wire [7:0] _04366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19737" *)
  wire [7:0] _04367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19747" *)
  wire [7:0] _04368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19757" *)
  wire [7:0] _04369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19767" *)
  wire [7:0] _04370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19777" *)
  wire [7:0] _04371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19787" *)
  wire [7:0] _04372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19797" *)
  wire [7:0] _04373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19807" *)
  wire [7:0] _04374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19817" *)
  wire [7:0] _04375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19827" *)
  wire [7:0] _04376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19837" *)
  wire [7:0] _04377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19847" *)
  wire [7:0] _04378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19857" *)
  wire [7:0] _04379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19867" *)
  wire [7:0] _04380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19877" *)
  wire [7:0] _04381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19887" *)
  wire [7:0] _04382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19897" *)
  wire [7:0] _04383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19907" *)
  wire [7:0] _04384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19917" *)
  wire [7:0] _04385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19927" *)
  wire [7:0] _04386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19937" *)
  wire [7:0] _04387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19947" *)
  wire [7:0] _04388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19957" *)
  wire [7:0] _04389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19967" *)
  wire [7:0] _04390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20000" *)
  wire _04391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20010" *)
  wire _04392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20021" *)
  wire [7:0] _04393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20031" *)
  wire [7:0] _04394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20041" *)
  wire [7:0] _04395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20051" *)
  wire [7:0] _04396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20061" *)
  wire [7:0] _04397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20071" *)
  wire [7:0] _04398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20081" *)
  wire [7:0] _04399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20091" *)
  wire [7:0] _04400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20101" *)
  wire [7:0] _04401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20111" *)
  wire [7:0] _04402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20121" *)
  wire [7:0] _04403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20131" *)
  wire [7:0] _04404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20141" *)
  wire [7:0] _04405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20151" *)
  wire [7:0] _04406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20161" *)
  wire [7:0] _04407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20171" *)
  wire [7:0] _04408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20181" *)
  wire [7:0] _04409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20191" *)
  wire [7:0] _04410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20201" *)
  wire [7:0] _04411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20211" *)
  wire [7:0] _04412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20221" *)
  wire [7:0] _04413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20231" *)
  wire [7:0] _04414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20241" *)
  wire [7:0] _04415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20251" *)
  wire [7:0] _04416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20261" *)
  wire [7:0] _04417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20271" *)
  wire [7:0] _04418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20281" *)
  wire [7:0] _04419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20291" *)
  wire [7:0] _04420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20301" *)
  wire [7:0] _04421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20311" *)
  wire [7:0] _04422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20321" *)
  wire [7:0] _04423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20331" *)
  wire [7:0] _04424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20341" *)
  wire [7:0] _04425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20351" *)
  wire [7:0] _04426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20361" *)
  wire [7:0] _04427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20371" *)
  wire [7:0] _04428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20381" *)
  wire [7:0] _04429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20391" *)
  wire [7:0] _04430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20401" *)
  wire [7:0] _04431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20411" *)
  wire [7:0] _04432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20421" *)
  wire [7:0] _04433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20431" *)
  wire [7:0] _04434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20441" *)
  wire [7:0] _04435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20451" *)
  wire [7:0] _04436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20461" *)
  wire [7:0] _04437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20471" *)
  wire [7:0] _04438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20481" *)
  wire [7:0] _04439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20491" *)
  wire [7:0] _04440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20501" *)
  wire [7:0] _04441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20511" *)
  wire [7:0] _04442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20521" *)
  wire [7:0] _04443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20531" *)
  wire [7:0] _04444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20541" *)
  wire [7:0] _04445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20551" *)
  wire [7:0] _04446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20561" *)
  wire [7:0] _04447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20571" *)
  wire [7:0] _04448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20581" *)
  wire [7:0] _04449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20591" *)
  wire [7:0] _04450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20601" *)
  wire [7:0] _04451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20611" *)
  wire [7:0] _04452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20621" *)
  wire [7:0] _04453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20631" *)
  wire [7:0] _04454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20641" *)
  wire [7:0] _04455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20651" *)
  wire [7:0] _04456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20661" *)
  wire [7:0] _04457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20671" *)
  wire [7:0] _04458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20681" *)
  wire [7:0] _04459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20691" *)
  wire [7:0] _04460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20701" *)
  wire [7:0] _04461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20711" *)
  wire [7:0] _04462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20721" *)
  wire [7:0] _04463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20731" *)
  wire [7:0] _04464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20741" *)
  wire [7:0] _04465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20751" *)
  wire [7:0] _04466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20761" *)
  wire [7:0] _04467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20771" *)
  wire [7:0] _04468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20781" *)
  wire [7:0] _04469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20791" *)
  wire [7:0] _04470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20801" *)
  wire [7:0] _04471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20811" *)
  wire [7:0] _04472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20821" *)
  wire [7:0] _04473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20831" *)
  wire [7:0] _04474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20841" *)
  wire [7:0] _04475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20851" *)
  wire [7:0] _04476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20861" *)
  wire [7:0] _04477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20871" *)
  wire [7:0] _04478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20881" *)
  wire [7:0] _04479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20891" *)
  wire [7:0] _04480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20901" *)
  wire [7:0] _04481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20911" *)
  wire [7:0] _04482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20921" *)
  wire [7:0] _04483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20931" *)
  wire [7:0] _04484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20941" *)
  wire [7:0] _04485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20951" *)
  wire [7:0] _04486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20961" *)
  wire [7:0] _04487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20971" *)
  wire [7:0] _04488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20981" *)
  wire [7:0] _04489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20991" *)
  wire [7:0] _04490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21001" *)
  wire [7:0] _04491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21011" *)
  wire [7:0] _04492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21021" *)
  wire [7:0] _04493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21031" *)
  wire [7:0] _04494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21041" *)
  wire [7:0] _04495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21051" *)
  wire [7:0] _04496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21061" *)
  wire [7:0] _04497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21071" *)
  wire [7:0] _04498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21081" *)
  wire [7:0] _04499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21091" *)
  wire [7:0] _04500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21101" *)
  wire [7:0] _04501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21111" *)
  wire [7:0] _04502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21121" *)
  wire [7:0] _04503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21131" *)
  wire [7:0] _04504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21141" *)
  wire [7:0] _04505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21151" *)
  wire [7:0] _04506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21161" *)
  wire [7:0] _04507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21171" *)
  wire [7:0] _04508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21181" *)
  wire [7:0] _04509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21191" *)
  wire [7:0] _04510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21201" *)
  wire [7:0] _04511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21211" *)
  wire [7:0] _04512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21221" *)
  wire [7:0] _04513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21231" *)
  wire [7:0] _04514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21241" *)
  wire [7:0] _04515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21251" *)
  wire [7:0] _04516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21261" *)
  wire [7:0] _04517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21271" *)
  wire [7:0] _04518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21281" *)
  wire [7:0] _04519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21291" *)
  wire [7:0] _04520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21324" *)
  wire _04521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21334" *)
  wire _04522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21345" *)
  wire [7:0] _04523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21355" *)
  wire [7:0] _04524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21365" *)
  wire [7:0] _04525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21375" *)
  wire [7:0] _04526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21385" *)
  wire [7:0] _04527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21395" *)
  wire [7:0] _04528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21405" *)
  wire [7:0] _04529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21415" *)
  wire [7:0] _04530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21425" *)
  wire [7:0] _04531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21435" *)
  wire [7:0] _04532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21445" *)
  wire [7:0] _04533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21455" *)
  wire [7:0] _04534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21465" *)
  wire [7:0] _04535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21475" *)
  wire [7:0] _04536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21485" *)
  wire [7:0] _04537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21495" *)
  wire [7:0] _04538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21505" *)
  wire [7:0] _04539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21515" *)
  wire [7:0] _04540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21525" *)
  wire [7:0] _04541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21535" *)
  wire [7:0] _04542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21545" *)
  wire [7:0] _04543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21555" *)
  wire [7:0] _04544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21565" *)
  wire [7:0] _04545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21575" *)
  wire [7:0] _04546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21585" *)
  wire [7:0] _04547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21595" *)
  wire [7:0] _04548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21605" *)
  wire [7:0] _04549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21615" *)
  wire [7:0] _04550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21625" *)
  wire [7:0] _04551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21635" *)
  wire [7:0] _04552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21645" *)
  wire [7:0] _04553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21655" *)
  wire [7:0] _04554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21665" *)
  wire [7:0] _04555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21675" *)
  wire [7:0] _04556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21685" *)
  wire [7:0] _04557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21695" *)
  wire [7:0] _04558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21705" *)
  wire [7:0] _04559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21715" *)
  wire [7:0] _04560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21725" *)
  wire [7:0] _04561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21735" *)
  wire [7:0] _04562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21745" *)
  wire [7:0] _04563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21755" *)
  wire [7:0] _04564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21765" *)
  wire [7:0] _04565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21775" *)
  wire [7:0] _04566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21785" *)
  wire [7:0] _04567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21795" *)
  wire [7:0] _04568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21805" *)
  wire [7:0] _04569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21815" *)
  wire [7:0] _04570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21825" *)
  wire [7:0] _04571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21835" *)
  wire [7:0] _04572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21845" *)
  wire [7:0] _04573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21855" *)
  wire [7:0] _04574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21865" *)
  wire [7:0] _04575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21875" *)
  wire [7:0] _04576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21885" *)
  wire [7:0] _04577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21895" *)
  wire [7:0] _04578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21905" *)
  wire [7:0] _04579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21915" *)
  wire [7:0] _04580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21925" *)
  wire [7:0] _04581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21935" *)
  wire [7:0] _04582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21945" *)
  wire [7:0] _04583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21955" *)
  wire [7:0] _04584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21965" *)
  wire [7:0] _04585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21975" *)
  wire [7:0] _04586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21985" *)
  wire [7:0] _04587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21995" *)
  wire [7:0] _04588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22005" *)
  wire [7:0] _04589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22015" *)
  wire [7:0] _04590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22025" *)
  wire [7:0] _04591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22035" *)
  wire [7:0] _04592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22045" *)
  wire [7:0] _04593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22055" *)
  wire [7:0] _04594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22065" *)
  wire [7:0] _04595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22075" *)
  wire [7:0] _04596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22085" *)
  wire [7:0] _04597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22095" *)
  wire [7:0] _04598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22105" *)
  wire [7:0] _04599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22115" *)
  wire [7:0] _04600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22125" *)
  wire [7:0] _04601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22135" *)
  wire [7:0] _04602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22145" *)
  wire [7:0] _04603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22155" *)
  wire [7:0] _04604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22165" *)
  wire [7:0] _04605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22175" *)
  wire [7:0] _04606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22185" *)
  wire [7:0] _04607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22195" *)
  wire [7:0] _04608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22205" *)
  wire [7:0] _04609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22215" *)
  wire [7:0] _04610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22225" *)
  wire [7:0] _04611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22235" *)
  wire [7:0] _04612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22245" *)
  wire [7:0] _04613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22255" *)
  wire [7:0] _04614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22265" *)
  wire [7:0] _04615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22275" *)
  wire [7:0] _04616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22285" *)
  wire [7:0] _04617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22295" *)
  wire [7:0] _04618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22305" *)
  wire [7:0] _04619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22315" *)
  wire [7:0] _04620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22325" *)
  wire [7:0] _04621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22335" *)
  wire [7:0] _04622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22345" *)
  wire [7:0] _04623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22355" *)
  wire [7:0] _04624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22365" *)
  wire [7:0] _04625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22375" *)
  wire [7:0] _04626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22385" *)
  wire [7:0] _04627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22395" *)
  wire [7:0] _04628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22405" *)
  wire [7:0] _04629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22415" *)
  wire [7:0] _04630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22425" *)
  wire [7:0] _04631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22435" *)
  wire [7:0] _04632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22445" *)
  wire [7:0] _04633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22455" *)
  wire [7:0] _04634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22465" *)
  wire [7:0] _04635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22475" *)
  wire [7:0] _04636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22485" *)
  wire [7:0] _04637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22495" *)
  wire [7:0] _04638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22505" *)
  wire [7:0] _04639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22515" *)
  wire [7:0] _04640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22525" *)
  wire [7:0] _04641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22535" *)
  wire [7:0] _04642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22545" *)
  wire [7:0] _04643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22555" *)
  wire [7:0] _04644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22565" *)
  wire [7:0] _04645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22575" *)
  wire [7:0] _04646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22585" *)
  wire [7:0] _04647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22595" *)
  wire [7:0] _04648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22605" *)
  wire [7:0] _04649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22615" *)
  wire [7:0] _04650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22648" *)
  wire _04651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22658" *)
  wire _04652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22669" *)
  wire [7:0] _04653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22679" *)
  wire [7:0] _04654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22689" *)
  wire [7:0] _04655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22699" *)
  wire [7:0] _04656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22709" *)
  wire [7:0] _04657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22719" *)
  wire [7:0] _04658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22729" *)
  wire [7:0] _04659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22739" *)
  wire [7:0] _04660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22749" *)
  wire [7:0] _04661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22759" *)
  wire [7:0] _04662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22769" *)
  wire [7:0] _04663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22779" *)
  wire [7:0] _04664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22789" *)
  wire [7:0] _04665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22799" *)
  wire [7:0] _04666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22809" *)
  wire [7:0] _04667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22819" *)
  wire [7:0] _04668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22829" *)
  wire [7:0] _04669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22839" *)
  wire [7:0] _04670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22849" *)
  wire [7:0] _04671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22859" *)
  wire [7:0] _04672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22869" *)
  wire [7:0] _04673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22879" *)
  wire [7:0] _04674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22889" *)
  wire [7:0] _04675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22899" *)
  wire [7:0] _04676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22909" *)
  wire [7:0] _04677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22919" *)
  wire [7:0] _04678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22929" *)
  wire [7:0] _04679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22939" *)
  wire [7:0] _04680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22949" *)
  wire [7:0] _04681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22959" *)
  wire [7:0] _04682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22969" *)
  wire [7:0] _04683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22979" *)
  wire [7:0] _04684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22989" *)
  wire [7:0] _04685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22999" *)
  wire [7:0] _04686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23009" *)
  wire [7:0] _04687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23019" *)
  wire [7:0] _04688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23029" *)
  wire [7:0] _04689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23039" *)
  wire [7:0] _04690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23049" *)
  wire [7:0] _04691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23059" *)
  wire [7:0] _04692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23069" *)
  wire [7:0] _04693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23079" *)
  wire [7:0] _04694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23089" *)
  wire [7:0] _04695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23099" *)
  wire [7:0] _04696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23109" *)
  wire [7:0] _04697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23119" *)
  wire [7:0] _04698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23129" *)
  wire [7:0] _04699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23139" *)
  wire [7:0] _04700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23149" *)
  wire [7:0] _04701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23159" *)
  wire [7:0] _04702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23169" *)
  wire [7:0] _04703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23179" *)
  wire [7:0] _04704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23189" *)
  wire [7:0] _04705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23199" *)
  wire [7:0] _04706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23209" *)
  wire [7:0] _04707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23219" *)
  wire [7:0] _04708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23229" *)
  wire [7:0] _04709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23239" *)
  wire [7:0] _04710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23249" *)
  wire [7:0] _04711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23259" *)
  wire [7:0] _04712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23269" *)
  wire [7:0] _04713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23279" *)
  wire [7:0] _04714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23289" *)
  wire [7:0] _04715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23299" *)
  wire [7:0] _04716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23309" *)
  wire [7:0] _04717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23319" *)
  wire [7:0] _04718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23329" *)
  wire [7:0] _04719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23339" *)
  wire [7:0] _04720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23349" *)
  wire [7:0] _04721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23359" *)
  wire [7:0] _04722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23369" *)
  wire [7:0] _04723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23379" *)
  wire [7:0] _04724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23389" *)
  wire [7:0] _04725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23399" *)
  wire [7:0] _04726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23409" *)
  wire [7:0] _04727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23419" *)
  wire [7:0] _04728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23429" *)
  wire [7:0] _04729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23439" *)
  wire [7:0] _04730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23449" *)
  wire [7:0] _04731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23459" *)
  wire [7:0] _04732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23469" *)
  wire [7:0] _04733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23479" *)
  wire [7:0] _04734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23489" *)
  wire [7:0] _04735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23499" *)
  wire [7:0] _04736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23509" *)
  wire [7:0] _04737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23519" *)
  wire [7:0] _04738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23529" *)
  wire [7:0] _04739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23539" *)
  wire [7:0] _04740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23549" *)
  wire [7:0] _04741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23559" *)
  wire [7:0] _04742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23569" *)
  wire [7:0] _04743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23579" *)
  wire [7:0] _04744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23589" *)
  wire [7:0] _04745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23599" *)
  wire [7:0] _04746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23609" *)
  wire [7:0] _04747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23619" *)
  wire [7:0] _04748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23629" *)
  wire [7:0] _04749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23639" *)
  wire [7:0] _04750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23649" *)
  wire [7:0] _04751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23659" *)
  wire [7:0] _04752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23669" *)
  wire [7:0] _04753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23679" *)
  wire [7:0] _04754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23689" *)
  wire [7:0] _04755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23699" *)
  wire [7:0] _04756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23709" *)
  wire [7:0] _04757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23719" *)
  wire [7:0] _04758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23729" *)
  wire [7:0] _04759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23739" *)
  wire [7:0] _04760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23749" *)
  wire [7:0] _04761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23759" *)
  wire [7:0] _04762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23769" *)
  wire [7:0] _04763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23779" *)
  wire [7:0] _04764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23789" *)
  wire [7:0] _04765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23799" *)
  wire [7:0] _04766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23809" *)
  wire [7:0] _04767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23819" *)
  wire [7:0] _04768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23829" *)
  wire [7:0] _04769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23839" *)
  wire [7:0] _04770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23849" *)
  wire [7:0] _04771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23859" *)
  wire [7:0] _04772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23869" *)
  wire [7:0] _04773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23879" *)
  wire [7:0] _04774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23889" *)
  wire [7:0] _04775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23899" *)
  wire [7:0] _04776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23909" *)
  wire [7:0] _04777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23919" *)
  wire [7:0] _04778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23929" *)
  wire [7:0] _04779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23939" *)
  wire [7:0] _04780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23972" *)
  wire _04781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23982" *)
  wire _04782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23993" *)
  wire [7:0] _04783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24003" *)
  wire [7:0] _04784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24013" *)
  wire [7:0] _04785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24023" *)
  wire [7:0] _04786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24033" *)
  wire [7:0] _04787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24043" *)
  wire [7:0] _04788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24053" *)
  wire [7:0] _04789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24063" *)
  wire [7:0] _04790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24073" *)
  wire [7:0] _04791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24083" *)
  wire [7:0] _04792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24093" *)
  wire [7:0] _04793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24103" *)
  wire [7:0] _04794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24113" *)
  wire [7:0] _04795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24123" *)
  wire [7:0] _04796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24133" *)
  wire [7:0] _04797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24143" *)
  wire [7:0] _04798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24153" *)
  wire [7:0] _04799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24163" *)
  wire [7:0] _04800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24173" *)
  wire [7:0] _04801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24183" *)
  wire [7:0] _04802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24193" *)
  wire [7:0] _04803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24203" *)
  wire [7:0] _04804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24213" *)
  wire [7:0] _04805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24223" *)
  wire [7:0] _04806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24233" *)
  wire [7:0] _04807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24243" *)
  wire [7:0] _04808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24253" *)
  wire [7:0] _04809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24263" *)
  wire [7:0] _04810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24273" *)
  wire [7:0] _04811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24283" *)
  wire [7:0] _04812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24293" *)
  wire [7:0] _04813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24303" *)
  wire [7:0] _04814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24313" *)
  wire [7:0] _04815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24323" *)
  wire [7:0] _04816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24333" *)
  wire [7:0] _04817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24343" *)
  wire [7:0] _04818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24353" *)
  wire [7:0] _04819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24363" *)
  wire [7:0] _04820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24373" *)
  wire [7:0] _04821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24383" *)
  wire [7:0] _04822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24393" *)
  wire [7:0] _04823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24403" *)
  wire [7:0] _04824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24413" *)
  wire [7:0] _04825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24423" *)
  wire [7:0] _04826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24433" *)
  wire [7:0] _04827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24443" *)
  wire [7:0] _04828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24453" *)
  wire [7:0] _04829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24463" *)
  wire [7:0] _04830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24473" *)
  wire [7:0] _04831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24483" *)
  wire [7:0] _04832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24493" *)
  wire [7:0] _04833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24503" *)
  wire [7:0] _04834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24513" *)
  wire [7:0] _04835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24523" *)
  wire [7:0] _04836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24533" *)
  wire [7:0] _04837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24543" *)
  wire [7:0] _04838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24553" *)
  wire [7:0] _04839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24563" *)
  wire [7:0] _04840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24573" *)
  wire [7:0] _04841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24583" *)
  wire [7:0] _04842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24593" *)
  wire [7:0] _04843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24603" *)
  wire [7:0] _04844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24613" *)
  wire [7:0] _04845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24623" *)
  wire [7:0] _04846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24633" *)
  wire [7:0] _04847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24643" *)
  wire [7:0] _04848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24653" *)
  wire [7:0] _04849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24663" *)
  wire [7:0] _04850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24673" *)
  wire [7:0] _04851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24683" *)
  wire [7:0] _04852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24693" *)
  wire [7:0] _04853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24703" *)
  wire [7:0] _04854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24713" *)
  wire [7:0] _04855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24723" *)
  wire [7:0] _04856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24733" *)
  wire [7:0] _04857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24743" *)
  wire [7:0] _04858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24753" *)
  wire [7:0] _04859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24763" *)
  wire [7:0] _04860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24773" *)
  wire [7:0] _04861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24783" *)
  wire [7:0] _04862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24793" *)
  wire [7:0] _04863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24803" *)
  wire [7:0] _04864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24813" *)
  wire [7:0] _04865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24823" *)
  wire [7:0] _04866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24833" *)
  wire [7:0] _04867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24843" *)
  wire [7:0] _04868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24853" *)
  wire [7:0] _04869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24863" *)
  wire [7:0] _04870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24873" *)
  wire [7:0] _04871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24883" *)
  wire [7:0] _04872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24893" *)
  wire [7:0] _04873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24903" *)
  wire [7:0] _04874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24913" *)
  wire [7:0] _04875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24923" *)
  wire [7:0] _04876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24933" *)
  wire [7:0] _04877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24943" *)
  wire [7:0] _04878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24953" *)
  wire [7:0] _04879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24963" *)
  wire [7:0] _04880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24973" *)
  wire [7:0] _04881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24983" *)
  wire [7:0] _04882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24993" *)
  wire [7:0] _04883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25003" *)
  wire [7:0] _04884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25013" *)
  wire [7:0] _04885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25023" *)
  wire [7:0] _04886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25033" *)
  wire [7:0] _04887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25043" *)
  wire [7:0] _04888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25053" *)
  wire [7:0] _04889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25063" *)
  wire [7:0] _04890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25073" *)
  wire [7:0] _04891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25083" *)
  wire [7:0] _04892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25093" *)
  wire [7:0] _04893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25103" *)
  wire [7:0] _04894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25113" *)
  wire [7:0] _04895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25123" *)
  wire [7:0] _04896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25133" *)
  wire [7:0] _04897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25143" *)
  wire [7:0] _04898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25153" *)
  wire [7:0] _04899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25163" *)
  wire [7:0] _04900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25173" *)
  wire [7:0] _04901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25183" *)
  wire [7:0] _04902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25193" *)
  wire [7:0] _04903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25203" *)
  wire [7:0] _04904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25213" *)
  wire [7:0] _04905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25223" *)
  wire [7:0] _04906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25233" *)
  wire [7:0] _04907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25243" *)
  wire [7:0] _04908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25253" *)
  wire [7:0] _04909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25263" *)
  wire [7:0] _04910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25296" *)
  wire _04911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25306" *)
  wire _04912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25317" *)
  wire [7:0] _04913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25327" *)
  wire [7:0] _04914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25337" *)
  wire [7:0] _04915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25347" *)
  wire [7:0] _04916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25357" *)
  wire [7:0] _04917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25367" *)
  wire [7:0] _04918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25377" *)
  wire [7:0] _04919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25387" *)
  wire [7:0] _04920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25397" *)
  wire [7:0] _04921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25407" *)
  wire [7:0] _04922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25417" *)
  wire [7:0] _04923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25427" *)
  wire [7:0] _04924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25437" *)
  wire [7:0] _04925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25447" *)
  wire [7:0] _04926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25457" *)
  wire [7:0] _04927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25467" *)
  wire [7:0] _04928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25477" *)
  wire [7:0] _04929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25487" *)
  wire [7:0] _04930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25497" *)
  wire [7:0] _04931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25507" *)
  wire [7:0] _04932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25517" *)
  wire [7:0] _04933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25527" *)
  wire [7:0] _04934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25537" *)
  wire [7:0] _04935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25547" *)
  wire [7:0] _04936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25557" *)
  wire [7:0] _04937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25567" *)
  wire [7:0] _04938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25577" *)
  wire [7:0] _04939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25587" *)
  wire [7:0] _04940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25597" *)
  wire [7:0] _04941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25607" *)
  wire [7:0] _04942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25617" *)
  wire [7:0] _04943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25627" *)
  wire [7:0] _04944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25637" *)
  wire [7:0] _04945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25647" *)
  wire [7:0] _04946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25657" *)
  wire [7:0] _04947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25667" *)
  wire [7:0] _04948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25677" *)
  wire [7:0] _04949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25687" *)
  wire [7:0] _04950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25697" *)
  wire [7:0] _04951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25707" *)
  wire [7:0] _04952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25717" *)
  wire [7:0] _04953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25727" *)
  wire [7:0] _04954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25737" *)
  wire [7:0] _04955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25747" *)
  wire [7:0] _04956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25757" *)
  wire [7:0] _04957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25767" *)
  wire [7:0] _04958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25777" *)
  wire [7:0] _04959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25787" *)
  wire [7:0] _04960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25797" *)
  wire [7:0] _04961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25807" *)
  wire [7:0] _04962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25817" *)
  wire [7:0] _04963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25827" *)
  wire [7:0] _04964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25837" *)
  wire [7:0] _04965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25847" *)
  wire [7:0] _04966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25857" *)
  wire [7:0] _04967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25867" *)
  wire [7:0] _04968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25877" *)
  wire [7:0] _04969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *)
  wire _04970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *)
  wire _04971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25887" *)
  wire [7:0] _04972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *)
  wire _04973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *)
  wire _04974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25897" *)
  wire [7:0] _04975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *)
  wire _04976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *)
  wire _04977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25907" *)
  wire [7:0] _04978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *)
  wire _04979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *)
  wire _04980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25917" *)
  wire [7:0] _04981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *)
  wire _04982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *)
  wire _04983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25927" *)
  wire [7:0] _04984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *)
  wire _04985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *)
  wire _04986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25937" *)
  wire [7:0] _04987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *)
  wire _04988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *)
  wire _04989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25947" *)
  wire [7:0] _04990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *)
  wire _04991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *)
  wire _04992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25957" *)
  wire [7:0] _04993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *)
  wire _04994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *)
  wire _04995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25967" *)
  wire [7:0] _04996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *)
  wire _04997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *)
  wire _04998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25977" *)
  wire [7:0] _04999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *)
  wire _05000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *)
  wire _05001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25987" *)
  wire [7:0] _05002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *)
  wire _05003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *)
  wire _05004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25997" *)
  wire [7:0] _05005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *)
  wire _05006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *)
  wire _05007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26007" *)
  wire [7:0] _05008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *)
  wire _05009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *)
  wire _05010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26017" *)
  wire [7:0] _05011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *)
  wire _05012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *)
  wire _05013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26027" *)
  wire [7:0] _05014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *)
  wire _05015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *)
  wire _05016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26037" *)
  wire [7:0] _05017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *)
  wire _05018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *)
  wire _05019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26047" *)
  wire [7:0] _05020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *)
  wire _05021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *)
  wire _05022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26057" *)
  wire [7:0] _05023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *)
  wire _05024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *)
  wire _05025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26067" *)
  wire [7:0] _05026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *)
  wire _05027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *)
  wire _05028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26077" *)
  wire [7:0] _05029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *)
  wire _05030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *)
  wire _05031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26087" *)
  wire [7:0] _05032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *)
  wire _05033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *)
  wire _05034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26097" *)
  wire [7:0] _05035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *)
  wire _05036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *)
  wire _05037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26107" *)
  wire [7:0] _05038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *)
  wire _05039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *)
  wire _05040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26117" *)
  wire [7:0] _05041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *)
  wire _05042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *)
  wire _05043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26127" *)
  wire [7:0] _05044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *)
  wire _05045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *)
  wire _05046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26137" *)
  wire [7:0] _05047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *)
  wire _05048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *)
  wire _05049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26147" *)
  wire [7:0] _05050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *)
  wire _05051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *)
  wire _05052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26157" *)
  wire [7:0] _05053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *)
  wire _05054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *)
  wire _05055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26167" *)
  wire [7:0] _05056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *)
  wire _05057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *)
  wire _05058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26177" *)
  wire [7:0] _05059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *)
  wire _05060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *)
  wire _05061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26187" *)
  wire [7:0] _05062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *)
  wire _05063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *)
  wire _05064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26197" *)
  wire [7:0] _05065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *)
  wire _05066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *)
  wire _05067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26207" *)
  wire [7:0] _05068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *)
  wire _05069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *)
  wire _05070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26217" *)
  wire [7:0] _05071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *)
  wire _05072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *)
  wire _05073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26227" *)
  wire [7:0] _05074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *)
  wire _05075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *)
  wire _05076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26237" *)
  wire [7:0] _05077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *)
  wire _05078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *)
  wire _05079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26247" *)
  wire [7:0] _05080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *)
  wire _05081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *)
  wire _05082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26257" *)
  wire [7:0] _05083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *)
  wire _05084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *)
  wire _05085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26267" *)
  wire [7:0] _05086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *)
  wire _05087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *)
  wire _05088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26277" *)
  wire [7:0] _05089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *)
  wire _05090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *)
  wire _05091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26287" *)
  wire [7:0] _05092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *)
  wire _05093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *)
  wire _05094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26297" *)
  wire [7:0] _05095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *)
  wire _05096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *)
  wire _05097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26307" *)
  wire [7:0] _05098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *)
  wire _05099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *)
  wire _05100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26317" *)
  wire [7:0] _05101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *)
  wire _05102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *)
  wire _05103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26327" *)
  wire [7:0] _05104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *)
  wire _05105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *)
  wire _05106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26337" *)
  wire [7:0] _05107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *)
  wire _05108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *)
  wire _05109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26347" *)
  wire [7:0] _05110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *)
  wire _05111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *)
  wire _05112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26357" *)
  wire [7:0] _05113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *)
  wire _05114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *)
  wire _05115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26367" *)
  wire [7:0] _05116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *)
  wire _05117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *)
  wire _05118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26377" *)
  wire [7:0] _05119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *)
  wire _05120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *)
  wire _05121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26387" *)
  wire [7:0] _05122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *)
  wire _05123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *)
  wire _05124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26397" *)
  wire [7:0] _05125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *)
  wire _05126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *)
  wire _05127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26407" *)
  wire [7:0] _05128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *)
  wire _05129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *)
  wire _05130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26417" *)
  wire [7:0] _05131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *)
  wire _05132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *)
  wire _05133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26427" *)
  wire [7:0] _05134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *)
  wire _05135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *)
  wire _05136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26437" *)
  wire [7:0] _05137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *)
  wire _05138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *)
  wire _05139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26447" *)
  wire [7:0] _05140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *)
  wire _05141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *)
  wire _05142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26457" *)
  wire [7:0] _05143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *)
  wire _05144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *)
  wire _05145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26467" *)
  wire [7:0] _05146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *)
  wire _05147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *)
  wire _05148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26477" *)
  wire [7:0] _05149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *)
  wire _05150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *)
  wire _05151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26487" *)
  wire [7:0] _05152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *)
  wire _05153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *)
  wire _05154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26497" *)
  wire [7:0] _05155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *)
  wire _05156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *)
  wire _05157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26507" *)
  wire [7:0] _05158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *)
  wire _05159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *)
  wire _05160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26517" *)
  wire [7:0] _05161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26527" *)
  wire [7:0] _05162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26537" *)
  wire [7:0] _05163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26547" *)
  wire [7:0] _05164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26557" *)
  wire [7:0] _05165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26567" *)
  wire [7:0] _05166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26577" *)
  wire [7:0] _05167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2658" *)
  wire _05168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26587" *)
  wire [7:0] _05169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2659" *)
  wire _05170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2660" *)
  wire _05171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2661" *)
  wire _05172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2662" *)
  wire _05173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2663" *)
  wire _05174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2664" *)
  wire _05175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2665" *)
  wire _05176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2666" *)
  wire _05177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2667" *)
  wire _05178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2668" *)
  wire _05179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2669" *)
  wire _05180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2670" *)
  wire _05181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2671" *)
  wire _05182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2672" *)
  wire _05183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2673" *)
  wire _05184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2674" *)
  wire _05185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2675" *)
  wire _05186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2676" *)
  wire _05187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2677" *)
  wire _05188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2678" *)
  wire _05189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2679" *)
  wire _05190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2680" *)
  wire _05191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2681" *)
  wire _05192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2682" *)
  wire _05193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2683" *)
  wire _05194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2684" *)
  wire _05195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2685" *)
  wire _05196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2686" *)
  wire _05197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2687" *)
  wire _05198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2688" *)
  wire _05199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2689" *)
  wire _05200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2690" *)
  wire _05201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2691" *)
  wire _05202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2692" *)
  wire _05203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2693" *)
  wire _05204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2694" *)
  wire _05205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2695" *)
  wire _05206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2696" *)
  wire _05207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2697" *)
  wire _05208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2698" *)
  wire _05209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2699" *)
  wire _05210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2700" *)
  wire _05211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2701" *)
  wire _05212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2702" *)
  wire _05213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2703" *)
  wire _05214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2704" *)
  wire _05215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2705" *)
  wire _05216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2706" *)
  wire _05217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2707" *)
  wire _05218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2708" *)
  wire _05219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2709" *)
  wire _05220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2710" *)
  wire _05221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2711" *)
  wire _05222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2712" *)
  wire _05223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2713" *)
  wire _05224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2714" *)
  wire _05225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2715" *)
  wire _05226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2716" *)
  wire _05227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2717" *)
  wire _05228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2718" *)
  wire _05229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2719" *)
  wire _05230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2720" *)
  wire _05231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2721" *)
  wire _05232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *)
  wire _05233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *)
  wire _05234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *)
  wire _05235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *)
  wire _05236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *)
  wire _05237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *)
  wire _05238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *)
  wire _05239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *)
  wire _05240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *)
  wire _05241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *)
  wire _05242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *)
  wire _05243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *)
  wire _05244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *)
  wire _05245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *)
  wire _05246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *)
  wire _05247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *)
  wire _05248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *)
  wire _05249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *)
  wire _05250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *)
  wire _05251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *)
  wire _05252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *)
  wire _05253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *)
  wire _05254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *)
  wire _05255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *)
  wire _05256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *)
  wire _05257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *)
  wire _05258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *)
  wire _05259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *)
  wire _05260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *)
  wire _05261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *)
  wire _05262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *)
  wire _05263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *)
  wire _05264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *)
  wire _05265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *)
  wire _05266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *)
  wire _05267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *)
  wire _05268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *)
  wire _05269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *)
  wire _05270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *)
  wire _05271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *)
  wire _05272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *)
  wire _05273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *)
  wire _05274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *)
  wire _05275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *)
  wire _05276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *)
  wire _05277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *)
  wire _05278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *)
  wire _05279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *)
  wire _05280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *)
  wire _05281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *)
  wire _05282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *)
  wire _05283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *)
  wire _05284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *)
  wire _05285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *)
  wire _05286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *)
  wire _05287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *)
  wire _05288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *)
  wire _05289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *)
  wire _05290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *)
  wire _05291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *)
  wire _05292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *)
  wire _05293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *)
  wire _05294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *)
  wire _05295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *)
  wire _05296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *)
  wire _05297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *)
  wire _05298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *)
  wire _05299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *)
  wire _05300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *)
  wire _05301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *)
  wire _05302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *)
  wire _05303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *)
  wire _05304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *)
  wire _05305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *)
  wire _05306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *)
  wire _05307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *)
  wire _05308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *)
  wire _05309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *)
  wire _05310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *)
  wire _05311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *)
  wire _05312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *)
  wire _05313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *)
  wire _05314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *)
  wire _05315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *)
  wire _05316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *)
  wire _05317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *)
  wire _05318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *)
  wire _05319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *)
  wire _05320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *)
  wire _05321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *)
  wire _05322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *)
  wire _05323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *)
  wire _05324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *)
  wire _05325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *)
  wire _05326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *)
  wire _05327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *)
  wire _05328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *)
  wire _05329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *)
  wire _05330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *)
  wire _05331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *)
  wire _05332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *)
  wire _05333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *)
  wire _05334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *)
  wire _05335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *)
  wire _05336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *)
  wire _05337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *)
  wire _05338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *)
  wire _05339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *)
  wire _05340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *)
  wire _05341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *)
  wire _05342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *)
  wire _05343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *)
  wire _05344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *)
  wire _05345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *)
  wire _05346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *)
  wire _05347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *)
  wire _05348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *)
  wire _05349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *)
  wire _05350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *)
  wire _05351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *)
  wire _05352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *)
  wire _05353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *)
  wire _05354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *)
  wire _05355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *)
  wire _05356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *)
  wire _05357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *)
  wire _05358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *)
  wire _05359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *)
  wire _05360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27731" *)
  wire _05361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27732" *)
  wire _05362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27733" *)
  wire _05363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27734" *)
  wire _05364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27735" *)
  wire _05365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27736" *)
  wire _05366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27737" *)
  wire _05367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27738" *)
  wire _05368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27739" *)
  wire _05369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27740" *)
  wire _05370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27741" *)
  wire _05371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27742" *)
  wire _05372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27743" *)
  wire _05373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27744" *)
  wire _05374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27745" *)
  wire _05375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27746" *)
  wire _05376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27747" *)
  wire _05377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27748" *)
  wire _05378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27749" *)
  wire _05379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27750" *)
  wire _05380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27751" *)
  wire _05381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27752" *)
  wire _05382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27753" *)
  wire _05383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27754" *)
  wire _05384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27755" *)
  wire _05385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27756" *)
  wire _05386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27757" *)
  wire _05387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27758" *)
  wire _05388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27759" *)
  wire _05389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27760" *)
  wire _05390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27761" *)
  wire _05391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27762" *)
  wire _05392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27763" *)
  wire _05393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27764" *)
  wire _05394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27765" *)
  wire _05395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27766" *)
  wire _05396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27767" *)
  wire _05397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27768" *)
  wire _05398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27769" *)
  wire _05399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27770" *)
  wire _05400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27771" *)
  wire _05401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27772" *)
  wire _05402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27773" *)
  wire _05403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27774" *)
  wire _05404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27775" *)
  wire _05405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27776" *)
  wire _05406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27777" *)
  wire _05407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27778" *)
  wire _05408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27779" *)
  wire _05409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27780" *)
  wire _05410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27781" *)
  wire _05411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27782" *)
  wire _05412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27783" *)
  wire _05413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27784" *)
  wire _05414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27785" *)
  wire _05415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27786" *)
  wire _05416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27787" *)
  wire _05417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27788" *)
  wire _05418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27789" *)
  wire _05419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27790" *)
  wire _05420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27791" *)
  wire _05421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27792" *)
  wire _05422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27793" *)
  wire _05423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27794" *)
  wire _05424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29041" *)
  wire [127:0] _05425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29076" *)
  wire _05426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29086" *)
  wire _05427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29096" *)
  wire _05428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29106" *)
  wire _05429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29116" *)
  wire _05430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29126" *)
  wire _05431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29136" *)
  wire _05432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29146" *)
  wire _05433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29156" *)
  wire _05434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29166" *)
  wire _05435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29176" *)
  wire _05436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29186" *)
  wire _05437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29196" *)
  wire _05438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29206" *)
  wire _05439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29216" *)
  wire _05440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29226" *)
  wire _05441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29236" *)
  wire _05442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29246" *)
  wire _05443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29256" *)
  wire _05444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29266" *)
  wire _05445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29276" *)
  wire _05446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29286" *)
  wire _05447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29296" *)
  wire _05448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29306" *)
  wire _05449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29316" *)
  wire _05450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29326" *)
  wire _05451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29336" *)
  wire _05452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29346" *)
  wire _05453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29356" *)
  wire _05454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29366" *)
  wire _05455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29376" *)
  wire _05456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29386" *)
  wire _05457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29396" *)
  wire _05458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29406" *)
  wire _05459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29416" *)
  wire _05460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29426" *)
  wire _05461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29436" *)
  wire _05462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29446" *)
  wire _05463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29456" *)
  wire _05464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29466" *)
  wire _05465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29476" *)
  wire _05466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29486" *)
  wire _05467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29496" *)
  wire _05468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29506" *)
  wire _05469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29516" *)
  wire _05470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29526" *)
  wire _05471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29536" *)
  wire _05472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29546" *)
  wire _05473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29556" *)
  wire _05474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29566" *)
  wire _05475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29576" *)
  wire _05476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29586" *)
  wire _05477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29596" *)
  wire _05478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29606" *)
  wire _05479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29616" *)
  wire _05480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29626" *)
  wire _05481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29636" *)
  wire _05482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29646" *)
  wire _05483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29656" *)
  wire _05484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29666" *)
  wire _05485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29676" *)
  wire _05486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29686" *)
  wire _05487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29696" *)
  wire _05488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29706" *)
  wire _05489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29716" *)
  wire _05490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29726" *)
  wire _05491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29736" *)
  wire _05492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29746" *)
  wire _05493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29756" *)
  wire _05494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29766" *)
  wire _05495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29776" *)
  wire _05496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29786" *)
  wire _05497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29796" *)
  wire _05498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29806" *)
  wire _05499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29816" *)
  wire _05500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29826" *)
  wire _05501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29836" *)
  wire _05502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29846" *)
  wire _05503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29856" *)
  wire _05504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29866" *)
  wire _05505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29876" *)
  wire _05506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29886" *)
  wire _05507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29896" *)
  wire _05508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29906" *)
  wire _05509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29916" *)
  wire _05510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29926" *)
  wire _05511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29936" *)
  wire _05512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29946" *)
  wire _05513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29956" *)
  wire _05514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29966" *)
  wire _05515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29976" *)
  wire _05516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29986" *)
  wire _05517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29996" *)
  wire _05518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30006" *)
  wire _05519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30016" *)
  wire _05520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30026" *)
  wire _05521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30036" *)
  wire _05522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30046" *)
  wire _05523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30056" *)
  wire _05524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30066" *)
  wire _05525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30076" *)
  wire _05526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30086" *)
  wire _05527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30096" *)
  wire _05528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30106" *)
  wire _05529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30116" *)
  wire _05530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30126" *)
  wire _05531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30136" *)
  wire _05532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30146" *)
  wire _05533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30156" *)
  wire _05534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30166" *)
  wire _05535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30176" *)
  wire _05536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30186" *)
  wire _05537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30196" *)
  wire _05538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30206" *)
  wire _05539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30216" *)
  wire _05540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30226" *)
  wire _05541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30236" *)
  wire _05542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30246" *)
  wire _05543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30256" *)
  wire _05544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30266" *)
  wire _05545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30276" *)
  wire _05546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30286" *)
  wire _05547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30296" *)
  wire _05548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30306" *)
  wire _05549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30316" *)
  wire _05550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30326" *)
  wire _05551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30336" *)
  wire _05552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30346" *)
  wire _05553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30356" *)
  wire _05554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30380" *)
  wire _05555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30400" *)
  wire _05556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30420" *)
  wire _05557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30440" *)
  wire _05558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30460" *)
  wire _05559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30480" *)
  wire _05560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30500" *)
  wire _05561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30520" *)
  wire _05562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30664" *)
  wire _05563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30674" *)
  wire _05564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30684" *)
  wire _05565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30694" *)
  wire _05566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30704" *)
  wire _05567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30714" *)
  wire _05568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30724" *)
  wire _05569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30734" *)
  wire _05570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30744" *)
  wire _05571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30754" *)
  wire _05572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30764" *)
  wire _05573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30774" *)
  wire _05574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30784" *)
  wire _05575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30794" *)
  wire _05576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30804" *)
  wire _05577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30814" *)
  wire _05578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30824" *)
  wire _05579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30834" *)
  wire _05580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30844" *)
  wire _05581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30854" *)
  wire _05582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30864" *)
  wire _05583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30874" *)
  wire _05584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30884" *)
  wire _05585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30894" *)
  wire _05586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30904" *)
  wire _05587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30914" *)
  wire _05588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30924" *)
  wire _05589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30934" *)
  wire _05590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30944" *)
  wire _05591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30954" *)
  wire _05592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30964" *)
  wire _05593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30974" *)
  wire _05594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30984" *)
  wire _05595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30994" *)
  wire _05596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31004" *)
  wire _05597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31014" *)
  wire _05598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31024" *)
  wire _05599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31034" *)
  wire _05600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31044" *)
  wire _05601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31054" *)
  wire _05602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31064" *)
  wire _05603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31074" *)
  wire _05604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31084" *)
  wire _05605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31094" *)
  wire _05606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31104" *)
  wire _05607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31114" *)
  wire _05608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31124" *)
  wire _05609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31134" *)
  wire _05610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31144" *)
  wire _05611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31154" *)
  wire _05612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31164" *)
  wire _05613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31174" *)
  wire _05614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31184" *)
  wire _05615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31194" *)
  wire _05616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31204" *)
  wire _05617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31214" *)
  wire _05618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31224" *)
  wire _05619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31234" *)
  wire _05620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31244" *)
  wire _05621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31254" *)
  wire _05622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31264" *)
  wire _05623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31274" *)
  wire _05624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31284" *)
  wire _05625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31294" *)
  wire _05626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31304" *)
  wire _05627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31314" *)
  wire _05628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31324" *)
  wire _05629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31334" *)
  wire _05630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31344" *)
  wire _05631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31354" *)
  wire _05632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31364" *)
  wire _05633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31374" *)
  wire _05634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31384" *)
  wire _05635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31394" *)
  wire _05636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31404" *)
  wire _05637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31414" *)
  wire _05638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31424" *)
  wire _05639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31434" *)
  wire _05640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31444" *)
  wire _05641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31454" *)
  wire _05642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31464" *)
  wire _05643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31474" *)
  wire _05644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31484" *)
  wire _05645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31494" *)
  wire _05646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31504" *)
  wire _05647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31514" *)
  wire _05648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31524" *)
  wire _05649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31534" *)
  wire _05650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31544" *)
  wire _05651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31554" *)
  wire _05652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31564" *)
  wire _05653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31574" *)
  wire _05654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31584" *)
  wire _05655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31594" *)
  wire _05656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31604" *)
  wire _05657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31614" *)
  wire _05658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31624" *)
  wire _05659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31634" *)
  wire _05660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31644" *)
  wire _05661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31654" *)
  wire _05662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31664" *)
  wire _05663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31674" *)
  wire _05664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31684" *)
  wire _05665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31694" *)
  wire _05666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31704" *)
  wire _05667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31714" *)
  wire _05668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31724" *)
  wire _05669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31734" *)
  wire _05670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31744" *)
  wire _05671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31754" *)
  wire _05672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31764" *)
  wire _05673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31774" *)
  wire _05674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31784" *)
  wire _05675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31794" *)
  wire _05676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31804" *)
  wire _05677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31814" *)
  wire _05678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31824" *)
  wire _05679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31834" *)
  wire _05680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31844" *)
  wire _05681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31854" *)
  wire _05682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31864" *)
  wire _05683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31874" *)
  wire _05684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31884" *)
  wire _05685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31894" *)
  wire _05686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31904" *)
  wire _05687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31914" *)
  wire _05688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31924" *)
  wire _05689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31934" *)
  wire _05690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31944" *)
  wire _05691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31971" *)
  wire _05692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33278" *)
  wire _05693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34585" *)
  wire _05694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35892" *)
  wire _05695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37199" *)
  wire _05696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38506" *)
  wire _05697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3968" *)
  wire [127:0] _05698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39813" *)
  wire _05699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4003" *)
  wire _05700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4033" *)
  wire _05701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4043" *)
  wire _05702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4053" *)
  wire _05703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4063" *)
  wire _05704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4073" *)
  wire _05705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4083" *)
  wire _05706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4093" *)
  wire _05707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4103" *)
  wire _05708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4113" *)
  wire _05709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4123" *)
  wire _05710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4133" *)
  wire _05711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4143" *)
  wire _05712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4153" *)
  wire _05713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4163" *)
  wire _05714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4173" *)
  wire _05715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4183" *)
  wire _05716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4193" *)
  wire _05717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4203" *)
  wire _05718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4213" *)
  wire _05719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4223" *)
  wire _05720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4233" *)
  wire _05721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4243" *)
  wire _05722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4253" *)
  wire _05723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4263" *)
  wire _05724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4273" *)
  wire _05725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4283" *)
  wire _05726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4293" *)
  wire _05727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4303" *)
  wire _05728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4313" *)
  wire _05729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4323" *)
  wire _05730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4333" *)
  wire _05731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4343" *)
  wire _05732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4353" *)
  wire _05733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4363" *)
  wire _05734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4373" *)
  wire _05735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4383" *)
  wire _05736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4393" *)
  wire _05737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4403" *)
  wire _05738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4413" *)
  wire _05739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4423" *)
  wire _05740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4433" *)
  wire _05741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4443" *)
  wire _05742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4453" *)
  wire _05743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4463" *)
  wire _05744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4473" *)
  wire _05745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4483" *)
  wire _05746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4493" *)
  wire _05747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4503" *)
  wire _05748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4513" *)
  wire _05749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4523" *)
  wire _05750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4533" *)
  wire _05751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4543" *)
  wire _05752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4553" *)
  wire _05753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4563" *)
  wire _05754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4573" *)
  wire _05755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4583" *)
  wire _05756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4593" *)
  wire _05757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4603" *)
  wire _05758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4613" *)
  wire _05759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4623" *)
  wire _05760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4633" *)
  wire _05761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4643" *)
  wire _05762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4653" *)
  wire _05763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4663" *)
  wire _05764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4673" *)
  wire _05765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4683" *)
  wire _05766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4693" *)
  wire _05767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4703" *)
  wire _05768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4713" *)
  wire _05769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4723" *)
  wire _05770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4733" *)
  wire _05771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4743" *)
  wire _05772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4753" *)
  wire _05773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4763" *)
  wire _05774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4773" *)
  wire _05775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4783" *)
  wire _05776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4793" *)
  wire _05777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4803" *)
  wire _05778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4813" *)
  wire _05779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4823" *)
  wire _05780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4833" *)
  wire _05781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4843" *)
  wire _05782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4853" *)
  wire _05783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4863" *)
  wire _05784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4873" *)
  wire _05785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4883" *)
  wire _05786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4893" *)
  wire _05787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4903" *)
  wire _05788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4913" *)
  wire _05789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4923" *)
  wire _05790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4933" *)
  wire _05791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4943" *)
  wire _05792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4953" *)
  wire _05793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4963" *)
  wire _05794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4973" *)
  wire _05795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4983" *)
  wire _05796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4993" *)
  wire _05797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5003" *)
  wire _05798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5013" *)
  wire _05799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5023" *)
  wire _05800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5033" *)
  wire _05801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5043" *)
  wire _05802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5053" *)
  wire _05803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5063" *)
  wire _05804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5073" *)
  wire _05805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5083" *)
  wire _05806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5093" *)
  wire _05807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5103" *)
  wire _05808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5113" *)
  wire _05809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5123" *)
  wire _05810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5133" *)
  wire _05811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5143" *)
  wire _05812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5153" *)
  wire _05813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5163" *)
  wire _05814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5173" *)
  wire _05815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5183" *)
  wire _05816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5193" *)
  wire _05817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5203" *)
  wire _05818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5213" *)
  wire _05819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5223" *)
  wire _05820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5233" *)
  wire _05821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5243" *)
  wire _05822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5253" *)
  wire _05823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5263" *)
  wire _05824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5273" *)
  wire _05825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5283" *)
  wire _05826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5293" *)
  wire _05827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5303" *)
  wire _05828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5342" *)
  wire _05829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5372" *)
  wire _05830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5382" *)
  wire _05831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5392" *)
  wire _05832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5402" *)
  wire _05833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5412" *)
  wire _05834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5422" *)
  wire _05835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5432" *)
  wire _05836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5442" *)
  wire _05837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5452" *)
  wire _05838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5462" *)
  wire _05839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5472" *)
  wire _05840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5482" *)
  wire _05841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5492" *)
  wire _05842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5502" *)
  wire _05843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5512" *)
  wire _05844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5522" *)
  wire _05845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5532" *)
  wire _05846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5542" *)
  wire _05847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5552" *)
  wire _05848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5562" *)
  wire _05849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5572" *)
  wire _05850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5582" *)
  wire _05851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5592" *)
  wire _05852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5602" *)
  wire _05853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5612" *)
  wire _05854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5622" *)
  wire _05855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5632" *)
  wire _05856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5642" *)
  wire _05857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5652" *)
  wire _05858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5662" *)
  wire _05859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5672" *)
  wire _05860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5682" *)
  wire _05861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5692" *)
  wire _05862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5702" *)
  wire _05863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5712" *)
  wire _05864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5722" *)
  wire _05865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5732" *)
  wire _05866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5742" *)
  wire _05867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5752" *)
  wire _05868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5762" *)
  wire _05869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5772" *)
  wire _05870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5782" *)
  wire _05871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5792" *)
  wire _05872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5802" *)
  wire _05873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5812" *)
  wire _05874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5822" *)
  wire _05875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5832" *)
  wire _05876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5842" *)
  wire _05877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5852" *)
  wire _05878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5862" *)
  wire _05879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5872" *)
  wire _05880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5882" *)
  wire _05881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5892" *)
  wire _05882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5902" *)
  wire _05883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5912" *)
  wire _05884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5922" *)
  wire _05885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5932" *)
  wire _05886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5942" *)
  wire _05887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5952" *)
  wire _05888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5962" *)
  wire _05889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5972" *)
  wire _05890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5982" *)
  wire _05891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5992" *)
  wire _05892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6002" *)
  wire _05893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6012" *)
  wire _05894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6022" *)
  wire _05895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6032" *)
  wire _05896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6042" *)
  wire _05897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6052" *)
  wire _05898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6062" *)
  wire _05899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6072" *)
  wire _05900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6082" *)
  wire _05901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6092" *)
  wire _05902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6102" *)
  wire _05903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6112" *)
  wire _05904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6122" *)
  wire _05905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6132" *)
  wire _05906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6142" *)
  wire _05907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6152" *)
  wire _05908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6162" *)
  wire _05909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6172" *)
  wire _05910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6182" *)
  wire _05911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6192" *)
  wire _05912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6202" *)
  wire _05913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6212" *)
  wire _05914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6222" *)
  wire _05915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6232" *)
  wire _05916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6242" *)
  wire _05917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6252" *)
  wire _05918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6262" *)
  wire _05919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6272" *)
  wire _05920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6282" *)
  wire _05921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6292" *)
  wire _05922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6302" *)
  wire _05923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6312" *)
  wire _05924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6322" *)
  wire _05925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6332" *)
  wire _05926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6342" *)
  wire _05927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6352" *)
  wire _05928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6362" *)
  wire _05929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6372" *)
  wire _05930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6382" *)
  wire _05931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6392" *)
  wire _05932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6402" *)
  wire _05933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6412" *)
  wire _05934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6422" *)
  wire _05935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6432" *)
  wire _05936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6442" *)
  wire _05937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6452" *)
  wire _05938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6462" *)
  wire _05939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6472" *)
  wire _05940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6482" *)
  wire _05941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6492" *)
  wire _05942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6502" *)
  wire _05943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6512" *)
  wire _05944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6522" *)
  wire _05945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6532" *)
  wire _05946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6542" *)
  wire _05947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6552" *)
  wire _05948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6562" *)
  wire _05949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6572" *)
  wire _05950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6582" *)
  wire _05951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6592" *)
  wire _05952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6602" *)
  wire _05953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6612" *)
  wire _05954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6622" *)
  wire _05955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6632" *)
  wire _05956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6642" *)
  wire _05957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6678" *)
  wire _05958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6708" *)
  wire _05959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6718" *)
  wire _05960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6728" *)
  wire _05961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6738" *)
  wire _05962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6748" *)
  wire _05963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6758" *)
  wire _05964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6768" *)
  wire _05965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6778" *)
  wire _05966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6788" *)
  wire _05967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6798" *)
  wire _05968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6808" *)
  wire _05969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6818" *)
  wire _05970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6828" *)
  wire _05971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6838" *)
  wire _05972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6848" *)
  wire _05973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6858" *)
  wire _05974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6868" *)
  wire _05975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6878" *)
  wire _05976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6888" *)
  wire _05977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6898" *)
  wire _05978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6908" *)
  wire _05979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6918" *)
  wire _05980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6928" *)
  wire _05981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6938" *)
  wire _05982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6948" *)
  wire _05983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6958" *)
  wire _05984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6968" *)
  wire _05985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6978" *)
  wire _05986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6988" *)
  wire _05987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6998" *)
  wire _05988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7008" *)
  wire _05989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7018" *)
  wire _05990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7028" *)
  wire _05991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7038" *)
  wire _05992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7048" *)
  wire _05993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7058" *)
  wire _05994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7068" *)
  wire _05995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7078" *)
  wire _05996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7088" *)
  wire _05997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7098" *)
  wire _05998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7108" *)
  wire _05999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7118" *)
  wire _06000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7128" *)
  wire _06001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7138" *)
  wire _06002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7148" *)
  wire _06003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7158" *)
  wire _06004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7168" *)
  wire _06005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7178" *)
  wire _06006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7188" *)
  wire _06007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7198" *)
  wire _06008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7208" *)
  wire _06009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7218" *)
  wire _06010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7228" *)
  wire _06011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7238" *)
  wire _06012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7248" *)
  wire _06013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7258" *)
  wire _06014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7268" *)
  wire _06015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7278" *)
  wire _06016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7288" *)
  wire _06017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7298" *)
  wire _06018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7308" *)
  wire _06019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7318" *)
  wire _06020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7328" *)
  wire _06021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7338" *)
  wire _06022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7348" *)
  wire _06023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7358" *)
  wire _06024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7368" *)
  wire _06025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7378" *)
  wire _06026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7388" *)
  wire _06027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7398" *)
  wire _06028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7408" *)
  wire _06029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7418" *)
  wire _06030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7428" *)
  wire _06031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7438" *)
  wire _06032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7448" *)
  wire _06033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7458" *)
  wire _06034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7468" *)
  wire _06035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7478" *)
  wire _06036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7488" *)
  wire _06037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7498" *)
  wire _06038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7508" *)
  wire _06039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7518" *)
  wire _06040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7528" *)
  wire _06041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7538" *)
  wire _06042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7548" *)
  wire _06043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7558" *)
  wire _06044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7568" *)
  wire _06045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7578" *)
  wire _06046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7588" *)
  wire _06047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7598" *)
  wire _06048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7608" *)
  wire _06049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7618" *)
  wire _06050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7628" *)
  wire _06051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7638" *)
  wire _06052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7648" *)
  wire _06053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7658" *)
  wire _06054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7668" *)
  wire _06055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7678" *)
  wire _06056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7688" *)
  wire _06057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7698" *)
  wire _06058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7708" *)
  wire _06059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7718" *)
  wire _06060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7728" *)
  wire _06061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7738" *)
  wire _06062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7748" *)
  wire _06063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7758" *)
  wire _06064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7768" *)
  wire _06065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7778" *)
  wire _06066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7788" *)
  wire _06067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7798" *)
  wire _06068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7808" *)
  wire _06069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7818" *)
  wire _06070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7828" *)
  wire _06071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7838" *)
  wire _06072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7848" *)
  wire _06073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7858" *)
  wire _06074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7868" *)
  wire _06075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7878" *)
  wire _06076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7888" *)
  wire _06077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7898" *)
  wire _06078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7908" *)
  wire _06079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7918" *)
  wire _06080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7928" *)
  wire _06081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7938" *)
  wire _06082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7948" *)
  wire _06083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7958" *)
  wire _06084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7968" *)
  wire _06085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7978" *)
  wire _06086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8014" *)
  wire _06087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8044" *)
  wire _06088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8054" *)
  wire _06089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8064" *)
  wire _06090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8074" *)
  wire _06091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8084" *)
  wire _06092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8094" *)
  wire _06093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8104" *)
  wire _06094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8114" *)
  wire _06095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8124" *)
  wire _06096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8134" *)
  wire _06097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8144" *)
  wire _06098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8154" *)
  wire _06099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8164" *)
  wire _06100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8174" *)
  wire _06101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8184" *)
  wire _06102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8194" *)
  wire _06103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8204" *)
  wire _06104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8214" *)
  wire _06105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8224" *)
  wire _06106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8234" *)
  wire _06107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8244" *)
  wire _06108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8254" *)
  wire _06109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8264" *)
  wire _06110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8274" *)
  wire _06111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8284" *)
  wire _06112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8294" *)
  wire _06113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8304" *)
  wire _06114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8314" *)
  wire _06115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8324" *)
  wire _06116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8334" *)
  wire _06117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8344" *)
  wire _06118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8354" *)
  wire _06119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8364" *)
  wire _06120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8374" *)
  wire _06121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8384" *)
  wire _06122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8394" *)
  wire _06123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8404" *)
  wire _06124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8414" *)
  wire _06125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8424" *)
  wire _06126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8434" *)
  wire _06127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8444" *)
  wire _06128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8454" *)
  wire _06129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8464" *)
  wire _06130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8474" *)
  wire _06131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8484" *)
  wire _06132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8494" *)
  wire _06133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8504" *)
  wire _06134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8514" *)
  wire _06135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8524" *)
  wire _06136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8534" *)
  wire _06137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8544" *)
  wire _06138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8554" *)
  wire _06139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8564" *)
  wire _06140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8574" *)
  wire _06141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8584" *)
  wire _06142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8594" *)
  wire _06143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8604" *)
  wire _06144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8614" *)
  wire _06145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8624" *)
  wire _06146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8634" *)
  wire _06147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8644" *)
  wire _06148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8654" *)
  wire _06149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8664" *)
  wire _06150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8674" *)
  wire _06151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8684" *)
  wire _06152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8694" *)
  wire _06153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8704" *)
  wire _06154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8714" *)
  wire _06155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8724" *)
  wire _06156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8734" *)
  wire _06157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8744" *)
  wire _06158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8754" *)
  wire _06159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8764" *)
  wire _06160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8774" *)
  wire _06161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8784" *)
  wire _06162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8794" *)
  wire _06163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8804" *)
  wire _06164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8814" *)
  wire _06165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8824" *)
  wire _06166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8834" *)
  wire _06167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8844" *)
  wire _06168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8854" *)
  wire _06169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8864" *)
  wire _06170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8874" *)
  wire _06171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8884" *)
  wire _06172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8894" *)
  wire _06173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8904" *)
  wire _06174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8914" *)
  wire _06175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8924" *)
  wire _06176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8934" *)
  wire _06177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8944" *)
  wire _06178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8954" *)
  wire _06179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8964" *)
  wire _06180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8974" *)
  wire _06181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8984" *)
  wire _06182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8994" *)
  wire _06183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9004" *)
  wire _06184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9014" *)
  wire _06185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9024" *)
  wire _06186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9034" *)
  wire _06187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9044" *)
  wire _06188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9054" *)
  wire _06189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9064" *)
  wire _06190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9074" *)
  wire _06191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9084" *)
  wire _06192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9094" *)
  wire _06193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9104" *)
  wire _06194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9114" *)
  wire _06195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9124" *)
  wire _06196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9134" *)
  wire _06197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9144" *)
  wire _06198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9154" *)
  wire _06199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9164" *)
  wire _06200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9174" *)
  wire _06201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9184" *)
  wire _06202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9194" *)
  wire _06203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9204" *)
  wire _06204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9214" *)
  wire _06205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9224" *)
  wire _06206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9234" *)
  wire _06207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9244" *)
  wire _06208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9254" *)
  wire _06209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9264" *)
  wire _06210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9274" *)
  wire _06211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9284" *)
  wire _06212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9294" *)
  wire _06213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9304" *)
  wire _06214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9314" *)
  wire _06215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9350" *)
  wire _06216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9380" *)
  wire _06217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9390" *)
  wire _06218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9400" *)
  wire _06219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9410" *)
  wire _06220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9420" *)
  wire _06221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9430" *)
  wire _06222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9440" *)
  wire _06223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9450" *)
  wire _06224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9460" *)
  wire _06225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9470" *)
  wire _06226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9480" *)
  wire _06227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9490" *)
  wire _06228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9500" *)
  wire _06229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9510" *)
  wire _06230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9520" *)
  wire _06231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9530" *)
  wire _06232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9540" *)
  wire _06233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9550" *)
  wire _06234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9560" *)
  wire _06235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9570" *)
  wire _06236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9580" *)
  wire _06237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9590" *)
  wire _06238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9600" *)
  wire _06239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9610" *)
  wire _06240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9620" *)
  wire _06241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9630" *)
  wire _06242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9640" *)
  wire _06243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9650" *)
  wire _06244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9660" *)
  wire _06245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9670" *)
  wire _06246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9680" *)
  wire _06247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9690" *)
  wire _06248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9700" *)
  wire _06249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9710" *)
  wire _06250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9720" *)
  wire _06251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9730" *)
  wire _06252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9740" *)
  wire _06253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9750" *)
  wire _06254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9760" *)
  wire _06255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9770" *)
  wire _06256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9780" *)
  wire _06257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9790" *)
  wire _06258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9800" *)
  wire _06259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9810" *)
  wire _06260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9820" *)
  wire _06261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9830" *)
  wire _06262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9840" *)
  wire _06263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9850" *)
  wire _06264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9860" *)
  wire _06265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9870" *)
  wire _06266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9880" *)
  wire _06267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9890" *)
  wire _06268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9900" *)
  wire _06269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9910" *)
  wire _06270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9920" *)
  wire _06271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9930" *)
  wire _06272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9940" *)
  wire _06273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9950" *)
  wire _06274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9960" *)
  wire _06275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9970" *)
  wire _06276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9980" *)
  wire _06277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9990" *)
  wire _06278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27872" *)
  wire [11:0] _06279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27881" *)
  wire [11:0] _06280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27890" *)
  wire [11:0] _06281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27899" *)
  wire [11:0] _06282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27908" *)
  wire [11:0] _06283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27917" *)
  wire [11:0] _06284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27926" *)
  wire [11:0] _06285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27935" *)
  wire [11:0] _06286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27944" *)
  wire [11:0] _06287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27953" *)
  wire [11:0] _06288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27962" *)
  wire [11:0] _06289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27971" *)
  wire [11:0] _06290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27980" *)
  wire [11:0] _06291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27989" *)
  wire [11:0] _06292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2799" *)
  wire [11:0] _06293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27998" *)
  wire [11:0] _06294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28007" *)
  wire [11:0] _06295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28016" *)
  wire [11:0] _06296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28025" *)
  wire [11:0] _06297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28034" *)
  wire [11:0] _06298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28043" *)
  wire [11:0] _06299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28052" *)
  wire [11:0] _06300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28061" *)
  wire [11:0] _06301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28070" *)
  wire [11:0] _06302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28079" *)
  wire [11:0] _06303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2808" *)
  wire [11:0] _06304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28088" *)
  wire [11:0] _06305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28097" *)
  wire [11:0] _06306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28106" *)
  wire [11:0] _06307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28115" *)
  wire [11:0] _06308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28124" *)
  wire [11:0] _06309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28133" *)
  wire [11:0] _06310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28142" *)
  wire [11:0] _06311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28151" *)
  wire [11:0] _06312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28160" *)
  wire [11:0] _06313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28169" *)
  wire [11:0] _06314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2817" *)
  wire [11:0] _06315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28178" *)
  wire [11:0] _06316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28187" *)
  wire [11:0] _06317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28196" *)
  wire [11:0] _06318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28205" *)
  wire [11:0] _06319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28214" *)
  wire [11:0] _06320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28223" *)
  wire [11:0] _06321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28232" *)
  wire [11:0] _06322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28241" *)
  wire [11:0] _06323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28250" *)
  wire [11:0] _06324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28259" *)
  wire [11:0] _06325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2826" *)
  wire [11:0] _06326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28268" *)
  wire [11:0] _06327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28277" *)
  wire [11:0] _06328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28286" *)
  wire [11:0] _06329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28295" *)
  wire [11:0] _06330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28304" *)
  wire [11:0] _06331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28313" *)
  wire [11:0] _06332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28322" *)
  wire [11:0] _06333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28331" *)
  wire [11:0] _06334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28340" *)
  wire [11:0] _06335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28349" *)
  wire [11:0] _06336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2835" *)
  wire [11:0] _06337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28358" *)
  wire [11:0] _06338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28367" *)
  wire [11:0] _06339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28376" *)
  wire [11:0] _06340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28385" *)
  wire [11:0] _06341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28394" *)
  wire [11:0] _06342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28403" *)
  wire [11:0] _06343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28412" *)
  wire [11:0] _06344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28421" *)
  wire [11:0] _06345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28430" *)
  wire [11:0] _06346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28439" *)
  wire [11:0] _06347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2844" *)
  wire [11:0] _06348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2853" *)
  wire [11:0] _06349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2862" *)
  wire [11:0] _06350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2871" *)
  wire [11:0] _06351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2880" *)
  wire [11:0] _06352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2889" *)
  wire [11:0] _06353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2898" *)
  wire [11:0] _06354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2907" *)
  wire [11:0] _06355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2916" *)
  wire [11:0] _06356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2925" *)
  wire [11:0] _06357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2934" *)
  wire [11:0] _06358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2943" *)
  wire [11:0] _06359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2952" *)
  wire [11:0] _06360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2961" *)
  wire [11:0] _06361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2970" *)
  wire [11:0] _06362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2979" *)
  wire [11:0] _06363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2988" *)
  wire [11:0] _06364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2997" *)
  wire [11:0] _06365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3006" *)
  wire [11:0] _06366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3015" *)
  wire [11:0] _06367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3024" *)
  wire [11:0] _06368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3033" *)
  wire [11:0] _06369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3042" *)
  wire [11:0] _06370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3051" *)
  wire [11:0] _06371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3060" *)
  wire [11:0] _06372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3069" *)
  wire [11:0] _06373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3078" *)
  wire [11:0] _06374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3087" *)
  wire [11:0] _06375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3096" *)
  wire [11:0] _06376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3105" *)
  wire [11:0] _06377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3114" *)
  wire [11:0] _06378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3123" *)
  wire [11:0] _06379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3132" *)
  wire [11:0] _06380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3141" *)
  wire [11:0] _06381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3150" *)
  wire [11:0] _06382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3159" *)
  wire [11:0] _06383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3168" *)
  wire [11:0] _06384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3177" *)
  wire [11:0] _06385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3186" *)
  wire [11:0] _06386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3195" *)
  wire [11:0] _06387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3204" *)
  wire [11:0] _06388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3213" *)
  wire [11:0] _06389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3222" *)
  wire [11:0] _06390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3231" *)
  wire [11:0] _06391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3240" *)
  wire [11:0] _06392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3249" *)
  wire [11:0] _06393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3258" *)
  wire [11:0] _06394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3267" *)
  wire [11:0] _06395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3276" *)
  wire [11:0] _06396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3285" *)
  wire [11:0] _06397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3294" *)
  wire [11:0] _06398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3303" *)
  wire [11:0] _06399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3312" *)
  wire [11:0] _06400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3321" *)
  wire [11:0] _06401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3330" *)
  wire [11:0] _06402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3339" *)
  wire [11:0] _06403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3348" *)
  wire [11:0] _06404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3357" *)
  wire [11:0] _06405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3366" *)
  wire [11:0] _06406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29041" *)
  wire _06407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3968" *)
  wire _06408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10000" *)
  wire _06409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10010" *)
  wire _06410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10020" *)
  wire _06411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10030" *)
  wire _06412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10040" *)
  wire _06413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10050" *)
  wire _06414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10060" *)
  wire _06415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10070" *)
  wire _06416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10080" *)
  wire _06417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10090" *)
  wire _06418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10100" *)
  wire _06419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10110" *)
  wire _06420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10120" *)
  wire _06421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10130" *)
  wire _06422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10140" *)
  wire _06423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10150" *)
  wire _06424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10160" *)
  wire _06425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10170" *)
  wire _06426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10180" *)
  wire _06427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10190" *)
  wire _06428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10200" *)
  wire _06429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10210" *)
  wire _06430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10220" *)
  wire _06431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10230" *)
  wire _06432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10240" *)
  wire _06433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10250" *)
  wire _06434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10260" *)
  wire _06435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10270" *)
  wire _06436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10280" *)
  wire _06437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10290" *)
  wire _06438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10300" *)
  wire _06439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10310" *)
  wire _06440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10320" *)
  wire _06441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10330" *)
  wire _06442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10340" *)
  wire _06443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10350" *)
  wire _06444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10360" *)
  wire _06445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10370" *)
  wire _06446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10380" *)
  wire _06447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10390" *)
  wire _06448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10400" *)
  wire _06449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10410" *)
  wire _06450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10420" *)
  wire _06451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10430" *)
  wire _06452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10440" *)
  wire _06453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10450" *)
  wire _06454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10460" *)
  wire _06455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10470" *)
  wire _06456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10480" *)
  wire _06457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10490" *)
  wire _06458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10500" *)
  wire _06459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10510" *)
  wire _06460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10520" *)
  wire _06461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10530" *)
  wire _06462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10540" *)
  wire _06463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10550" *)
  wire _06464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10560" *)
  wire _06465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10570" *)
  wire _06466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10580" *)
  wire _06467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10590" *)
  wire _06468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10600" *)
  wire _06469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10610" *)
  wire _06470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10620" *)
  wire _06471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10630" *)
  wire _06472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10640" *)
  wire _06473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10650" *)
  wire _06474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10716" *)
  wire _06475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10726" *)
  wire _06476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10736" *)
  wire _06477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10746" *)
  wire _06478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10756" *)
  wire _06479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10766" *)
  wire _06480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10776" *)
  wire _06481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10786" *)
  wire _06482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10796" *)
  wire _06483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10806" *)
  wire _06484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10816" *)
  wire _06485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10826" *)
  wire _06486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10836" *)
  wire _06487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10846" *)
  wire _06488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10856" *)
  wire _06489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10866" *)
  wire _06490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10876" *)
  wire _06491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10886" *)
  wire _06492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10896" *)
  wire _06493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10906" *)
  wire _06494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10916" *)
  wire _06495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10926" *)
  wire _06496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10936" *)
  wire _06497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10946" *)
  wire _06498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10956" *)
  wire _06499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10966" *)
  wire _06500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10976" *)
  wire _06501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10986" *)
  wire _06502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10996" *)
  wire _06503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11006" *)
  wire _06504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11016" *)
  wire _06505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11026" *)
  wire _06506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11036" *)
  wire _06507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11046" *)
  wire _06508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11056" *)
  wire _06509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11066" *)
  wire _06510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11076" *)
  wire _06511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11086" *)
  wire _06512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11096" *)
  wire _06513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11106" *)
  wire _06514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11116" *)
  wire _06515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11126" *)
  wire _06516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11136" *)
  wire _06517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11146" *)
  wire _06518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11156" *)
  wire _06519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11166" *)
  wire _06520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11176" *)
  wire _06521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11186" *)
  wire _06522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11196" *)
  wire _06523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11206" *)
  wire _06524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11216" *)
  wire _06525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11226" *)
  wire _06526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11236" *)
  wire _06527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11246" *)
  wire _06528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11256" *)
  wire _06529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11266" *)
  wire _06530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11276" *)
  wire _06531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11286" *)
  wire _06532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11296" *)
  wire _06533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11306" *)
  wire _06534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11316" *)
  wire _06535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11326" *)
  wire _06536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16049" *)
  wire _06537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16059" *)
  wire _06538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16069" *)
  wire _06539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16079" *)
  wire _06540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16089" *)
  wire _06541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16099" *)
  wire _06542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16109" *)
  wire _06543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16119" *)
  wire _06544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16129" *)
  wire _06545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16139" *)
  wire _06546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16149" *)
  wire _06547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16159" *)
  wire _06548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16169" *)
  wire _06549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16179" *)
  wire _06550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16189" *)
  wire _06551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16199" *)
  wire _06552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16209" *)
  wire _06553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16219" *)
  wire _06554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16229" *)
  wire _06555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16239" *)
  wire _06556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16249" *)
  wire _06557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16259" *)
  wire _06558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16269" *)
  wire _06559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16279" *)
  wire _06560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16289" *)
  wire _06561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16299" *)
  wire _06562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16309" *)
  wire _06563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16319" *)
  wire _06564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16329" *)
  wire _06565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16339" *)
  wire _06566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16349" *)
  wire _06567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16359" *)
  wire _06568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16369" *)
  wire _06569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16379" *)
  wire _06570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16389" *)
  wire _06571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16399" *)
  wire _06572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16409" *)
  wire _06573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16419" *)
  wire _06574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16429" *)
  wire _06575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16439" *)
  wire _06576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16449" *)
  wire _06577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16459" *)
  wire _06578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16469" *)
  wire _06579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16479" *)
  wire _06580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16489" *)
  wire _06581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16499" *)
  wire _06582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16509" *)
  wire _06583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16519" *)
  wire _06584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16529" *)
  wire _06585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16539" *)
  wire _06586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16549" *)
  wire _06587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16559" *)
  wire _06588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16569" *)
  wire _06589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16579" *)
  wire _06590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16589" *)
  wire _06591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16599" *)
  wire _06592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16609" *)
  wire _06593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16619" *)
  wire _06594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16629" *)
  wire _06595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16639" *)
  wire _06596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16649" *)
  wire _06597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16659" *)
  wire _06598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16669" *)
  wire _06599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16679" *)
  wire _06600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16689" *)
  wire _06601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16699" *)
  wire _06602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16709" *)
  wire _06603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16719" *)
  wire _06604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16729" *)
  wire _06605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16739" *)
  wire _06606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16749" *)
  wire _06607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16759" *)
  wire _06608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16769" *)
  wire _06609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16779" *)
  wire _06610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16789" *)
  wire _06611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16799" *)
  wire _06612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16809" *)
  wire _06613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16819" *)
  wire _06614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16829" *)
  wire _06615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16839" *)
  wire _06616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16849" *)
  wire _06617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16859" *)
  wire _06618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16869" *)
  wire _06619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16879" *)
  wire _06620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16889" *)
  wire _06621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16899" *)
  wire _06622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16909" *)
  wire _06623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16919" *)
  wire _06624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16929" *)
  wire _06625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16939" *)
  wire _06626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16949" *)
  wire _06627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16959" *)
  wire _06628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16969" *)
  wire _06629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16979" *)
  wire _06630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16989" *)
  wire _06631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16999" *)
  wire _06632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17009" *)
  wire _06633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17019" *)
  wire _06634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17029" *)
  wire _06635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17039" *)
  wire _06636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17049" *)
  wire _06637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17059" *)
  wire _06638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17069" *)
  wire _06639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17079" *)
  wire _06640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17089" *)
  wire _06641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17099" *)
  wire _06642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17109" *)
  wire _06643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17119" *)
  wire _06644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17129" *)
  wire _06645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17139" *)
  wire _06646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17149" *)
  wire _06647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17159" *)
  wire _06648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17169" *)
  wire _06649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17179" *)
  wire _06650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17189" *)
  wire _06651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17199" *)
  wire _06652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17209" *)
  wire _06653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17219" *)
  wire _06654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17229" *)
  wire _06655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17239" *)
  wire _06656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17249" *)
  wire _06657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17259" *)
  wire _06658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17269" *)
  wire _06659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17279" *)
  wire _06660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17289" *)
  wire _06661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17299" *)
  wire _06662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17309" *)
  wire _06663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17319" *)
  wire _06664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17373" *)
  wire _06665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17383" *)
  wire _06666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17393" *)
  wire _06667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17403" *)
  wire _06668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17413" *)
  wire _06669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17423" *)
  wire _06670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17433" *)
  wire _06671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17443" *)
  wire _06672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17453" *)
  wire _06673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17463" *)
  wire _06674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17473" *)
  wire _06675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17483" *)
  wire _06676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17493" *)
  wire _06677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17503" *)
  wire _06678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17513" *)
  wire _06679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17523" *)
  wire _06680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17533" *)
  wire _06681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17543" *)
  wire _06682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17553" *)
  wire _06683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17563" *)
  wire _06684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17573" *)
  wire _06685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17583" *)
  wire _06686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17593" *)
  wire _06687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17603" *)
  wire _06688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17613" *)
  wire _06689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17623" *)
  wire _06690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17633" *)
  wire _06691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17643" *)
  wire _06692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17653" *)
  wire _06693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17663" *)
  wire _06694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17673" *)
  wire _06695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17683" *)
  wire _06696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17693" *)
  wire _06697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17703" *)
  wire _06698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17713" *)
  wire _06699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17723" *)
  wire _06700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17733" *)
  wire _06701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17743" *)
  wire _06702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17753" *)
  wire _06703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17763" *)
  wire _06704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17773" *)
  wire _06705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17783" *)
  wire _06706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17793" *)
  wire _06707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17803" *)
  wire _06708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17813" *)
  wire _06709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17823" *)
  wire _06710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17833" *)
  wire _06711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17843" *)
  wire _06712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17853" *)
  wire _06713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17863" *)
  wire _06714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17873" *)
  wire _06715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17883" *)
  wire _06716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17893" *)
  wire _06717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17903" *)
  wire _06718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17913" *)
  wire _06719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17923" *)
  wire _06720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17933" *)
  wire _06721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17943" *)
  wire _06722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17953" *)
  wire _06723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17963" *)
  wire _06724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17973" *)
  wire _06725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17983" *)
  wire _06726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17993" *)
  wire _06727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18003" *)
  wire _06728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18013" *)
  wire _06729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18023" *)
  wire _06730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18033" *)
  wire _06731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18043" *)
  wire _06732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18053" *)
  wire _06733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18063" *)
  wire _06734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18073" *)
  wire _06735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18083" *)
  wire _06736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18093" *)
  wire _06737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18103" *)
  wire _06738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18113" *)
  wire _06739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18123" *)
  wire _06740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18133" *)
  wire _06741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18143" *)
  wire _06742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18153" *)
  wire _06743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18163" *)
  wire _06744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18173" *)
  wire _06745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18183" *)
  wire _06746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18193" *)
  wire _06747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18203" *)
  wire _06748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18213" *)
  wire _06749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18223" *)
  wire _06750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18233" *)
  wire _06751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18243" *)
  wire _06752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18253" *)
  wire _06753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18263" *)
  wire _06754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18273" *)
  wire _06755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18283" *)
  wire _06756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18293" *)
  wire _06757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18303" *)
  wire _06758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18313" *)
  wire _06759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18323" *)
  wire _06760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18333" *)
  wire _06761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18343" *)
  wire _06762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18353" *)
  wire _06763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18363" *)
  wire _06764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18373" *)
  wire _06765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18383" *)
  wire _06766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18393" *)
  wire _06767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18403" *)
  wire _06768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18413" *)
  wire _06769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18423" *)
  wire _06770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18433" *)
  wire _06771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18443" *)
  wire _06772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18453" *)
  wire _06773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18463" *)
  wire _06774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18473" *)
  wire _06775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18483" *)
  wire _06776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18493" *)
  wire _06777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18503" *)
  wire _06778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18513" *)
  wire _06779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18523" *)
  wire _06780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18533" *)
  wire _06781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18543" *)
  wire _06782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18553" *)
  wire _06783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18563" *)
  wire _06784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18573" *)
  wire _06785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18583" *)
  wire _06786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18593" *)
  wire _06787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18603" *)
  wire _06788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18613" *)
  wire _06789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18623" *)
  wire _06790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18633" *)
  wire _06791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18643" *)
  wire _06792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18697" *)
  wire _06793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18707" *)
  wire _06794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18717" *)
  wire _06795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18727" *)
  wire _06796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18737" *)
  wire _06797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18747" *)
  wire _06798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18757" *)
  wire _06799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18767" *)
  wire _06800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18777" *)
  wire _06801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18787" *)
  wire _06802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18797" *)
  wire _06803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18807" *)
  wire _06804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18817" *)
  wire _06805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18827" *)
  wire _06806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18837" *)
  wire _06807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18847" *)
  wire _06808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18857" *)
  wire _06809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18867" *)
  wire _06810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18877" *)
  wire _06811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18887" *)
  wire _06812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18897" *)
  wire _06813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18907" *)
  wire _06814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18917" *)
  wire _06815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18927" *)
  wire _06816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18937" *)
  wire _06817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18947" *)
  wire _06818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18957" *)
  wire _06819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18967" *)
  wire _06820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18977" *)
  wire _06821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18987" *)
  wire _06822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18997" *)
  wire _06823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19007" *)
  wire _06824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19017" *)
  wire _06825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19027" *)
  wire _06826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19037" *)
  wire _06827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19047" *)
  wire _06828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19057" *)
  wire _06829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19067" *)
  wire _06830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19077" *)
  wire _06831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19087" *)
  wire _06832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19097" *)
  wire _06833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19107" *)
  wire _06834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19117" *)
  wire _06835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19127" *)
  wire _06836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19137" *)
  wire _06837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19147" *)
  wire _06838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19157" *)
  wire _06839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19167" *)
  wire _06840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19177" *)
  wire _06841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19187" *)
  wire _06842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19197" *)
  wire _06843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19207" *)
  wire _06844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19217" *)
  wire _06845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19227" *)
  wire _06846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19237" *)
  wire _06847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19247" *)
  wire _06848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19257" *)
  wire _06849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19267" *)
  wire _06850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19277" *)
  wire _06851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19287" *)
  wire _06852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19297" *)
  wire _06853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19307" *)
  wire _06854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19317" *)
  wire _06855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19327" *)
  wire _06856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19337" *)
  wire _06857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19347" *)
  wire _06858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19357" *)
  wire _06859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19367" *)
  wire _06860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19377" *)
  wire _06861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19387" *)
  wire _06862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19397" *)
  wire _06863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19407" *)
  wire _06864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19417" *)
  wire _06865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19427" *)
  wire _06866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19437" *)
  wire _06867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19447" *)
  wire _06868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19457" *)
  wire _06869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19467" *)
  wire _06870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19477" *)
  wire _06871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19487" *)
  wire _06872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19497" *)
  wire _06873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19507" *)
  wire _06874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19517" *)
  wire _06875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19527" *)
  wire _06876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19537" *)
  wire _06877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19547" *)
  wire _06878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19557" *)
  wire _06879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19567" *)
  wire _06880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19577" *)
  wire _06881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19587" *)
  wire _06882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19597" *)
  wire _06883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19607" *)
  wire _06884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19617" *)
  wire _06885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19627" *)
  wire _06886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19637" *)
  wire _06887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19647" *)
  wire _06888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19657" *)
  wire _06889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19667" *)
  wire _06890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19677" *)
  wire _06891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19687" *)
  wire _06892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19697" *)
  wire _06893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19707" *)
  wire _06894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19717" *)
  wire _06895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19727" *)
  wire _06896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19737" *)
  wire _06897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19747" *)
  wire _06898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19757" *)
  wire _06899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19767" *)
  wire _06900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19777" *)
  wire _06901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19787" *)
  wire _06902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19797" *)
  wire _06903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19807" *)
  wire _06904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19817" *)
  wire _06905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19827" *)
  wire _06906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19837" *)
  wire _06907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19847" *)
  wire _06908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19857" *)
  wire _06909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19867" *)
  wire _06910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19877" *)
  wire _06911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19887" *)
  wire _06912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19897" *)
  wire _06913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19907" *)
  wire _06914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19917" *)
  wire _06915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19927" *)
  wire _06916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19937" *)
  wire _06917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19947" *)
  wire _06918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19957" *)
  wire _06919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19967" *)
  wire _06920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20021" *)
  wire _06921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20031" *)
  wire _06922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20041" *)
  wire _06923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20051" *)
  wire _06924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20061" *)
  wire _06925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20071" *)
  wire _06926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20081" *)
  wire _06927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20091" *)
  wire _06928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20101" *)
  wire _06929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20111" *)
  wire _06930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20121" *)
  wire _06931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20131" *)
  wire _06932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20141" *)
  wire _06933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20151" *)
  wire _06934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20161" *)
  wire _06935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20171" *)
  wire _06936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20181" *)
  wire _06937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20191" *)
  wire _06938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20201" *)
  wire _06939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20211" *)
  wire _06940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20221" *)
  wire _06941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20231" *)
  wire _06942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20241" *)
  wire _06943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20251" *)
  wire _06944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20261" *)
  wire _06945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20271" *)
  wire _06946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20281" *)
  wire _06947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20291" *)
  wire _06948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20301" *)
  wire _06949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20311" *)
  wire _06950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20321" *)
  wire _06951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20331" *)
  wire _06952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20341" *)
  wire _06953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20351" *)
  wire _06954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20361" *)
  wire _06955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20371" *)
  wire _06956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20381" *)
  wire _06957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20391" *)
  wire _06958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20401" *)
  wire _06959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20411" *)
  wire _06960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20421" *)
  wire _06961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20431" *)
  wire _06962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20441" *)
  wire _06963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20451" *)
  wire _06964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20461" *)
  wire _06965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20471" *)
  wire _06966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20481" *)
  wire _06967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20491" *)
  wire _06968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20501" *)
  wire _06969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20511" *)
  wire _06970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20521" *)
  wire _06971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20531" *)
  wire _06972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20541" *)
  wire _06973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20551" *)
  wire _06974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20561" *)
  wire _06975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20571" *)
  wire _06976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20581" *)
  wire _06977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20591" *)
  wire _06978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20601" *)
  wire _06979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20611" *)
  wire _06980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20621" *)
  wire _06981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20631" *)
  wire _06982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20641" *)
  wire _06983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20651" *)
  wire _06984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20661" *)
  wire _06985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20671" *)
  wire _06986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20681" *)
  wire _06987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20691" *)
  wire _06988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20701" *)
  wire _06989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20711" *)
  wire _06990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20721" *)
  wire _06991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20731" *)
  wire _06992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20741" *)
  wire _06993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20751" *)
  wire _06994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20761" *)
  wire _06995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20771" *)
  wire _06996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20781" *)
  wire _06997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20791" *)
  wire _06998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20801" *)
  wire _06999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20811" *)
  wire _07000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20821" *)
  wire _07001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20831" *)
  wire _07002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20841" *)
  wire _07003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20851" *)
  wire _07004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20861" *)
  wire _07005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20871" *)
  wire _07006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20881" *)
  wire _07007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20891" *)
  wire _07008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20901" *)
  wire _07009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20911" *)
  wire _07010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20921" *)
  wire _07011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20931" *)
  wire _07012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20941" *)
  wire _07013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20951" *)
  wire _07014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20961" *)
  wire _07015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20971" *)
  wire _07016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20981" *)
  wire _07017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20991" *)
  wire _07018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21001" *)
  wire _07019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21011" *)
  wire _07020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21021" *)
  wire _07021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21031" *)
  wire _07022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21041" *)
  wire _07023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21051" *)
  wire _07024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21061" *)
  wire _07025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21071" *)
  wire _07026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21081" *)
  wire _07027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21091" *)
  wire _07028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21101" *)
  wire _07029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21111" *)
  wire _07030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21121" *)
  wire _07031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21131" *)
  wire _07032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21141" *)
  wire _07033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21151" *)
  wire _07034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21161" *)
  wire _07035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21171" *)
  wire _07036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21181" *)
  wire _07037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21191" *)
  wire _07038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21201" *)
  wire _07039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21211" *)
  wire _07040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21221" *)
  wire _07041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21231" *)
  wire _07042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21241" *)
  wire _07043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21251" *)
  wire _07044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21261" *)
  wire _07045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21271" *)
  wire _07046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21281" *)
  wire _07047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21291" *)
  wire _07048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21345" *)
  wire _07049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21355" *)
  wire _07050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21365" *)
  wire _07051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21375" *)
  wire _07052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21385" *)
  wire _07053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21395" *)
  wire _07054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21405" *)
  wire _07055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21415" *)
  wire _07056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21425" *)
  wire _07057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21435" *)
  wire _07058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21445" *)
  wire _07059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21455" *)
  wire _07060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21465" *)
  wire _07061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21475" *)
  wire _07062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21485" *)
  wire _07063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21495" *)
  wire _07064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21505" *)
  wire _07065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21515" *)
  wire _07066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21525" *)
  wire _07067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21535" *)
  wire _07068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21545" *)
  wire _07069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21555" *)
  wire _07070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21565" *)
  wire _07071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21575" *)
  wire _07072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21585" *)
  wire _07073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21595" *)
  wire _07074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21605" *)
  wire _07075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21615" *)
  wire _07076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21625" *)
  wire _07077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21635" *)
  wire _07078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21645" *)
  wire _07079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21655" *)
  wire _07080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21665" *)
  wire _07081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21675" *)
  wire _07082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21685" *)
  wire _07083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21695" *)
  wire _07084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21705" *)
  wire _07085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21715" *)
  wire _07086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21725" *)
  wire _07087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21735" *)
  wire _07088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21745" *)
  wire _07089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21755" *)
  wire _07090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21765" *)
  wire _07091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21775" *)
  wire _07092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21785" *)
  wire _07093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21795" *)
  wire _07094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21805" *)
  wire _07095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21815" *)
  wire _07096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21825" *)
  wire _07097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21835" *)
  wire _07098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21845" *)
  wire _07099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21855" *)
  wire _07100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21865" *)
  wire _07101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21875" *)
  wire _07102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21885" *)
  wire _07103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21895" *)
  wire _07104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21905" *)
  wire _07105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21915" *)
  wire _07106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21925" *)
  wire _07107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21935" *)
  wire _07108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21945" *)
  wire _07109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21955" *)
  wire _07110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21965" *)
  wire _07111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21975" *)
  wire _07112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21985" *)
  wire _07113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21995" *)
  wire _07114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22005" *)
  wire _07115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22015" *)
  wire _07116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22025" *)
  wire _07117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22035" *)
  wire _07118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22045" *)
  wire _07119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22055" *)
  wire _07120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22065" *)
  wire _07121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22075" *)
  wire _07122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22085" *)
  wire _07123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22095" *)
  wire _07124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22105" *)
  wire _07125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22115" *)
  wire _07126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22125" *)
  wire _07127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22135" *)
  wire _07128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22145" *)
  wire _07129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22155" *)
  wire _07130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22165" *)
  wire _07131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22175" *)
  wire _07132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22185" *)
  wire _07133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22195" *)
  wire _07134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22205" *)
  wire _07135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22215" *)
  wire _07136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22225" *)
  wire _07137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22235" *)
  wire _07138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22245" *)
  wire _07139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22255" *)
  wire _07140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22265" *)
  wire _07141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22275" *)
  wire _07142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22285" *)
  wire _07143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22295" *)
  wire _07144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22305" *)
  wire _07145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22315" *)
  wire _07146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22325" *)
  wire _07147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22335" *)
  wire _07148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22345" *)
  wire _07149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22355" *)
  wire _07150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22365" *)
  wire _07151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22375" *)
  wire _07152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22385" *)
  wire _07153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22395" *)
  wire _07154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22405" *)
  wire _07155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22415" *)
  wire _07156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22425" *)
  wire _07157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22435" *)
  wire _07158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22445" *)
  wire _07159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22455" *)
  wire _07160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22465" *)
  wire _07161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22475" *)
  wire _07162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22485" *)
  wire _07163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22495" *)
  wire _07164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22505" *)
  wire _07165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22515" *)
  wire _07166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22525" *)
  wire _07167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22535" *)
  wire _07168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22545" *)
  wire _07169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22555" *)
  wire _07170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22565" *)
  wire _07171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22575" *)
  wire _07172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22585" *)
  wire _07173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22595" *)
  wire _07174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22605" *)
  wire _07175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22615" *)
  wire _07176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22669" *)
  wire _07177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22679" *)
  wire _07178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22689" *)
  wire _07179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22699" *)
  wire _07180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22709" *)
  wire _07181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22719" *)
  wire _07182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22729" *)
  wire _07183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22739" *)
  wire _07184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22749" *)
  wire _07185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22759" *)
  wire _07186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22769" *)
  wire _07187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22779" *)
  wire _07188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22789" *)
  wire _07189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22799" *)
  wire _07190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22809" *)
  wire _07191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22819" *)
  wire _07192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22829" *)
  wire _07193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22839" *)
  wire _07194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22849" *)
  wire _07195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22859" *)
  wire _07196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22869" *)
  wire _07197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22879" *)
  wire _07198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22889" *)
  wire _07199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22899" *)
  wire _07200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22909" *)
  wire _07201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22919" *)
  wire _07202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22929" *)
  wire _07203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22939" *)
  wire _07204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22949" *)
  wire _07205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22959" *)
  wire _07206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22969" *)
  wire _07207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22979" *)
  wire _07208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22989" *)
  wire _07209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22999" *)
  wire _07210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23009" *)
  wire _07211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23019" *)
  wire _07212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23029" *)
  wire _07213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23039" *)
  wire _07214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23049" *)
  wire _07215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23059" *)
  wire _07216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23069" *)
  wire _07217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23079" *)
  wire _07218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23089" *)
  wire _07219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23099" *)
  wire _07220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23109" *)
  wire _07221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23119" *)
  wire _07222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23129" *)
  wire _07223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23139" *)
  wire _07224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23149" *)
  wire _07225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23159" *)
  wire _07226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23169" *)
  wire _07227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23179" *)
  wire _07228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23189" *)
  wire _07229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23199" *)
  wire _07230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23209" *)
  wire _07231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23219" *)
  wire _07232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23229" *)
  wire _07233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23239" *)
  wire _07234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23249" *)
  wire _07235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23259" *)
  wire _07236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23269" *)
  wire _07237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23279" *)
  wire _07238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23289" *)
  wire _07239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23299" *)
  wire _07240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23309" *)
  wire _07241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23319" *)
  wire _07242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23329" *)
  wire _07243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23339" *)
  wire _07244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23349" *)
  wire _07245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23359" *)
  wire _07246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23369" *)
  wire _07247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23379" *)
  wire _07248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23389" *)
  wire _07249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23399" *)
  wire _07250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23409" *)
  wire _07251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23419" *)
  wire _07252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23429" *)
  wire _07253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23439" *)
  wire _07254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23449" *)
  wire _07255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23459" *)
  wire _07256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23469" *)
  wire _07257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23479" *)
  wire _07258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23489" *)
  wire _07259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23499" *)
  wire _07260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23509" *)
  wire _07261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23519" *)
  wire _07262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23529" *)
  wire _07263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23539" *)
  wire _07264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23549" *)
  wire _07265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23559" *)
  wire _07266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23569" *)
  wire _07267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23579" *)
  wire _07268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23589" *)
  wire _07269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23599" *)
  wire _07270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23609" *)
  wire _07271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23619" *)
  wire _07272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23629" *)
  wire _07273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23639" *)
  wire _07274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23649" *)
  wire _07275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23659" *)
  wire _07276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23669" *)
  wire _07277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23679" *)
  wire _07278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23689" *)
  wire _07279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23699" *)
  wire _07280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23709" *)
  wire _07281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23719" *)
  wire _07282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23729" *)
  wire _07283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23739" *)
  wire _07284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23749" *)
  wire _07285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23759" *)
  wire _07286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23769" *)
  wire _07287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23779" *)
  wire _07288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23789" *)
  wire _07289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23799" *)
  wire _07290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23809" *)
  wire _07291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23819" *)
  wire _07292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23829" *)
  wire _07293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23839" *)
  wire _07294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23849" *)
  wire _07295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23859" *)
  wire _07296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23869" *)
  wire _07297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23879" *)
  wire _07298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23889" *)
  wire _07299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23899" *)
  wire _07300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23909" *)
  wire _07301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23919" *)
  wire _07302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23929" *)
  wire _07303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23939" *)
  wire _07304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23993" *)
  wire _07305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24003" *)
  wire _07306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24013" *)
  wire _07307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24023" *)
  wire _07308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24033" *)
  wire _07309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24043" *)
  wire _07310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24053" *)
  wire _07311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24063" *)
  wire _07312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24073" *)
  wire _07313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24083" *)
  wire _07314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24093" *)
  wire _07315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24103" *)
  wire _07316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24113" *)
  wire _07317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24123" *)
  wire _07318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24133" *)
  wire _07319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24143" *)
  wire _07320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24153" *)
  wire _07321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24163" *)
  wire _07322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24173" *)
  wire _07323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24183" *)
  wire _07324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24193" *)
  wire _07325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24203" *)
  wire _07326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24213" *)
  wire _07327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24223" *)
  wire _07328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24233" *)
  wire _07329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24243" *)
  wire _07330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24253" *)
  wire _07331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24263" *)
  wire _07332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24273" *)
  wire _07333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24283" *)
  wire _07334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24293" *)
  wire _07335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24303" *)
  wire _07336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24313" *)
  wire _07337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24323" *)
  wire _07338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24333" *)
  wire _07339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24343" *)
  wire _07340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24353" *)
  wire _07341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24363" *)
  wire _07342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24373" *)
  wire _07343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24383" *)
  wire _07344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24393" *)
  wire _07345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24403" *)
  wire _07346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24413" *)
  wire _07347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24423" *)
  wire _07348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24433" *)
  wire _07349_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24443" *)
  wire _07350_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24453" *)
  wire _07351_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24463" *)
  wire _07352_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24473" *)
  wire _07353_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24483" *)
  wire _07354_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24493" *)
  wire _07355_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24503" *)
  wire _07356_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24513" *)
  wire _07357_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24523" *)
  wire _07358_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24533" *)
  wire _07359_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24543" *)
  wire _07360_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24553" *)
  wire _07361_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24563" *)
  wire _07362_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24573" *)
  wire _07363_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24583" *)
  wire _07364_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24593" *)
  wire _07365_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24603" *)
  wire _07366_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24613" *)
  wire _07367_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24623" *)
  wire _07368_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24633" *)
  wire _07369_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24643" *)
  wire _07370_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24653" *)
  wire _07371_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24663" *)
  wire _07372_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24673" *)
  wire _07373_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24683" *)
  wire _07374_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24693" *)
  wire _07375_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24703" *)
  wire _07376_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24713" *)
  wire _07377_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24723" *)
  wire _07378_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24733" *)
  wire _07379_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24743" *)
  wire _07380_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24753" *)
  wire _07381_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24763" *)
  wire _07382_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24773" *)
  wire _07383_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24783" *)
  wire _07384_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24793" *)
  wire _07385_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24803" *)
  wire _07386_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24813" *)
  wire _07387_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24823" *)
  wire _07388_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24833" *)
  wire _07389_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24843" *)
  wire _07390_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24853" *)
  wire _07391_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24863" *)
  wire _07392_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24873" *)
  wire _07393_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24883" *)
  wire _07394_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24893" *)
  wire _07395_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24903" *)
  wire _07396_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24913" *)
  wire _07397_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24923" *)
  wire _07398_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24933" *)
  wire _07399_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24943" *)
  wire _07400_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24953" *)
  wire _07401_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24963" *)
  wire _07402_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24973" *)
  wire _07403_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24983" *)
  wire _07404_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24993" *)
  wire _07405_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25003" *)
  wire _07406_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25013" *)
  wire _07407_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25023" *)
  wire _07408_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25033" *)
  wire _07409_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25043" *)
  wire _07410_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25053" *)
  wire _07411_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25063" *)
  wire _07412_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25073" *)
  wire _07413_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25083" *)
  wire _07414_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25093" *)
  wire _07415_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25103" *)
  wire _07416_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25113" *)
  wire _07417_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25123" *)
  wire _07418_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25133" *)
  wire _07419_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25143" *)
  wire _07420_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25153" *)
  wire _07421_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25163" *)
  wire _07422_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25173" *)
  wire _07423_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25183" *)
  wire _07424_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25193" *)
  wire _07425_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25203" *)
  wire _07426_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25213" *)
  wire _07427_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25223" *)
  wire _07428_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25233" *)
  wire _07429_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25243" *)
  wire _07430_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25253" *)
  wire _07431_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25263" *)
  wire _07432_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25317" *)
  wire _07433_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25327" *)
  wire _07434_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25337" *)
  wire _07435_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25347" *)
  wire _07436_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25357" *)
  wire _07437_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25367" *)
  wire _07438_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25377" *)
  wire _07439_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25387" *)
  wire _07440_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25397" *)
  wire _07441_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25407" *)
  wire _07442_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25417" *)
  wire _07443_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25427" *)
  wire _07444_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25437" *)
  wire _07445_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25447" *)
  wire _07446_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25457" *)
  wire _07447_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25467" *)
  wire _07448_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25477" *)
  wire _07449_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25487" *)
  wire _07450_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25497" *)
  wire _07451_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25507" *)
  wire _07452_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25517" *)
  wire _07453_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25527" *)
  wire _07454_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25537" *)
  wire _07455_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25547" *)
  wire _07456_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25557" *)
  wire _07457_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25567" *)
  wire _07458_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25577" *)
  wire _07459_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25587" *)
  wire _07460_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25597" *)
  wire _07461_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25607" *)
  wire _07462_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25617" *)
  wire _07463_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25627" *)
  wire _07464_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25637" *)
  wire _07465_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25647" *)
  wire _07466_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25657" *)
  wire _07467_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25667" *)
  wire _07468_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25677" *)
  wire _07469_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25687" *)
  wire _07470_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25697" *)
  wire _07471_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25707" *)
  wire _07472_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25717" *)
  wire _07473_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25727" *)
  wire _07474_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25737" *)
  wire _07475_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25747" *)
  wire _07476_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25757" *)
  wire _07477_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25767" *)
  wire _07478_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25777" *)
  wire _07479_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25787" *)
  wire _07480_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25797" *)
  wire _07481_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25807" *)
  wire _07482_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25817" *)
  wire _07483_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25827" *)
  wire _07484_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25837" *)
  wire _07485_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25847" *)
  wire _07486_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25857" *)
  wire _07487_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25867" *)
  wire _07488_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25877" *)
  wire _07489_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25887" *)
  wire _07490_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25897" *)
  wire _07491_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25907" *)
  wire _07492_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25917" *)
  wire _07493_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25927" *)
  wire _07494_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25937" *)
  wire _07495_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25947" *)
  wire _07496_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25957" *)
  wire _07497_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25967" *)
  wire _07498_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25977" *)
  wire _07499_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25987" *)
  wire _07500_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25997" *)
  wire _07501_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26007" *)
  wire _07502_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26017" *)
  wire _07503_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26027" *)
  wire _07504_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26037" *)
  wire _07505_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26047" *)
  wire _07506_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26057" *)
  wire _07507_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26067" *)
  wire _07508_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26077" *)
  wire _07509_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26087" *)
  wire _07510_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26097" *)
  wire _07511_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26107" *)
  wire _07512_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26117" *)
  wire _07513_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26127" *)
  wire _07514_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26137" *)
  wire _07515_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26147" *)
  wire _07516_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26157" *)
  wire _07517_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26167" *)
  wire _07518_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26177" *)
  wire _07519_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26187" *)
  wire _07520_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26197" *)
  wire _07521_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26207" *)
  wire _07522_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26217" *)
  wire _07523_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26227" *)
  wire _07524_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26237" *)
  wire _07525_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26247" *)
  wire _07526_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26257" *)
  wire _07527_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26267" *)
  wire _07528_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26277" *)
  wire _07529_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26287" *)
  wire _07530_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26297" *)
  wire _07531_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26307" *)
  wire _07532_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26317" *)
  wire _07533_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26327" *)
  wire _07534_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26337" *)
  wire _07535_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26347" *)
  wire _07536_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26357" *)
  wire _07537_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26367" *)
  wire _07538_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26377" *)
  wire _07539_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26387" *)
  wire _07540_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26397" *)
  wire _07541_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26407" *)
  wire _07542_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26417" *)
  wire _07543_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26427" *)
  wire _07544_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26437" *)
  wire _07545_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26447" *)
  wire _07546_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26457" *)
  wire _07547_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26467" *)
  wire _07548_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26477" *)
  wire _07549_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26487" *)
  wire _07550_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26497" *)
  wire _07551_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26507" *)
  wire _07552_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26517" *)
  wire _07553_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26527" *)
  wire _07554_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26537" *)
  wire _07555_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26547" *)
  wire _07556_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26557" *)
  wire _07557_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26567" *)
  wire _07558_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26577" *)
  wire _07559_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26587" *)
  wire _07560_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29032" *)
  wire [1023:0] _07561_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29086" *)
  wire _07562_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29096" *)
  wire _07563_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29106" *)
  wire _07564_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29116" *)
  wire _07565_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29126" *)
  wire _07566_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29136" *)
  wire _07567_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29146" *)
  wire _07568_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29156" *)
  wire _07569_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29166" *)
  wire _07570_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29176" *)
  wire _07571_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29186" *)
  wire _07572_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29196" *)
  wire _07573_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29206" *)
  wire _07574_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29216" *)
  wire _07575_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29226" *)
  wire _07576_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29236" *)
  wire _07577_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29246" *)
  wire _07578_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29256" *)
  wire _07579_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29266" *)
  wire _07580_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29276" *)
  wire _07581_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29286" *)
  wire _07582_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29296" *)
  wire _07583_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29306" *)
  wire _07584_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29316" *)
  wire _07585_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29326" *)
  wire _07586_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29336" *)
  wire _07587_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29346" *)
  wire _07588_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29356" *)
  wire _07589_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29366" *)
  wire _07590_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29376" *)
  wire _07591_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29386" *)
  wire _07592_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29396" *)
  wire _07593_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29406" *)
  wire _07594_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29416" *)
  wire _07595_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29426" *)
  wire _07596_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29436" *)
  wire _07597_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29446" *)
  wire _07598_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29456" *)
  wire _07599_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29466" *)
  wire _07600_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29476" *)
  wire _07601_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29486" *)
  wire _07602_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29496" *)
  wire _07603_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29506" *)
  wire _07604_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29516" *)
  wire _07605_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29526" *)
  wire _07606_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29536" *)
  wire _07607_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29546" *)
  wire _07608_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29556" *)
  wire _07609_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29566" *)
  wire _07610_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29576" *)
  wire _07611_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29586" *)
  wire _07612_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29596" *)
  wire _07613_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29606" *)
  wire _07614_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29616" *)
  wire _07615_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29626" *)
  wire _07616_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29636" *)
  wire _07617_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29646" *)
  wire _07618_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29656" *)
  wire _07619_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29666" *)
  wire _07620_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29676" *)
  wire _07621_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29686" *)
  wire _07622_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29696" *)
  wire _07623_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29706" *)
  wire _07624_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29716" *)
  wire _07625_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29726" *)
  wire _07626_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29736" *)
  wire _07627_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29746" *)
  wire _07628_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29756" *)
  wire _07629_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29766" *)
  wire _07630_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29776" *)
  wire _07631_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29786" *)
  wire _07632_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29796" *)
  wire _07633_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29806" *)
  wire _07634_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29816" *)
  wire _07635_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29826" *)
  wire _07636_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29836" *)
  wire _07637_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29846" *)
  wire _07638_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29856" *)
  wire _07639_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29866" *)
  wire _07640_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29876" *)
  wire _07641_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29886" *)
  wire _07642_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29896" *)
  wire _07643_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29906" *)
  wire _07644_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29916" *)
  wire _07645_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29926" *)
  wire _07646_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29936" *)
  wire _07647_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29946" *)
  wire _07648_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29956" *)
  wire _07649_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29966" *)
  wire _07650_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29976" *)
  wire _07651_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29986" *)
  wire _07652_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29996" *)
  wire _07653_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30006" *)
  wire _07654_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30016" *)
  wire _07655_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30026" *)
  wire _07656_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30036" *)
  wire _07657_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30046" *)
  wire _07658_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30056" *)
  wire _07659_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30066" *)
  wire _07660_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30076" *)
  wire _07661_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30086" *)
  wire _07662_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30096" *)
  wire _07663_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30106" *)
  wire _07664_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30116" *)
  wire _07665_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30126" *)
  wire _07666_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30136" *)
  wire _07667_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30146" *)
  wire _07668_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30156" *)
  wire _07669_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30166" *)
  wire _07670_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30176" *)
  wire _07671_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30186" *)
  wire _07672_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30196" *)
  wire _07673_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30206" *)
  wire _07674_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30216" *)
  wire _07675_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30226" *)
  wire _07676_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30236" *)
  wire _07677_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30246" *)
  wire _07678_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30256" *)
  wire _07679_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30266" *)
  wire _07680_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30276" *)
  wire _07681_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30286" *)
  wire _07682_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30296" *)
  wire _07683_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30306" *)
  wire _07684_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30316" *)
  wire _07685_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30326" *)
  wire _07686_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30336" *)
  wire _07687_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30346" *)
  wire _07688_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30356" *)
  wire _07689_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30674" *)
  wire _07690_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30684" *)
  wire _07691_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30694" *)
  wire _07692_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30704" *)
  wire _07693_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30714" *)
  wire _07694_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30724" *)
  wire _07695_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30734" *)
  wire _07696_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30744" *)
  wire _07697_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30754" *)
  wire _07698_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30764" *)
  wire _07699_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30774" *)
  wire _07700_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30784" *)
  wire _07701_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30794" *)
  wire _07702_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30804" *)
  wire _07703_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30814" *)
  wire _07704_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30824" *)
  wire _07705_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30834" *)
  wire _07706_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30844" *)
  wire _07707_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30854" *)
  wire _07708_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30864" *)
  wire _07709_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30874" *)
  wire _07710_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30884" *)
  wire _07711_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30894" *)
  wire _07712_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30904" *)
  wire _07713_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30914" *)
  wire _07714_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30924" *)
  wire _07715_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30934" *)
  wire _07716_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30944" *)
  wire _07717_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30954" *)
  wire _07718_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30964" *)
  wire _07719_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30974" *)
  wire _07720_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30984" *)
  wire _07721_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30994" *)
  wire _07722_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31004" *)
  wire _07723_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31014" *)
  wire _07724_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31024" *)
  wire _07725_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31034" *)
  wire _07726_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31044" *)
  wire _07727_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31054" *)
  wire _07728_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31064" *)
  wire _07729_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31074" *)
  wire _07730_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31084" *)
  wire _07731_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31094" *)
  wire _07732_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31104" *)
  wire _07733_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31114" *)
  wire _07734_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31124" *)
  wire _07735_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31134" *)
  wire _07736_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31144" *)
  wire _07737_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31154" *)
  wire _07738_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31164" *)
  wire _07739_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31174" *)
  wire _07740_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31184" *)
  wire _07741_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31194" *)
  wire _07742_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31204" *)
  wire _07743_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31214" *)
  wire _07744_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31224" *)
  wire _07745_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31234" *)
  wire _07746_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31244" *)
  wire _07747_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31254" *)
  wire _07748_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31264" *)
  wire _07749_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31274" *)
  wire _07750_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31284" *)
  wire _07751_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31294" *)
  wire _07752_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31304" *)
  wire _07753_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31314" *)
  wire _07754_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31324" *)
  wire _07755_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31334" *)
  wire _07756_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31344" *)
  wire _07757_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31354" *)
  wire _07758_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31364" *)
  wire _07759_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31374" *)
  wire _07760_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31384" *)
  wire _07761_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31394" *)
  wire _07762_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31404" *)
  wire _07763_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31414" *)
  wire _07764_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31424" *)
  wire _07765_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31434" *)
  wire _07766_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31444" *)
  wire _07767_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31454" *)
  wire _07768_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31464" *)
  wire _07769_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31474" *)
  wire _07770_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31484" *)
  wire _07771_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31494" *)
  wire _07772_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31504" *)
  wire _07773_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31514" *)
  wire _07774_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31524" *)
  wire _07775_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31534" *)
  wire _07776_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31544" *)
  wire _07777_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31554" *)
  wire _07778_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31564" *)
  wire _07779_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31574" *)
  wire _07780_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31584" *)
  wire _07781_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31594" *)
  wire _07782_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31604" *)
  wire _07783_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31614" *)
  wire _07784_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31624" *)
  wire _07785_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31634" *)
  wire _07786_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31644" *)
  wire _07787_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31654" *)
  wire _07788_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31664" *)
  wire _07789_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31674" *)
  wire _07790_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31684" *)
  wire _07791_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31694" *)
  wire _07792_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31704" *)
  wire _07793_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31714" *)
  wire _07794_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31724" *)
  wire _07795_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31734" *)
  wire _07796_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31744" *)
  wire _07797_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31754" *)
  wire _07798_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31764" *)
  wire _07799_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31774" *)
  wire _07800_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31784" *)
  wire _07801_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31794" *)
  wire _07802_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31804" *)
  wire _07803_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31814" *)
  wire _07804_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31824" *)
  wire _07805_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31834" *)
  wire _07806_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31844" *)
  wire _07807_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31854" *)
  wire _07808_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31864" *)
  wire _07809_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31874" *)
  wire _07810_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31884" *)
  wire _07811_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31894" *)
  wire _07812_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31904" *)
  wire _07813_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31914" *)
  wire _07814_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31924" *)
  wire _07815_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31934" *)
  wire _07816_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31944" *)
  wire _07817_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3959" *)
  wire [1023:0] _07818_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4033" *)
  wire _07819_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4043" *)
  wire _07820_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4053" *)
  wire _07821_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4063" *)
  wire _07822_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4073" *)
  wire _07823_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4083" *)
  wire _07824_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4093" *)
  wire _07825_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4103" *)
  wire _07826_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4113" *)
  wire _07827_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4123" *)
  wire _07828_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4133" *)
  wire _07829_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4143" *)
  wire _07830_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4153" *)
  wire _07831_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4163" *)
  wire _07832_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4173" *)
  wire _07833_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4183" *)
  wire _07834_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4193" *)
  wire _07835_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4203" *)
  wire _07836_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4213" *)
  wire _07837_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4223" *)
  wire _07838_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4233" *)
  wire _07839_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4243" *)
  wire _07840_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4253" *)
  wire _07841_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4263" *)
  wire _07842_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4273" *)
  wire _07843_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4283" *)
  wire _07844_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4293" *)
  wire _07845_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4303" *)
  wire _07846_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4313" *)
  wire _07847_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4323" *)
  wire _07848_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4333" *)
  wire _07849_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4343" *)
  wire _07850_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4353" *)
  wire _07851_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4363" *)
  wire _07852_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4373" *)
  wire _07853_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4383" *)
  wire _07854_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4393" *)
  wire _07855_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4403" *)
  wire _07856_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4413" *)
  wire _07857_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4423" *)
  wire _07858_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4433" *)
  wire _07859_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4443" *)
  wire _07860_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4453" *)
  wire _07861_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4463" *)
  wire _07862_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4473" *)
  wire _07863_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4483" *)
  wire _07864_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4493" *)
  wire _07865_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4503" *)
  wire _07866_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4513" *)
  wire _07867_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4523" *)
  wire _07868_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4533" *)
  wire _07869_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4543" *)
  wire _07870_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4553" *)
  wire _07871_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4563" *)
  wire _07872_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4573" *)
  wire _07873_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4583" *)
  wire _07874_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4593" *)
  wire _07875_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4603" *)
  wire _07876_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4613" *)
  wire _07877_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4623" *)
  wire _07878_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4633" *)
  wire _07879_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4643" *)
  wire _07880_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4653" *)
  wire _07881_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4663" *)
  wire _07882_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4673" *)
  wire _07883_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4683" *)
  wire _07884_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4693" *)
  wire _07885_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4703" *)
  wire _07886_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4713" *)
  wire _07887_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4723" *)
  wire _07888_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4733" *)
  wire _07889_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4743" *)
  wire _07890_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4753" *)
  wire _07891_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4763" *)
  wire _07892_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4773" *)
  wire _07893_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4783" *)
  wire _07894_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4793" *)
  wire _07895_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4803" *)
  wire _07896_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4813" *)
  wire _07897_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4823" *)
  wire _07898_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4833" *)
  wire _07899_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4843" *)
  wire _07900_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4853" *)
  wire _07901_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4863" *)
  wire _07902_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4873" *)
  wire _07903_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4883" *)
  wire _07904_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4893" *)
  wire _07905_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4903" *)
  wire _07906_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4913" *)
  wire _07907_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4923" *)
  wire _07908_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4933" *)
  wire _07909_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4943" *)
  wire _07910_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4953" *)
  wire _07911_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4963" *)
  wire _07912_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4973" *)
  wire _07913_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4983" *)
  wire _07914_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4993" *)
  wire _07915_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5003" *)
  wire _07916_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5013" *)
  wire _07917_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5023" *)
  wire _07918_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5033" *)
  wire _07919_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5043" *)
  wire _07920_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5053" *)
  wire _07921_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5063" *)
  wire _07922_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5073" *)
  wire _07923_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5083" *)
  wire _07924_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5093" *)
  wire _07925_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5103" *)
  wire _07926_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5113" *)
  wire _07927_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5123" *)
  wire _07928_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5133" *)
  wire _07929_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5143" *)
  wire _07930_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5153" *)
  wire _07931_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5163" *)
  wire _07932_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5173" *)
  wire _07933_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5183" *)
  wire _07934_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5193" *)
  wire _07935_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5203" *)
  wire _07936_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5213" *)
  wire _07937_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5223" *)
  wire _07938_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5233" *)
  wire _07939_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5243" *)
  wire _07940_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5253" *)
  wire _07941_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5263" *)
  wire _07942_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5273" *)
  wire _07943_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5283" *)
  wire _07944_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5293" *)
  wire _07945_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5303" *)
  wire _07946_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *)
  wire _07947_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *)
  wire _07948_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *)
  wire _07949_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *)
  wire _07950_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *)
  wire _07951_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *)
  wire _07952_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *)
  wire _07953_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *)
  wire _07954_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *)
  wire _07955_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *)
  wire _07956_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *)
  wire _07957_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *)
  wire _07958_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *)
  wire _07959_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *)
  wire _07960_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *)
  wire _07961_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *)
  wire _07962_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *)
  wire _07963_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *)
  wire _07964_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *)
  wire _07965_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *)
  wire _07966_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *)
  wire _07967_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *)
  wire _07968_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *)
  wire _07969_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *)
  wire _07970_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *)
  wire _07971_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *)
  wire _07972_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *)
  wire _07973_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *)
  wire _07974_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *)
  wire _07975_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *)
  wire _07976_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *)
  wire _07977_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *)
  wire _07978_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *)
  wire _07979_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *)
  wire _07980_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *)
  wire _07981_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *)
  wire _07982_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *)
  wire _07983_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *)
  wire _07984_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *)
  wire _07985_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *)
  wire _07986_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *)
  wire _07987_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *)
  wire _07988_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *)
  wire _07989_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *)
  wire _07990_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *)
  wire _07991_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *)
  wire _07992_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *)
  wire _07993_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *)
  wire _07994_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *)
  wire _07995_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *)
  wire _07996_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *)
  wire _07997_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *)
  wire _07998_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *)
  wire _07999_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *)
  wire _08000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *)
  wire _08001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *)
  wire _08002_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *)
  wire _08003_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *)
  wire _08004_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *)
  wire _08005_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *)
  wire _08006_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *)
  wire _08007_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *)
  wire _08008_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *)
  wire _08009_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *)
  wire _08010_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *)
  wire _08011_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *)
  wire _08012_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *)
  wire _08013_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *)
  wire _08014_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *)
  wire _08015_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *)
  wire _08016_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *)
  wire _08017_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *)
  wire _08018_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *)
  wire _08019_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *)
  wire _08020_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *)
  wire _08021_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *)
  wire _08022_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *)
  wire _08023_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *)
  wire _08024_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *)
  wire _08025_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *)
  wire _08026_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *)
  wire _08027_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *)
  wire _08028_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *)
  wire _08029_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *)
  wire _08030_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *)
  wire _08031_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *)
  wire _08032_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *)
  wire _08033_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *)
  wire _08034_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *)
  wire _08035_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *)
  wire _08036_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *)
  wire _08037_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *)
  wire _08038_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *)
  wire _08039_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *)
  wire _08040_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *)
  wire _08041_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *)
  wire _08042_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *)
  wire _08043_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *)
  wire _08044_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *)
  wire _08045_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *)
  wire _08046_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *)
  wire _08047_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *)
  wire _08048_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *)
  wire _08049_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *)
  wire _08050_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *)
  wire _08051_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *)
  wire _08052_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *)
  wire _08053_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *)
  wire _08054_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *)
  wire _08055_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *)
  wire _08056_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *)
  wire _08057_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *)
  wire _08058_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *)
  wire _08059_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *)
  wire _08060_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *)
  wire _08061_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *)
  wire _08062_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *)
  wire _08063_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *)
  wire _08064_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *)
  wire _08065_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *)
  wire _08066_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *)
  wire _08067_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *)
  wire _08068_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *)
  wire _08069_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *)
  wire _08070_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *)
  wire _08071_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *)
  wire _08072_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *)
  wire _08073_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *)
  wire _08074_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *)
  wire _08075_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *)
  wire _08076_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *)
  wire _08077_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *)
  wire _08078_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *)
  wire _08079_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *)
  wire _08080_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *)
  wire _08081_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *)
  wire _08082_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *)
  wire _08083_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *)
  wire _08084_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *)
  wire _08085_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *)
  wire _08086_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *)
  wire _08087_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *)
  wire _08088_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *)
  wire _08089_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *)
  wire _08090_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *)
  wire _08091_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *)
  wire _08092_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *)
  wire _08093_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *)
  wire _08094_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *)
  wire _08095_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *)
  wire _08096_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *)
  wire _08097_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *)
  wire _08098_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *)
  wire _08099_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *)
  wire _08100_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *)
  wire _08101_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *)
  wire _08102_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *)
  wire _08103_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *)
  wire _08104_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *)
  wire _08105_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *)
  wire _08106_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *)
  wire _08107_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *)
  wire _08108_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *)
  wire _08109_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *)
  wire _08110_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *)
  wire _08111_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *)
  wire _08112_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *)
  wire _08113_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *)
  wire _08114_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *)
  wire _08115_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *)
  wire _08116_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *)
  wire _08117_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *)
  wire _08118_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *)
  wire _08119_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *)
  wire _08120_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *)
  wire _08121_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *)
  wire _08122_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *)
  wire _08123_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *)
  wire _08124_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *)
  wire _08125_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *)
  wire _08126_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *)
  wire _08127_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *)
  wire _08128_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *)
  wire _08129_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *)
  wire _08130_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *)
  wire _08131_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *)
  wire _08132_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *)
  wire _08133_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *)
  wire _08134_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *)
  wire _08135_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *)
  wire _08136_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *)
  wire _08137_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *)
  wire _08138_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2727" *)
  wire _08139_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2728" *)
  wire _08140_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2729" *)
  wire _08141_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2730" *)
  wire _08142_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2731" *)
  wire _08143_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2732" *)
  wire _08144_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2733" *)
  wire _08145_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2734" *)
  wire _08146_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2735" *)
  wire _08147_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2736" *)
  wire _08148_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2737" *)
  wire _08149_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2738" *)
  wire _08150_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2739" *)
  wire _08151_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2740" *)
  wire _08152_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2741" *)
  wire _08153_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2742" *)
  wire _08154_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2743" *)
  wire _08155_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2744" *)
  wire _08156_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2745" *)
  wire _08157_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2746" *)
  wire _08158_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2747" *)
  wire _08159_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2748" *)
  wire _08160_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2749" *)
  wire _08161_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2750" *)
  wire _08162_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2751" *)
  wire _08163_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2752" *)
  wire _08164_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2753" *)
  wire _08165_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2754" *)
  wire _08166_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2755" *)
  wire _08167_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2756" *)
  wire _08168_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2757" *)
  wire _08169_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2758" *)
  wire _08170_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2759" *)
  wire _08171_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2760" *)
  wire _08172_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2761" *)
  wire _08173_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2762" *)
  wire _08174_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2763" *)
  wire _08175_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2764" *)
  wire _08176_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2765" *)
  wire _08177_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2766" *)
  wire _08178_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *)
  wire _08179_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *)
  wire _08180_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *)
  wire _08181_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *)
  wire _08182_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *)
  wire _08183_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *)
  wire _08184_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *)
  wire _08185_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *)
  wire _08186_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *)
  wire _08187_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2767" *)
  wire _08188_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *)
  wire _08189_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *)
  wire _08190_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *)
  wire _08191_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *)
  wire _08192_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *)
  wire _08193_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *)
  wire _08194_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *)
  wire _08195_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *)
  wire _08196_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *)
  wire _08197_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *)
  wire _08198_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2768" *)
  wire _08199_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *)
  wire _08200_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *)
  wire _08201_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *)
  wire _08202_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *)
  wire _08203_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *)
  wire _08204_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *)
  wire _08205_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *)
  wire _08206_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *)
  wire _08207_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *)
  wire _08208_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *)
  wire _08209_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2769" *)
  wire _08210_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *)
  wire _08211_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *)
  wire _08212_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *)
  wire _08213_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *)
  wire _08214_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *)
  wire _08215_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *)
  wire _08216_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *)
  wire _08217_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *)
  wire _08218_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *)
  wire _08219_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *)
  wire _08220_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2770" *)
  wire _08221_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *)
  wire _08222_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *)
  wire _08223_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *)
  wire _08224_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *)
  wire _08225_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *)
  wire _08226_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *)
  wire _08227_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *)
  wire _08228_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *)
  wire _08229_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *)
  wire _08230_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *)
  wire _08231_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2771" *)
  wire _08232_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *)
  wire _08233_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *)
  wire _08234_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *)
  wire _08235_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *)
  wire _08236_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *)
  wire _08237_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *)
  wire _08238_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *)
  wire _08239_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *)
  wire _08240_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *)
  wire _08241_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *)
  wire _08242_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2772" *)
  wire _08243_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *)
  wire _08244_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *)
  wire _08245_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *)
  wire _08246_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *)
  wire _08247_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *)
  wire _08248_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2773" *)
  wire _08249_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2774" *)
  wire _08250_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2775" *)
  wire _08251_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2776" *)
  wire _08252_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2777" *)
  wire _08253_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2778" *)
  wire _08254_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2779" *)
  wire _08255_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2780" *)
  wire _08256_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27800" *)
  wire _08257_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27801" *)
  wire _08258_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27802" *)
  wire _08259_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27803" *)
  wire _08260_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27804" *)
  wire _08261_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27805" *)
  wire _08262_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27806" *)
  wire _08263_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27807" *)
  wire _08264_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27808" *)
  wire _08265_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27809" *)
  wire _08266_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2781" *)
  wire _08267_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27810" *)
  wire _08268_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27811" *)
  wire _08269_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27812" *)
  wire _08270_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27813" *)
  wire _08271_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27814" *)
  wire _08272_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27815" *)
  wire _08273_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27816" *)
  wire _08274_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27817" *)
  wire _08275_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27818" *)
  wire _08276_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27819" *)
  wire _08277_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2782" *)
  wire _08278_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27820" *)
  wire _08279_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27821" *)
  wire _08280_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27822" *)
  wire _08281_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27823" *)
  wire _08282_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27824" *)
  wire _08283_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27825" *)
  wire _08284_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27826" *)
  wire _08285_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27827" *)
  wire _08286_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27828" *)
  wire _08287_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27829" *)
  wire _08288_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2783" *)
  wire _08289_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27830" *)
  wire _08290_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27831" *)
  wire _08291_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27832" *)
  wire _08292_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27833" *)
  wire _08293_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27834" *)
  wire _08294_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27835" *)
  wire _08295_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27836" *)
  wire _08296_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27837" *)
  wire _08297_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27838" *)
  wire _08298_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27839" *)
  wire _08299_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2784" *)
  wire _08300_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27840" *)
  wire _08301_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27841" *)
  wire _08302_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27842" *)
  wire _08303_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27843" *)
  wire _08304_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27844" *)
  wire _08305_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27845" *)
  wire _08306_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27846" *)
  wire _08307_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27847" *)
  wire _08308_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27848" *)
  wire _08309_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27849" *)
  wire _08310_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2785" *)
  wire _08311_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27850" *)
  wire _08312_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27851" *)
  wire _08313_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27852" *)
  wire _08314_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27853" *)
  wire _08315_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27854" *)
  wire _08316_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27855" *)
  wire _08317_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27856" *)
  wire _08318_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27857" *)
  wire _08319_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27858" *)
  wire _08320_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27859" *)
  wire _08321_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2786" *)
  wire _08322_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27860" *)
  wire _08323_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27861" *)
  wire _08324_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27862" *)
  wire _08325_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27863" *)
  wire _08326_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2787" *)
  wire _08327_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2788" *)
  wire _08328_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2789" *)
  wire _08329_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2790" *)
  wire _08330_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10666" *)
  wire _08331_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12002" *)
  wire _08332_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13338" *)
  wire _08333_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14674" *)
  wire _08334_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16011" *)
  wire _08335_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17335" *)
  wire _08336_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18659" *)
  wire _08337_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19983" *)
  wire _08338_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21307" *)
  wire _08339_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22631" *)
  wire _08340_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23955" *)
  wire _08341_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25279" *)
  wire _08342_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29043" *)
  wire [127:0] _08343_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3970" *)
  wire [127:0] _08344_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5322" *)
  wire _08345_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6658" *)
  wire _08346_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7994" *)
  wire _08347_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9330" *)
  wire _08348_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:410" *)
  input cfg_is_fp16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:805" *)
  reg [97:0] cfg_is_fp16_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:411" *)
  input cfg_is_int16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:806" *)
  reg [63:0] cfg_is_int16_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:412" *)
  input cfg_is_int8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:807" *)
  reg [64:0] cfg_is_int8_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:413" *)
  input cfg_reg_en;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:677" *)
  output [1023:0] dat0_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:678" *)
  output [63:0] dat0_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:679" *)
  output [127:0] dat0_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:680" *)
  output [103:0] dat0_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:681" *)
  output [191:0] dat0_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:682" *)
  output [63:0] dat0_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:683" *)
  output dat0_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:684" *)
  output dat0_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:685" *)
  output dat0_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:686" *)
  output [1023:0] dat1_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:687" *)
  output [63:0] dat1_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:688" *)
  output [127:0] dat1_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:689" *)
  output [103:0] dat1_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:690" *)
  output [191:0] dat1_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:691" *)
  output [63:0] dat1_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:692" *)
  output dat1_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:693" *)
  output dat1_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:694" *)
  output dat1_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:695" *)
  output [1023:0] dat2_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:696" *)
  output [63:0] dat2_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:697" *)
  output [127:0] dat2_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:698" *)
  output [103:0] dat2_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:699" *)
  output [191:0] dat2_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:700" *)
  output [63:0] dat2_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:701" *)
  output dat2_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:702" *)
  output dat2_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:703" *)
  output dat2_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:704" *)
  output [1023:0] dat3_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:705" *)
  output [63:0] dat3_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:706" *)
  output [127:0] dat3_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:707" *)
  output [103:0] dat3_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:708" *)
  output [191:0] dat3_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:709" *)
  output [63:0] dat3_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:710" *)
  output dat3_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:711" *)
  output dat3_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:712" *)
  output dat3_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:713" *)
  output [1023:0] dat4_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:714" *)
  output [63:0] dat4_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:715" *)
  output [127:0] dat4_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:716" *)
  output [103:0] dat4_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:717" *)
  output [191:0] dat4_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:718" *)
  output [63:0] dat4_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:719" *)
  output dat4_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:720" *)
  output dat4_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:721" *)
  output dat4_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:722" *)
  output [1023:0] dat5_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:723" *)
  output [63:0] dat5_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:724" *)
  output [127:0] dat5_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:725" *)
  output [103:0] dat5_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:726" *)
  output [191:0] dat5_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:727" *)
  output [63:0] dat5_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:728" *)
  output dat5_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:729" *)
  output dat5_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:730" *)
  output dat5_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:731" *)
  output [1023:0] dat6_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:732" *)
  output [63:0] dat6_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:733" *)
  output [127:0] dat6_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:734" *)
  output [103:0] dat6_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:735" *)
  output [191:0] dat6_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:736" *)
  output [63:0] dat6_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:737" *)
  output dat6_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:738" *)
  output dat6_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:739" *)
  output dat6_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:740" *)
  output [1023:0] dat7_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:741" *)
  output [63:0] dat7_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:742" *)
  output [127:0] dat7_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:743" *)
  output [103:0] dat7_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:744" *)
  output [191:0] dat7_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:745" *)
  output [63:0] dat7_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:746" *)
  output dat7_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:747" *)
  output dat7_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:748" *)
  output dat7_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:880" *)
  reg [1023:0] dat_actv_data_reg0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:881" *)
  reg [1023:0] dat_actv_data_reg1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:882" *)
  reg [1023:0] dat_actv_data_reg2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:883" *)
  reg [1023:0] dat_actv_data_reg3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:884" *)
  reg [1023:0] dat_actv_data_reg4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:885" *)
  reg [1023:0] dat_actv_data_reg5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:886" *)
  reg [1023:0] dat_actv_data_reg6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:887" *)
  reg [1023:0] dat_actv_data_reg7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:888" *)
  reg [63:0] dat_actv_nan_reg0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:889" *)
  reg [63:0] dat_actv_nan_reg1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:890" *)
  reg [63:0] dat_actv_nan_reg2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:891" *)
  reg [63:0] dat_actv_nan_reg3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:892" *)
  reg [63:0] dat_actv_nan_reg4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:893" *)
  reg [63:0] dat_actv_nan_reg5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:894" *)
  reg [63:0] dat_actv_nan_reg6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:895" *)
  reg [63:0] dat_actv_nan_reg7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:896" *)
  reg [127:0] dat_actv_nz_reg0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:897" *)
  reg [127:0] dat_actv_nz_reg1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:898" *)
  reg [127:0] dat_actv_nz_reg2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:899" *)
  reg [127:0] dat_actv_nz_reg3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:900" *)
  reg [127:0] dat_actv_nz_reg4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:901" *)
  reg [127:0] dat_actv_nz_reg5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:902" *)
  reg [127:0] dat_actv_nz_reg6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:903" *)
  reg [127:0] dat_actv_nz_reg7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:904" *)
  wire [103:0] dat_actv_pvld_reg0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:905" *)
  wire [103:0] dat_actv_pvld_reg1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:906" *)
  wire [103:0] dat_actv_pvld_reg2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:907" *)
  wire [103:0] dat_actv_pvld_reg3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:908" *)
  wire [103:0] dat_actv_pvld_reg4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:909" *)
  wire [103:0] dat_actv_pvld_reg5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:910" *)
  wire [103:0] dat_actv_pvld_reg6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:911" *)
  wire [103:0] dat_actv_pvld_reg7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:912" *)
  reg dat_actv_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:913" *)
  wire dat_has_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:914" *)
  reg [1023:0] dat_pre_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:915" *)
  wire [1023:0] dat_pre_data_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:916" *)
  reg [191:0] dat_pre_exp_reg0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:917" *)
  reg [191:0] dat_pre_exp_reg1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:918" *)
  reg [191:0] dat_pre_exp_reg2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:919" *)
  reg [191:0] dat_pre_exp_reg3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:920" *)
  reg [191:0] dat_pre_exp_reg4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:921" *)
  reg [191:0] dat_pre_exp_reg5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:922" *)
  reg [191:0] dat_pre_exp_reg6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:923" *)
  reg [191:0] dat_pre_exp_reg7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:924" *)
  wire [191:0] dat_pre_exp_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:925" *)
  reg [63:0] dat_pre_mask0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:926" *)
  reg [63:0] dat_pre_mask1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:927" *)
  reg [63:0] dat_pre_mask2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:928" *)
  reg [63:0] dat_pre_mask3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:929" *)
  reg [63:0] dat_pre_mask4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:930" *)
  reg [63:0] dat_pre_mask5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:931" *)
  reg [63:0] dat_pre_mask6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:932" *)
  reg [63:0] dat_pre_mask7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:933" *)
  wire [63:0] dat_pre_mask_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:934" *)
  reg [63:0] dat_pre_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:935" *)
  reg [127:0] dat_pre_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:936" *)
  wire [127:0] dat_pre_nz_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:937" *)
  wire [15:0] dat_pre_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:938" *)
  wire [8:0] dat_pre_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:939" *)
  wire [15:0] dat_pre_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:414" *)
  input [7:0] in_dat_data0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:415" *)
  input [7:0] in_dat_data1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:416" *)
  input [7:0] in_dat_data10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:417" *)
  input [7:0] in_dat_data100;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:418" *)
  input [7:0] in_dat_data101;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:419" *)
  input [7:0] in_dat_data102;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:420" *)
  input [7:0] in_dat_data103;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:421" *)
  input [7:0] in_dat_data104;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:422" *)
  input [7:0] in_dat_data105;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:423" *)
  input [7:0] in_dat_data106;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:424" *)
  input [7:0] in_dat_data107;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:425" *)
  input [7:0] in_dat_data108;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:426" *)
  input [7:0] in_dat_data109;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:427" *)
  input [7:0] in_dat_data11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:428" *)
  input [7:0] in_dat_data110;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:429" *)
  input [7:0] in_dat_data111;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:430" *)
  input [7:0] in_dat_data112;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:431" *)
  input [7:0] in_dat_data113;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:432" *)
  input [7:0] in_dat_data114;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:433" *)
  input [7:0] in_dat_data115;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:434" *)
  input [7:0] in_dat_data116;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:435" *)
  input [7:0] in_dat_data117;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:436" *)
  input [7:0] in_dat_data118;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:437" *)
  input [7:0] in_dat_data119;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:438" *)
  input [7:0] in_dat_data12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:439" *)
  input [7:0] in_dat_data120;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:440" *)
  input [7:0] in_dat_data121;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:441" *)
  input [7:0] in_dat_data122;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:442" *)
  input [7:0] in_dat_data123;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:443" *)
  input [7:0] in_dat_data124;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:444" *)
  input [7:0] in_dat_data125;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:445" *)
  input [7:0] in_dat_data126;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:446" *)
  input [7:0] in_dat_data127;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:447" *)
  input [7:0] in_dat_data13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:448" *)
  input [7:0] in_dat_data14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:449" *)
  input [7:0] in_dat_data15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:450" *)
  input [7:0] in_dat_data16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:451" *)
  input [7:0] in_dat_data17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:452" *)
  input [7:0] in_dat_data18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:453" *)
  input [7:0] in_dat_data19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:454" *)
  input [7:0] in_dat_data2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:455" *)
  input [7:0] in_dat_data20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:456" *)
  input [7:0] in_dat_data21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:457" *)
  input [7:0] in_dat_data22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:458" *)
  input [7:0] in_dat_data23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:459" *)
  input [7:0] in_dat_data24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:460" *)
  input [7:0] in_dat_data25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:461" *)
  input [7:0] in_dat_data26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:462" *)
  input [7:0] in_dat_data27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:463" *)
  input [7:0] in_dat_data28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:464" *)
  input [7:0] in_dat_data29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:465" *)
  input [7:0] in_dat_data3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:466" *)
  input [7:0] in_dat_data30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:467" *)
  input [7:0] in_dat_data31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:468" *)
  input [7:0] in_dat_data32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:469" *)
  input [7:0] in_dat_data33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:470" *)
  input [7:0] in_dat_data34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:471" *)
  input [7:0] in_dat_data35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:472" *)
  input [7:0] in_dat_data36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:473" *)
  input [7:0] in_dat_data37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:474" *)
  input [7:0] in_dat_data38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:475" *)
  input [7:0] in_dat_data39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:476" *)
  input [7:0] in_dat_data4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:477" *)
  input [7:0] in_dat_data40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:478" *)
  input [7:0] in_dat_data41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:479" *)
  input [7:0] in_dat_data42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:480" *)
  input [7:0] in_dat_data43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:481" *)
  input [7:0] in_dat_data44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:482" *)
  input [7:0] in_dat_data45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:483" *)
  input [7:0] in_dat_data46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:484" *)
  input [7:0] in_dat_data47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:485" *)
  input [7:0] in_dat_data48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:486" *)
  input [7:0] in_dat_data49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:487" *)
  input [7:0] in_dat_data5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:488" *)
  input [7:0] in_dat_data50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:489" *)
  input [7:0] in_dat_data51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:490" *)
  input [7:0] in_dat_data52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:491" *)
  input [7:0] in_dat_data53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:492" *)
  input [7:0] in_dat_data54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:493" *)
  input [7:0] in_dat_data55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:494" *)
  input [7:0] in_dat_data56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:495" *)
  input [7:0] in_dat_data57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:496" *)
  input [7:0] in_dat_data58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:497" *)
  input [7:0] in_dat_data59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:498" *)
  input [7:0] in_dat_data6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:499" *)
  input [7:0] in_dat_data60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:500" *)
  input [7:0] in_dat_data61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:501" *)
  input [7:0] in_dat_data62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:502" *)
  input [7:0] in_dat_data63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:503" *)
  input [7:0] in_dat_data64;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:504" *)
  input [7:0] in_dat_data65;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:505" *)
  input [7:0] in_dat_data66;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:506" *)
  input [7:0] in_dat_data67;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:507" *)
  input [7:0] in_dat_data68;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:508" *)
  input [7:0] in_dat_data69;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:509" *)
  input [7:0] in_dat_data7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:510" *)
  input [7:0] in_dat_data70;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:511" *)
  input [7:0] in_dat_data71;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:512" *)
  input [7:0] in_dat_data72;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:513" *)
  input [7:0] in_dat_data73;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:514" *)
  input [7:0] in_dat_data74;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:515" *)
  input [7:0] in_dat_data75;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:516" *)
  input [7:0] in_dat_data76;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:517" *)
  input [7:0] in_dat_data77;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:518" *)
  input [7:0] in_dat_data78;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:519" *)
  input [7:0] in_dat_data79;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:520" *)
  input [7:0] in_dat_data8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:521" *)
  input [7:0] in_dat_data80;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:522" *)
  input [7:0] in_dat_data81;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:523" *)
  input [7:0] in_dat_data82;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:524" *)
  input [7:0] in_dat_data83;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:525" *)
  input [7:0] in_dat_data84;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:526" *)
  input [7:0] in_dat_data85;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:527" *)
  input [7:0] in_dat_data86;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:528" *)
  input [7:0] in_dat_data87;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:529" *)
  input [7:0] in_dat_data88;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:530" *)
  input [7:0] in_dat_data89;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:531" *)
  input [7:0] in_dat_data9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:532" *)
  input [7:0] in_dat_data90;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:533" *)
  input [7:0] in_dat_data91;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:534" *)
  input [7:0] in_dat_data92;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:535" *)
  input [7:0] in_dat_data93;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:536" *)
  input [7:0] in_dat_data94;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:537" *)
  input [7:0] in_dat_data95;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:538" *)
  input [7:0] in_dat_data96;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:539" *)
  input [7:0] in_dat_data97;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:540" *)
  input [7:0] in_dat_data98;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:541" *)
  input [7:0] in_dat_data99;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:940" *)
  wire [1023:0] in_dat_data_fp16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:941" *)
  wire [15:0] in_dat_data_fp16_0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:942" *)
  wire [15:0] in_dat_data_fp16_1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:943" *)
  wire [15:0] in_dat_data_fp16_10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:944" *)
  wire [15:0] in_dat_data_fp16_11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:945" *)
  wire [15:0] in_dat_data_fp16_12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:946" *)
  wire [15:0] in_dat_data_fp16_13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:947" *)
  wire [15:0] in_dat_data_fp16_14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:948" *)
  wire [15:0] in_dat_data_fp16_15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:949" *)
  wire [15:0] in_dat_data_fp16_16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:950" *)
  wire [15:0] in_dat_data_fp16_17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:951" *)
  wire [15:0] in_dat_data_fp16_18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:952" *)
  wire [15:0] in_dat_data_fp16_19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:953" *)
  wire [15:0] in_dat_data_fp16_2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:954" *)
  wire [15:0] in_dat_data_fp16_20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:955" *)
  wire [15:0] in_dat_data_fp16_21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:956" *)
  wire [15:0] in_dat_data_fp16_22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:957" *)
  wire [15:0] in_dat_data_fp16_23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:958" *)
  wire [15:0] in_dat_data_fp16_24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:959" *)
  wire [15:0] in_dat_data_fp16_25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:960" *)
  wire [15:0] in_dat_data_fp16_26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:961" *)
  wire [15:0] in_dat_data_fp16_27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:962" *)
  wire [15:0] in_dat_data_fp16_28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:963" *)
  wire [15:0] in_dat_data_fp16_29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:964" *)
  wire [15:0] in_dat_data_fp16_3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:965" *)
  wire [15:0] in_dat_data_fp16_30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:966" *)
  wire [15:0] in_dat_data_fp16_31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:967" *)
  wire [15:0] in_dat_data_fp16_32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:968" *)
  wire [15:0] in_dat_data_fp16_33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:969" *)
  wire [15:0] in_dat_data_fp16_34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:970" *)
  wire [15:0] in_dat_data_fp16_35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:971" *)
  wire [15:0] in_dat_data_fp16_36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:972" *)
  wire [15:0] in_dat_data_fp16_37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:973" *)
  wire [15:0] in_dat_data_fp16_38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:974" *)
  wire [15:0] in_dat_data_fp16_39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:975" *)
  wire [15:0] in_dat_data_fp16_4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:976" *)
  wire [15:0] in_dat_data_fp16_40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:977" *)
  wire [15:0] in_dat_data_fp16_41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:978" *)
  wire [15:0] in_dat_data_fp16_42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:979" *)
  wire [15:0] in_dat_data_fp16_43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:980" *)
  wire [15:0] in_dat_data_fp16_44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:981" *)
  wire [15:0] in_dat_data_fp16_45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:982" *)
  wire [15:0] in_dat_data_fp16_46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:983" *)
  wire [15:0] in_dat_data_fp16_47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:984" *)
  wire [15:0] in_dat_data_fp16_48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:985" *)
  wire [15:0] in_dat_data_fp16_49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:986" *)
  wire [15:0] in_dat_data_fp16_5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:987" *)
  wire [15:0] in_dat_data_fp16_50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:988" *)
  wire [15:0] in_dat_data_fp16_51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:989" *)
  wire [15:0] in_dat_data_fp16_52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:990" *)
  wire [15:0] in_dat_data_fp16_53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:991" *)
  wire [15:0] in_dat_data_fp16_54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:992" *)
  wire [15:0] in_dat_data_fp16_55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:993" *)
  wire [15:0] in_dat_data_fp16_56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:994" *)
  wire [15:0] in_dat_data_fp16_57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:995" *)
  wire [15:0] in_dat_data_fp16_58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:996" *)
  wire [15:0] in_dat_data_fp16_59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:997" *)
  wire [15:0] in_dat_data_fp16_6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:998" *)
  wire [15:0] in_dat_data_fp16_60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:999" *)
  wire [15:0] in_dat_data_fp16_61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1000" *)
  wire [15:0] in_dat_data_fp16_62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1001" *)
  wire [15:0] in_dat_data_fp16_63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1002" *)
  wire [15:0] in_dat_data_fp16_7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1003" *)
  wire [15:0] in_dat_data_fp16_8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1004" *)
  wire [15:0] in_dat_data_fp16_9;
  wire [10:0] in_dat_data_fp16_mts_ori0;
  wire [10:0] in_dat_data_fp16_mts_ori1;
  wire [10:0] in_dat_data_fp16_mts_ori10;
  wire [10:0] in_dat_data_fp16_mts_ori11;
  wire [10:0] in_dat_data_fp16_mts_ori12;
  wire [10:0] in_dat_data_fp16_mts_ori13;
  wire [10:0] in_dat_data_fp16_mts_ori14;
  wire [10:0] in_dat_data_fp16_mts_ori15;
  wire [10:0] in_dat_data_fp16_mts_ori16;
  wire [10:0] in_dat_data_fp16_mts_ori17;
  wire [10:0] in_dat_data_fp16_mts_ori18;
  wire [10:0] in_dat_data_fp16_mts_ori19;
  wire [10:0] in_dat_data_fp16_mts_ori2;
  wire [10:0] in_dat_data_fp16_mts_ori20;
  wire [10:0] in_dat_data_fp16_mts_ori21;
  wire [10:0] in_dat_data_fp16_mts_ori22;
  wire [10:0] in_dat_data_fp16_mts_ori23;
  wire [10:0] in_dat_data_fp16_mts_ori24;
  wire [10:0] in_dat_data_fp16_mts_ori25;
  wire [10:0] in_dat_data_fp16_mts_ori26;
  wire [10:0] in_dat_data_fp16_mts_ori27;
  wire [10:0] in_dat_data_fp16_mts_ori28;
  wire [10:0] in_dat_data_fp16_mts_ori29;
  wire [10:0] in_dat_data_fp16_mts_ori3;
  wire [10:0] in_dat_data_fp16_mts_ori30;
  wire [10:0] in_dat_data_fp16_mts_ori31;
  wire [10:0] in_dat_data_fp16_mts_ori32;
  wire [10:0] in_dat_data_fp16_mts_ori33;
  wire [10:0] in_dat_data_fp16_mts_ori34;
  wire [10:0] in_dat_data_fp16_mts_ori35;
  wire [10:0] in_dat_data_fp16_mts_ori36;
  wire [10:0] in_dat_data_fp16_mts_ori37;
  wire [10:0] in_dat_data_fp16_mts_ori38;
  wire [10:0] in_dat_data_fp16_mts_ori39;
  wire [10:0] in_dat_data_fp16_mts_ori4;
  wire [10:0] in_dat_data_fp16_mts_ori40;
  wire [10:0] in_dat_data_fp16_mts_ori41;
  wire [10:0] in_dat_data_fp16_mts_ori42;
  wire [10:0] in_dat_data_fp16_mts_ori43;
  wire [10:0] in_dat_data_fp16_mts_ori44;
  wire [10:0] in_dat_data_fp16_mts_ori45;
  wire [10:0] in_dat_data_fp16_mts_ori46;
  wire [10:0] in_dat_data_fp16_mts_ori47;
  wire [10:0] in_dat_data_fp16_mts_ori48;
  wire [10:0] in_dat_data_fp16_mts_ori49;
  wire [10:0] in_dat_data_fp16_mts_ori5;
  wire [10:0] in_dat_data_fp16_mts_ori50;
  wire [10:0] in_dat_data_fp16_mts_ori51;
  wire [10:0] in_dat_data_fp16_mts_ori52;
  wire [10:0] in_dat_data_fp16_mts_ori53;
  wire [10:0] in_dat_data_fp16_mts_ori54;
  wire [10:0] in_dat_data_fp16_mts_ori55;
  wire [10:0] in_dat_data_fp16_mts_ori56;
  wire [10:0] in_dat_data_fp16_mts_ori57;
  wire [10:0] in_dat_data_fp16_mts_ori58;
  wire [10:0] in_dat_data_fp16_mts_ori59;
  wire [10:0] in_dat_data_fp16_mts_ori6;
  wire [10:0] in_dat_data_fp16_mts_ori60;
  wire [10:0] in_dat_data_fp16_mts_ori61;
  wire [10:0] in_dat_data_fp16_mts_ori62;
  wire [10:0] in_dat_data_fp16_mts_ori63;
  wire [10:0] in_dat_data_fp16_mts_ori7;
  wire [10:0] in_dat_data_fp16_mts_ori8;
  wire [10:0] in_dat_data_fp16_mts_ori9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1069" *)
  wire [14:0] in_dat_data_fp16_mts_sft0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1070" *)
  wire [14:0] in_dat_data_fp16_mts_sft1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1071" *)
  wire [14:0] in_dat_data_fp16_mts_sft10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1072" *)
  wire [14:0] in_dat_data_fp16_mts_sft11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1073" *)
  wire [14:0] in_dat_data_fp16_mts_sft12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1074" *)
  wire [14:0] in_dat_data_fp16_mts_sft13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1075" *)
  wire [14:0] in_dat_data_fp16_mts_sft14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1076" *)
  wire [14:0] in_dat_data_fp16_mts_sft15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1077" *)
  wire [14:0] in_dat_data_fp16_mts_sft16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1078" *)
  wire [14:0] in_dat_data_fp16_mts_sft17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1079" *)
  wire [14:0] in_dat_data_fp16_mts_sft18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1080" *)
  wire [14:0] in_dat_data_fp16_mts_sft19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1081" *)
  wire [14:0] in_dat_data_fp16_mts_sft2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1082" *)
  wire [14:0] in_dat_data_fp16_mts_sft20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1083" *)
  wire [14:0] in_dat_data_fp16_mts_sft21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1084" *)
  wire [14:0] in_dat_data_fp16_mts_sft22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1085" *)
  wire [14:0] in_dat_data_fp16_mts_sft23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1086" *)
  wire [14:0] in_dat_data_fp16_mts_sft24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1087" *)
  wire [14:0] in_dat_data_fp16_mts_sft25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1088" *)
  wire [14:0] in_dat_data_fp16_mts_sft26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1089" *)
  wire [14:0] in_dat_data_fp16_mts_sft27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1090" *)
  wire [14:0] in_dat_data_fp16_mts_sft28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1091" *)
  wire [14:0] in_dat_data_fp16_mts_sft29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1092" *)
  wire [14:0] in_dat_data_fp16_mts_sft3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1093" *)
  wire [14:0] in_dat_data_fp16_mts_sft30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1094" *)
  wire [14:0] in_dat_data_fp16_mts_sft31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1095" *)
  wire [14:0] in_dat_data_fp16_mts_sft32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1096" *)
  wire [14:0] in_dat_data_fp16_mts_sft33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1097" *)
  wire [14:0] in_dat_data_fp16_mts_sft34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1098" *)
  wire [14:0] in_dat_data_fp16_mts_sft35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1099" *)
  wire [14:0] in_dat_data_fp16_mts_sft36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1100" *)
  wire [14:0] in_dat_data_fp16_mts_sft37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1101" *)
  wire [14:0] in_dat_data_fp16_mts_sft38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1102" *)
  wire [14:0] in_dat_data_fp16_mts_sft39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1103" *)
  wire [14:0] in_dat_data_fp16_mts_sft4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1104" *)
  wire [14:0] in_dat_data_fp16_mts_sft40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1105" *)
  wire [14:0] in_dat_data_fp16_mts_sft41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1106" *)
  wire [14:0] in_dat_data_fp16_mts_sft42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1107" *)
  wire [14:0] in_dat_data_fp16_mts_sft43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1108" *)
  wire [14:0] in_dat_data_fp16_mts_sft44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1109" *)
  wire [14:0] in_dat_data_fp16_mts_sft45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1110" *)
  wire [14:0] in_dat_data_fp16_mts_sft46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1111" *)
  wire [14:0] in_dat_data_fp16_mts_sft47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1112" *)
  wire [14:0] in_dat_data_fp16_mts_sft48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1113" *)
  wire [14:0] in_dat_data_fp16_mts_sft49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1114" *)
  wire [14:0] in_dat_data_fp16_mts_sft5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1115" *)
  wire [14:0] in_dat_data_fp16_mts_sft50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1116" *)
  wire [14:0] in_dat_data_fp16_mts_sft51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1117" *)
  wire [14:0] in_dat_data_fp16_mts_sft52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1118" *)
  wire [14:0] in_dat_data_fp16_mts_sft53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1119" *)
  wire [14:0] in_dat_data_fp16_mts_sft54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1120" *)
  wire [14:0] in_dat_data_fp16_mts_sft55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1121" *)
  wire [14:0] in_dat_data_fp16_mts_sft56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1122" *)
  wire [14:0] in_dat_data_fp16_mts_sft57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1123" *)
  wire [14:0] in_dat_data_fp16_mts_sft58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1124" *)
  wire [14:0] in_dat_data_fp16_mts_sft59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1125" *)
  wire [14:0] in_dat_data_fp16_mts_sft6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1126" *)
  wire [14:0] in_dat_data_fp16_mts_sft60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1127" *)
  wire [14:0] in_dat_data_fp16_mts_sft61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1128" *)
  wire [14:0] in_dat_data_fp16_mts_sft62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1129" *)
  wire [14:0] in_dat_data_fp16_mts_sft63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1130" *)
  wire [14:0] in_dat_data_fp16_mts_sft7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1131" *)
  wire [14:0] in_dat_data_fp16_mts_sft8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1132" *)
  wire [14:0] in_dat_data_fp16_mts_sft9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1133" *)
  wire [1023:0] in_dat_data_int16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1134" *)
  wire [15:0] in_dat_data_int16_0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1135" *)
  wire [15:0] in_dat_data_int16_1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1136" *)
  wire [15:0] in_dat_data_int16_10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1137" *)
  wire [15:0] in_dat_data_int16_11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1138" *)
  wire [15:0] in_dat_data_int16_12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1139" *)
  wire [15:0] in_dat_data_int16_13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1140" *)
  wire [15:0] in_dat_data_int16_14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1141" *)
  wire [15:0] in_dat_data_int16_15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1142" *)
  wire [15:0] in_dat_data_int16_16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1143" *)
  wire [15:0] in_dat_data_int16_17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1144" *)
  wire [15:0] in_dat_data_int16_18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1145" *)
  wire [15:0] in_dat_data_int16_19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1146" *)
  wire [15:0] in_dat_data_int16_2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1147" *)
  wire [15:0] in_dat_data_int16_20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1148" *)
  wire [15:0] in_dat_data_int16_21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1149" *)
  wire [15:0] in_dat_data_int16_22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1150" *)
  wire [15:0] in_dat_data_int16_23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1151" *)
  wire [15:0] in_dat_data_int16_24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1152" *)
  wire [15:0] in_dat_data_int16_25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1153" *)
  wire [15:0] in_dat_data_int16_26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1154" *)
  wire [15:0] in_dat_data_int16_27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1155" *)
  wire [15:0] in_dat_data_int16_28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1156" *)
  wire [15:0] in_dat_data_int16_29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1157" *)
  wire [15:0] in_dat_data_int16_3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1158" *)
  wire [15:0] in_dat_data_int16_30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1159" *)
  wire [15:0] in_dat_data_int16_31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1160" *)
  wire [15:0] in_dat_data_int16_32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1161" *)
  wire [15:0] in_dat_data_int16_33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1162" *)
  wire [15:0] in_dat_data_int16_34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1163" *)
  wire [15:0] in_dat_data_int16_35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1164" *)
  wire [15:0] in_dat_data_int16_36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1165" *)
  wire [15:0] in_dat_data_int16_37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1166" *)
  wire [15:0] in_dat_data_int16_38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1167" *)
  wire [15:0] in_dat_data_int16_39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1168" *)
  wire [15:0] in_dat_data_int16_4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1169" *)
  wire [15:0] in_dat_data_int16_40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1170" *)
  wire [15:0] in_dat_data_int16_41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1171" *)
  wire [15:0] in_dat_data_int16_42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1172" *)
  wire [15:0] in_dat_data_int16_43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1173" *)
  wire [15:0] in_dat_data_int16_44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1174" *)
  wire [15:0] in_dat_data_int16_45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1175" *)
  wire [15:0] in_dat_data_int16_46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1176" *)
  wire [15:0] in_dat_data_int16_47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1177" *)
  wire [15:0] in_dat_data_int16_48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1178" *)
  wire [15:0] in_dat_data_int16_49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1179" *)
  wire [15:0] in_dat_data_int16_5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1180" *)
  wire [15:0] in_dat_data_int16_50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1181" *)
  wire [15:0] in_dat_data_int16_51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1182" *)
  wire [15:0] in_dat_data_int16_52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1183" *)
  wire [15:0] in_dat_data_int16_53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1184" *)
  wire [15:0] in_dat_data_int16_54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1185" *)
  wire [15:0] in_dat_data_int16_55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1186" *)
  wire [15:0] in_dat_data_int16_56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1187" *)
  wire [15:0] in_dat_data_int16_57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1188" *)
  wire [15:0] in_dat_data_int16_58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1189" *)
  wire [15:0] in_dat_data_int16_59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1190" *)
  wire [15:0] in_dat_data_int16_6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1191" *)
  wire [15:0] in_dat_data_int16_60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1192" *)
  wire [15:0] in_dat_data_int16_61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1193" *)
  wire [15:0] in_dat_data_int16_62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1194" *)
  wire [15:0] in_dat_data_int16_63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1195" *)
  wire [15:0] in_dat_data_int16_7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1196" *)
  wire [15:0] in_dat_data_int16_8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1197" *)
  wire [15:0] in_dat_data_int16_9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1198" *)
  wire [1023:0] in_dat_data_int8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1199" *)
  wire [15:0] in_dat_data_int8_0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1200" *)
  wire [15:0] in_dat_data_int8_1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1201" *)
  wire [15:0] in_dat_data_int8_10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1202" *)
  wire [15:0] in_dat_data_int8_11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1203" *)
  wire [15:0] in_dat_data_int8_12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1204" *)
  wire [15:0] in_dat_data_int8_13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1205" *)
  wire [15:0] in_dat_data_int8_14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1206" *)
  wire [15:0] in_dat_data_int8_15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1207" *)
  wire [15:0] in_dat_data_int8_16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1208" *)
  wire [15:0] in_dat_data_int8_17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1209" *)
  wire [15:0] in_dat_data_int8_18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1210" *)
  wire [15:0] in_dat_data_int8_19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1211" *)
  wire [15:0] in_dat_data_int8_2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1212" *)
  wire [15:0] in_dat_data_int8_20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1213" *)
  wire [15:0] in_dat_data_int8_21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1214" *)
  wire [15:0] in_dat_data_int8_22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1215" *)
  wire [15:0] in_dat_data_int8_23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1216" *)
  wire [15:0] in_dat_data_int8_24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1217" *)
  wire [15:0] in_dat_data_int8_25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1218" *)
  wire [15:0] in_dat_data_int8_26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1219" *)
  wire [15:0] in_dat_data_int8_27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1220" *)
  wire [15:0] in_dat_data_int8_28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1221" *)
  wire [15:0] in_dat_data_int8_29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1222" *)
  wire [15:0] in_dat_data_int8_3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1223" *)
  wire [15:0] in_dat_data_int8_30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1224" *)
  wire [15:0] in_dat_data_int8_31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1225" *)
  wire [15:0] in_dat_data_int8_32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1226" *)
  wire [15:0] in_dat_data_int8_33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1227" *)
  wire [15:0] in_dat_data_int8_34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1228" *)
  wire [15:0] in_dat_data_int8_35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1229" *)
  wire [15:0] in_dat_data_int8_36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1230" *)
  wire [15:0] in_dat_data_int8_37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1231" *)
  wire [15:0] in_dat_data_int8_38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1232" *)
  wire [15:0] in_dat_data_int8_39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1233" *)
  wire [15:0] in_dat_data_int8_4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1234" *)
  wire [15:0] in_dat_data_int8_40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1235" *)
  wire [15:0] in_dat_data_int8_41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1236" *)
  wire [15:0] in_dat_data_int8_42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1237" *)
  wire [15:0] in_dat_data_int8_43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1238" *)
  wire [15:0] in_dat_data_int8_44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1239" *)
  wire [15:0] in_dat_data_int8_45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1240" *)
  wire [15:0] in_dat_data_int8_46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1241" *)
  wire [15:0] in_dat_data_int8_47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1242" *)
  wire [15:0] in_dat_data_int8_48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1243" *)
  wire [15:0] in_dat_data_int8_49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1244" *)
  wire [15:0] in_dat_data_int8_5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1245" *)
  wire [15:0] in_dat_data_int8_50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1246" *)
  wire [15:0] in_dat_data_int8_51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1247" *)
  wire [15:0] in_dat_data_int8_52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1248" *)
  wire [15:0] in_dat_data_int8_53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1249" *)
  wire [15:0] in_dat_data_int8_54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1250" *)
  wire [15:0] in_dat_data_int8_55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1251" *)
  wire [15:0] in_dat_data_int8_56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1252" *)
  wire [15:0] in_dat_data_int8_57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1253" *)
  wire [15:0] in_dat_data_int8_58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1254" *)
  wire [15:0] in_dat_data_int8_59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1255" *)
  wire [15:0] in_dat_data_int8_6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1256" *)
  wire [15:0] in_dat_data_int8_60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1257" *)
  wire [15:0] in_dat_data_int8_61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1258" *)
  wire [15:0] in_dat_data_int8_62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1259" *)
  wire [15:0] in_dat_data_int8_63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1260" *)
  wire [15:0] in_dat_data_int8_7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1261" *)
  wire [15:0] in_dat_data_int8_8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1262" *)
  wire [15:0] in_dat_data_int8_9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1263" *)
  wire [1023:0] in_dat_data_pack;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1264" *)
  wire [191:0] in_dat_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:542" *)
  input [127:0] in_dat_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1265" *)
  wire [127:0] in_dat_mask_int8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1266" *)
  wire [63:0] in_dat_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1267" *)
  wire [63:0] in_dat_norm;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:543" *)
  input in_dat_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:544" *)
  input in_dat_stripe_end;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:545" *)
  input in_dat_stripe_st;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:546" *)
  input [7:0] in_wt_data0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:547" *)
  input [7:0] in_wt_data1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:548" *)
  input [7:0] in_wt_data10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:549" *)
  input [7:0] in_wt_data100;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:550" *)
  input [7:0] in_wt_data101;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:551" *)
  input [7:0] in_wt_data102;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:552" *)
  input [7:0] in_wt_data103;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:553" *)
  input [7:0] in_wt_data104;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:554" *)
  input [7:0] in_wt_data105;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:555" *)
  input [7:0] in_wt_data106;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:556" *)
  input [7:0] in_wt_data107;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:557" *)
  input [7:0] in_wt_data108;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:558" *)
  input [7:0] in_wt_data109;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:559" *)
  input [7:0] in_wt_data11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:560" *)
  input [7:0] in_wt_data110;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:561" *)
  input [7:0] in_wt_data111;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:562" *)
  input [7:0] in_wt_data112;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:563" *)
  input [7:0] in_wt_data113;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:564" *)
  input [7:0] in_wt_data114;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:565" *)
  input [7:0] in_wt_data115;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:566" *)
  input [7:0] in_wt_data116;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:567" *)
  input [7:0] in_wt_data117;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:568" *)
  input [7:0] in_wt_data118;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:569" *)
  input [7:0] in_wt_data119;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:570" *)
  input [7:0] in_wt_data12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:571" *)
  input [7:0] in_wt_data120;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:572" *)
  input [7:0] in_wt_data121;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:573" *)
  input [7:0] in_wt_data122;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:574" *)
  input [7:0] in_wt_data123;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:575" *)
  input [7:0] in_wt_data124;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:576" *)
  input [7:0] in_wt_data125;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:577" *)
  input [7:0] in_wt_data126;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:578" *)
  input [7:0] in_wt_data127;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:579" *)
  input [7:0] in_wt_data13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:580" *)
  input [7:0] in_wt_data14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:581" *)
  input [7:0] in_wt_data15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:582" *)
  input [7:0] in_wt_data16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:583" *)
  input [7:0] in_wt_data17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:584" *)
  input [7:0] in_wt_data18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:585" *)
  input [7:0] in_wt_data19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:586" *)
  input [7:0] in_wt_data2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:587" *)
  input [7:0] in_wt_data20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:588" *)
  input [7:0] in_wt_data21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:589" *)
  input [7:0] in_wt_data22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:590" *)
  input [7:0] in_wt_data23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:591" *)
  input [7:0] in_wt_data24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:592" *)
  input [7:0] in_wt_data25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:593" *)
  input [7:0] in_wt_data26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:594" *)
  input [7:0] in_wt_data27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:595" *)
  input [7:0] in_wt_data28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:596" *)
  input [7:0] in_wt_data29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:597" *)
  input [7:0] in_wt_data3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:598" *)
  input [7:0] in_wt_data30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:599" *)
  input [7:0] in_wt_data31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:600" *)
  input [7:0] in_wt_data32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:601" *)
  input [7:0] in_wt_data33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:602" *)
  input [7:0] in_wt_data34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:603" *)
  input [7:0] in_wt_data35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:604" *)
  input [7:0] in_wt_data36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:605" *)
  input [7:0] in_wt_data37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:606" *)
  input [7:0] in_wt_data38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:607" *)
  input [7:0] in_wt_data39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:608" *)
  input [7:0] in_wt_data4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:609" *)
  input [7:0] in_wt_data40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:610" *)
  input [7:0] in_wt_data41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:611" *)
  input [7:0] in_wt_data42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:612" *)
  input [7:0] in_wt_data43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:613" *)
  input [7:0] in_wt_data44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:614" *)
  input [7:0] in_wt_data45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:615" *)
  input [7:0] in_wt_data46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:616" *)
  input [7:0] in_wt_data47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:617" *)
  input [7:0] in_wt_data48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:618" *)
  input [7:0] in_wt_data49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:619" *)
  input [7:0] in_wt_data5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:620" *)
  input [7:0] in_wt_data50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:621" *)
  input [7:0] in_wt_data51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:622" *)
  input [7:0] in_wt_data52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:623" *)
  input [7:0] in_wt_data53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:624" *)
  input [7:0] in_wt_data54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:625" *)
  input [7:0] in_wt_data55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:626" *)
  input [7:0] in_wt_data56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:627" *)
  input [7:0] in_wt_data57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:628" *)
  input [7:0] in_wt_data58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:629" *)
  input [7:0] in_wt_data59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:630" *)
  input [7:0] in_wt_data6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:631" *)
  input [7:0] in_wt_data60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:632" *)
  input [7:0] in_wt_data61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:633" *)
  input [7:0] in_wt_data62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:634" *)
  input [7:0] in_wt_data63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:635" *)
  input [7:0] in_wt_data64;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:636" *)
  input [7:0] in_wt_data65;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:637" *)
  input [7:0] in_wt_data66;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:638" *)
  input [7:0] in_wt_data67;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:639" *)
  input [7:0] in_wt_data68;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:640" *)
  input [7:0] in_wt_data69;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:641" *)
  input [7:0] in_wt_data7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:642" *)
  input [7:0] in_wt_data70;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:643" *)
  input [7:0] in_wt_data71;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:644" *)
  input [7:0] in_wt_data72;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:645" *)
  input [7:0] in_wt_data73;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:646" *)
  input [7:0] in_wt_data74;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:647" *)
  input [7:0] in_wt_data75;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:648" *)
  input [7:0] in_wt_data76;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:649" *)
  input [7:0] in_wt_data77;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:650" *)
  input [7:0] in_wt_data78;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:651" *)
  input [7:0] in_wt_data79;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:652" *)
  input [7:0] in_wt_data8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:653" *)
  input [7:0] in_wt_data80;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:654" *)
  input [7:0] in_wt_data81;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:655" *)
  input [7:0] in_wt_data82;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:656" *)
  input [7:0] in_wt_data83;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:657" *)
  input [7:0] in_wt_data84;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:658" *)
  input [7:0] in_wt_data85;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:659" *)
  input [7:0] in_wt_data86;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:660" *)
  input [7:0] in_wt_data87;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:661" *)
  input [7:0] in_wt_data88;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:662" *)
  input [7:0] in_wt_data89;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:663" *)
  input [7:0] in_wt_data9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:664" *)
  input [7:0] in_wt_data90;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:665" *)
  input [7:0] in_wt_data91;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:666" *)
  input [7:0] in_wt_data92;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:667" *)
  input [7:0] in_wt_data93;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:668" *)
  input [7:0] in_wt_data94;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:669" *)
  input [7:0] in_wt_data95;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:670" *)
  input [7:0] in_wt_data96;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:671" *)
  input [7:0] in_wt_data97;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:672" *)
  input [7:0] in_wt_data98;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:673" *)
  input [7:0] in_wt_data99;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1268" *)
  wire [1023:0] in_wt_data_fp16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1269" *)
  wire [15:0] in_wt_data_fp16_0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1270" *)
  wire [15:0] in_wt_data_fp16_1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1271" *)
  wire [15:0] in_wt_data_fp16_10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1272" *)
  wire [15:0] in_wt_data_fp16_11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1273" *)
  wire [15:0] in_wt_data_fp16_12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1274" *)
  wire [15:0] in_wt_data_fp16_13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1275" *)
  wire [15:0] in_wt_data_fp16_14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1276" *)
  wire [15:0] in_wt_data_fp16_15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1277" *)
  wire [15:0] in_wt_data_fp16_16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1278" *)
  wire [15:0] in_wt_data_fp16_17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1279" *)
  wire [15:0] in_wt_data_fp16_18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1280" *)
  wire [15:0] in_wt_data_fp16_19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1281" *)
  wire [15:0] in_wt_data_fp16_2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1282" *)
  wire [15:0] in_wt_data_fp16_20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1283" *)
  wire [15:0] in_wt_data_fp16_21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1284" *)
  wire [15:0] in_wt_data_fp16_22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1285" *)
  wire [15:0] in_wt_data_fp16_23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1286" *)
  wire [15:0] in_wt_data_fp16_24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1287" *)
  wire [15:0] in_wt_data_fp16_25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1288" *)
  wire [15:0] in_wt_data_fp16_26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1289" *)
  wire [15:0] in_wt_data_fp16_27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1290" *)
  wire [15:0] in_wt_data_fp16_28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1291" *)
  wire [15:0] in_wt_data_fp16_29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1292" *)
  wire [15:0] in_wt_data_fp16_3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1293" *)
  wire [15:0] in_wt_data_fp16_30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1294" *)
  wire [15:0] in_wt_data_fp16_31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1295" *)
  wire [15:0] in_wt_data_fp16_32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1296" *)
  wire [15:0] in_wt_data_fp16_33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1297" *)
  wire [15:0] in_wt_data_fp16_34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1298" *)
  wire [15:0] in_wt_data_fp16_35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1299" *)
  wire [15:0] in_wt_data_fp16_36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1300" *)
  wire [15:0] in_wt_data_fp16_37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1301" *)
  wire [15:0] in_wt_data_fp16_38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1302" *)
  wire [15:0] in_wt_data_fp16_39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1303" *)
  wire [15:0] in_wt_data_fp16_4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1304" *)
  wire [15:0] in_wt_data_fp16_40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1305" *)
  wire [15:0] in_wt_data_fp16_41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1306" *)
  wire [15:0] in_wt_data_fp16_42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1307" *)
  wire [15:0] in_wt_data_fp16_43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1308" *)
  wire [15:0] in_wt_data_fp16_44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1309" *)
  wire [15:0] in_wt_data_fp16_45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1310" *)
  wire [15:0] in_wt_data_fp16_46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1311" *)
  wire [15:0] in_wt_data_fp16_47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1312" *)
  wire [15:0] in_wt_data_fp16_48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1313" *)
  wire [15:0] in_wt_data_fp16_49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1314" *)
  wire [15:0] in_wt_data_fp16_5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1315" *)
  wire [15:0] in_wt_data_fp16_50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1316" *)
  wire [15:0] in_wt_data_fp16_51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1317" *)
  wire [15:0] in_wt_data_fp16_52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1318" *)
  wire [15:0] in_wt_data_fp16_53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1319" *)
  wire [15:0] in_wt_data_fp16_54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1320" *)
  wire [15:0] in_wt_data_fp16_55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1321" *)
  wire [15:0] in_wt_data_fp16_56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1322" *)
  wire [15:0] in_wt_data_fp16_57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1323" *)
  wire [15:0] in_wt_data_fp16_58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1324" *)
  wire [15:0] in_wt_data_fp16_59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1325" *)
  wire [15:0] in_wt_data_fp16_6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1326" *)
  wire [15:0] in_wt_data_fp16_60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1327" *)
  wire [15:0] in_wt_data_fp16_61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1328" *)
  wire [15:0] in_wt_data_fp16_62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1329" *)
  wire [15:0] in_wt_data_fp16_63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1330" *)
  wire [15:0] in_wt_data_fp16_7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1331" *)
  wire [15:0] in_wt_data_fp16_8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1332" *)
  wire [15:0] in_wt_data_fp16_9;
  wire [10:0] in_wt_data_fp16_mts_ori0;
  wire [10:0] in_wt_data_fp16_mts_ori1;
  wire [10:0] in_wt_data_fp16_mts_ori10;
  wire [10:0] in_wt_data_fp16_mts_ori11;
  wire [10:0] in_wt_data_fp16_mts_ori12;
  wire [10:0] in_wt_data_fp16_mts_ori13;
  wire [10:0] in_wt_data_fp16_mts_ori14;
  wire [10:0] in_wt_data_fp16_mts_ori15;
  wire [10:0] in_wt_data_fp16_mts_ori16;
  wire [10:0] in_wt_data_fp16_mts_ori17;
  wire [10:0] in_wt_data_fp16_mts_ori18;
  wire [10:0] in_wt_data_fp16_mts_ori19;
  wire [10:0] in_wt_data_fp16_mts_ori2;
  wire [10:0] in_wt_data_fp16_mts_ori20;
  wire [10:0] in_wt_data_fp16_mts_ori21;
  wire [10:0] in_wt_data_fp16_mts_ori22;
  wire [10:0] in_wt_data_fp16_mts_ori23;
  wire [10:0] in_wt_data_fp16_mts_ori24;
  wire [10:0] in_wt_data_fp16_mts_ori25;
  wire [10:0] in_wt_data_fp16_mts_ori26;
  wire [10:0] in_wt_data_fp16_mts_ori27;
  wire [10:0] in_wt_data_fp16_mts_ori28;
  wire [10:0] in_wt_data_fp16_mts_ori29;
  wire [10:0] in_wt_data_fp16_mts_ori3;
  wire [10:0] in_wt_data_fp16_mts_ori30;
  wire [10:0] in_wt_data_fp16_mts_ori31;
  wire [10:0] in_wt_data_fp16_mts_ori32;
  wire [10:0] in_wt_data_fp16_mts_ori33;
  wire [10:0] in_wt_data_fp16_mts_ori34;
  wire [10:0] in_wt_data_fp16_mts_ori35;
  wire [10:0] in_wt_data_fp16_mts_ori36;
  wire [10:0] in_wt_data_fp16_mts_ori37;
  wire [10:0] in_wt_data_fp16_mts_ori38;
  wire [10:0] in_wt_data_fp16_mts_ori39;
  wire [10:0] in_wt_data_fp16_mts_ori4;
  wire [10:0] in_wt_data_fp16_mts_ori40;
  wire [10:0] in_wt_data_fp16_mts_ori41;
  wire [10:0] in_wt_data_fp16_mts_ori42;
  wire [10:0] in_wt_data_fp16_mts_ori43;
  wire [10:0] in_wt_data_fp16_mts_ori44;
  wire [10:0] in_wt_data_fp16_mts_ori45;
  wire [10:0] in_wt_data_fp16_mts_ori46;
  wire [10:0] in_wt_data_fp16_mts_ori47;
  wire [10:0] in_wt_data_fp16_mts_ori48;
  wire [10:0] in_wt_data_fp16_mts_ori49;
  wire [10:0] in_wt_data_fp16_mts_ori5;
  wire [10:0] in_wt_data_fp16_mts_ori50;
  wire [10:0] in_wt_data_fp16_mts_ori51;
  wire [10:0] in_wt_data_fp16_mts_ori52;
  wire [10:0] in_wt_data_fp16_mts_ori53;
  wire [10:0] in_wt_data_fp16_mts_ori54;
  wire [10:0] in_wt_data_fp16_mts_ori55;
  wire [10:0] in_wt_data_fp16_mts_ori56;
  wire [10:0] in_wt_data_fp16_mts_ori57;
  wire [10:0] in_wt_data_fp16_mts_ori58;
  wire [10:0] in_wt_data_fp16_mts_ori59;
  wire [10:0] in_wt_data_fp16_mts_ori6;
  wire [10:0] in_wt_data_fp16_mts_ori60;
  wire [10:0] in_wt_data_fp16_mts_ori61;
  wire [10:0] in_wt_data_fp16_mts_ori62;
  wire [10:0] in_wt_data_fp16_mts_ori63;
  wire [10:0] in_wt_data_fp16_mts_ori7;
  wire [10:0] in_wt_data_fp16_mts_ori8;
  wire [10:0] in_wt_data_fp16_mts_ori9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1397" *)
  wire [14:0] in_wt_data_fp16_mts_sft0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1398" *)
  wire [14:0] in_wt_data_fp16_mts_sft1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1399" *)
  wire [14:0] in_wt_data_fp16_mts_sft10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1400" *)
  wire [14:0] in_wt_data_fp16_mts_sft11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1401" *)
  wire [14:0] in_wt_data_fp16_mts_sft12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1402" *)
  wire [14:0] in_wt_data_fp16_mts_sft13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1403" *)
  wire [14:0] in_wt_data_fp16_mts_sft14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1404" *)
  wire [14:0] in_wt_data_fp16_mts_sft15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1405" *)
  wire [14:0] in_wt_data_fp16_mts_sft16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1406" *)
  wire [14:0] in_wt_data_fp16_mts_sft17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1407" *)
  wire [14:0] in_wt_data_fp16_mts_sft18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1408" *)
  wire [14:0] in_wt_data_fp16_mts_sft19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1409" *)
  wire [14:0] in_wt_data_fp16_mts_sft2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1410" *)
  wire [14:0] in_wt_data_fp16_mts_sft20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1411" *)
  wire [14:0] in_wt_data_fp16_mts_sft21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1412" *)
  wire [14:0] in_wt_data_fp16_mts_sft22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1413" *)
  wire [14:0] in_wt_data_fp16_mts_sft23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1414" *)
  wire [14:0] in_wt_data_fp16_mts_sft24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1415" *)
  wire [14:0] in_wt_data_fp16_mts_sft25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1416" *)
  wire [14:0] in_wt_data_fp16_mts_sft26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1417" *)
  wire [14:0] in_wt_data_fp16_mts_sft27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1418" *)
  wire [14:0] in_wt_data_fp16_mts_sft28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1419" *)
  wire [14:0] in_wt_data_fp16_mts_sft29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1420" *)
  wire [14:0] in_wt_data_fp16_mts_sft3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1421" *)
  wire [14:0] in_wt_data_fp16_mts_sft30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1422" *)
  wire [14:0] in_wt_data_fp16_mts_sft31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1423" *)
  wire [14:0] in_wt_data_fp16_mts_sft32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1424" *)
  wire [14:0] in_wt_data_fp16_mts_sft33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1425" *)
  wire [14:0] in_wt_data_fp16_mts_sft34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1426" *)
  wire [14:0] in_wt_data_fp16_mts_sft35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1427" *)
  wire [14:0] in_wt_data_fp16_mts_sft36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1428" *)
  wire [14:0] in_wt_data_fp16_mts_sft37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1429" *)
  wire [14:0] in_wt_data_fp16_mts_sft38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1430" *)
  wire [14:0] in_wt_data_fp16_mts_sft39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1431" *)
  wire [14:0] in_wt_data_fp16_mts_sft4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1432" *)
  wire [14:0] in_wt_data_fp16_mts_sft40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1433" *)
  wire [14:0] in_wt_data_fp16_mts_sft41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1434" *)
  wire [14:0] in_wt_data_fp16_mts_sft42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1435" *)
  wire [14:0] in_wt_data_fp16_mts_sft43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1436" *)
  wire [14:0] in_wt_data_fp16_mts_sft44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1437" *)
  wire [14:0] in_wt_data_fp16_mts_sft45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1438" *)
  wire [14:0] in_wt_data_fp16_mts_sft46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1439" *)
  wire [14:0] in_wt_data_fp16_mts_sft47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1440" *)
  wire [14:0] in_wt_data_fp16_mts_sft48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1441" *)
  wire [14:0] in_wt_data_fp16_mts_sft49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1442" *)
  wire [14:0] in_wt_data_fp16_mts_sft5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1443" *)
  wire [14:0] in_wt_data_fp16_mts_sft50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1444" *)
  wire [14:0] in_wt_data_fp16_mts_sft51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1445" *)
  wire [14:0] in_wt_data_fp16_mts_sft52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1446" *)
  wire [14:0] in_wt_data_fp16_mts_sft53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1447" *)
  wire [14:0] in_wt_data_fp16_mts_sft54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1448" *)
  wire [14:0] in_wt_data_fp16_mts_sft55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1449" *)
  wire [14:0] in_wt_data_fp16_mts_sft56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1450" *)
  wire [14:0] in_wt_data_fp16_mts_sft57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1451" *)
  wire [14:0] in_wt_data_fp16_mts_sft58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1452" *)
  wire [14:0] in_wt_data_fp16_mts_sft59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1453" *)
  wire [14:0] in_wt_data_fp16_mts_sft6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1454" *)
  wire [14:0] in_wt_data_fp16_mts_sft60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1455" *)
  wire [14:0] in_wt_data_fp16_mts_sft61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1456" *)
  wire [14:0] in_wt_data_fp16_mts_sft62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1457" *)
  wire [14:0] in_wt_data_fp16_mts_sft63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1458" *)
  wire [14:0] in_wt_data_fp16_mts_sft7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1459" *)
  wire [14:0] in_wt_data_fp16_mts_sft8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1460" *)
  wire [14:0] in_wt_data_fp16_mts_sft9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1461" *)
  wire [1023:0] in_wt_data_int16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1462" *)
  wire [15:0] in_wt_data_int16_0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1463" *)
  wire [15:0] in_wt_data_int16_1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1464" *)
  wire [15:0] in_wt_data_int16_10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1465" *)
  wire [15:0] in_wt_data_int16_11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1466" *)
  wire [15:0] in_wt_data_int16_12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1467" *)
  wire [15:0] in_wt_data_int16_13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1468" *)
  wire [15:0] in_wt_data_int16_14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1469" *)
  wire [15:0] in_wt_data_int16_15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1470" *)
  wire [15:0] in_wt_data_int16_16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1471" *)
  wire [15:0] in_wt_data_int16_17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1472" *)
  wire [15:0] in_wt_data_int16_18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1473" *)
  wire [15:0] in_wt_data_int16_19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1474" *)
  wire [15:0] in_wt_data_int16_2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1475" *)
  wire [15:0] in_wt_data_int16_20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1476" *)
  wire [15:0] in_wt_data_int16_21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1477" *)
  wire [15:0] in_wt_data_int16_22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1478" *)
  wire [15:0] in_wt_data_int16_23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1479" *)
  wire [15:0] in_wt_data_int16_24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1480" *)
  wire [15:0] in_wt_data_int16_25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1481" *)
  wire [15:0] in_wt_data_int16_26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1482" *)
  wire [15:0] in_wt_data_int16_27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1483" *)
  wire [15:0] in_wt_data_int16_28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1484" *)
  wire [15:0] in_wt_data_int16_29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1485" *)
  wire [15:0] in_wt_data_int16_3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1486" *)
  wire [15:0] in_wt_data_int16_30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1487" *)
  wire [15:0] in_wt_data_int16_31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1488" *)
  wire [15:0] in_wt_data_int16_32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1489" *)
  wire [15:0] in_wt_data_int16_33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1490" *)
  wire [15:0] in_wt_data_int16_34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1491" *)
  wire [15:0] in_wt_data_int16_35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1492" *)
  wire [15:0] in_wt_data_int16_36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1493" *)
  wire [15:0] in_wt_data_int16_37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1494" *)
  wire [15:0] in_wt_data_int16_38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1495" *)
  wire [15:0] in_wt_data_int16_39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1496" *)
  wire [15:0] in_wt_data_int16_4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1497" *)
  wire [15:0] in_wt_data_int16_40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1498" *)
  wire [15:0] in_wt_data_int16_41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1499" *)
  wire [15:0] in_wt_data_int16_42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1500" *)
  wire [15:0] in_wt_data_int16_43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1501" *)
  wire [15:0] in_wt_data_int16_44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1502" *)
  wire [15:0] in_wt_data_int16_45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1503" *)
  wire [15:0] in_wt_data_int16_46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1504" *)
  wire [15:0] in_wt_data_int16_47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1505" *)
  wire [15:0] in_wt_data_int16_48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1506" *)
  wire [15:0] in_wt_data_int16_49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1507" *)
  wire [15:0] in_wt_data_int16_5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1508" *)
  wire [15:0] in_wt_data_int16_50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1509" *)
  wire [15:0] in_wt_data_int16_51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1510" *)
  wire [15:0] in_wt_data_int16_52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1511" *)
  wire [15:0] in_wt_data_int16_53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1512" *)
  wire [15:0] in_wt_data_int16_54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1513" *)
  wire [15:0] in_wt_data_int16_55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1514" *)
  wire [15:0] in_wt_data_int16_56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1515" *)
  wire [15:0] in_wt_data_int16_57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1516" *)
  wire [15:0] in_wt_data_int16_58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1517" *)
  wire [15:0] in_wt_data_int16_59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1518" *)
  wire [15:0] in_wt_data_int16_6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1519" *)
  wire [15:0] in_wt_data_int16_60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1520" *)
  wire [15:0] in_wt_data_int16_61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1521" *)
  wire [15:0] in_wt_data_int16_62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1522" *)
  wire [15:0] in_wt_data_int16_63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1523" *)
  wire [15:0] in_wt_data_int16_7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1524" *)
  wire [15:0] in_wt_data_int16_8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1525" *)
  wire [15:0] in_wt_data_int16_9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1526" *)
  wire [1023:0] in_wt_data_int8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1527" *)
  wire [15:0] in_wt_data_int8_0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1528" *)
  wire [15:0] in_wt_data_int8_1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1529" *)
  wire [15:0] in_wt_data_int8_10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1530" *)
  wire [15:0] in_wt_data_int8_11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1531" *)
  wire [15:0] in_wt_data_int8_12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1532" *)
  wire [15:0] in_wt_data_int8_13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1533" *)
  wire [15:0] in_wt_data_int8_14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1534" *)
  wire [15:0] in_wt_data_int8_15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1535" *)
  wire [15:0] in_wt_data_int8_16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1536" *)
  wire [15:0] in_wt_data_int8_17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1537" *)
  wire [15:0] in_wt_data_int8_18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1538" *)
  wire [15:0] in_wt_data_int8_19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1539" *)
  wire [15:0] in_wt_data_int8_2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1540" *)
  wire [15:0] in_wt_data_int8_20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1541" *)
  wire [15:0] in_wt_data_int8_21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1542" *)
  wire [15:0] in_wt_data_int8_22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1543" *)
  wire [15:0] in_wt_data_int8_23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1544" *)
  wire [15:0] in_wt_data_int8_24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1545" *)
  wire [15:0] in_wt_data_int8_25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1546" *)
  wire [15:0] in_wt_data_int8_26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1547" *)
  wire [15:0] in_wt_data_int8_27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1548" *)
  wire [15:0] in_wt_data_int8_28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1549" *)
  wire [15:0] in_wt_data_int8_29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1550" *)
  wire [15:0] in_wt_data_int8_3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1551" *)
  wire [15:0] in_wt_data_int8_30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1552" *)
  wire [15:0] in_wt_data_int8_31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1553" *)
  wire [15:0] in_wt_data_int8_32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1554" *)
  wire [15:0] in_wt_data_int8_33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1555" *)
  wire [15:0] in_wt_data_int8_34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1556" *)
  wire [15:0] in_wt_data_int8_35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1557" *)
  wire [15:0] in_wt_data_int8_36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1558" *)
  wire [15:0] in_wt_data_int8_37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1559" *)
  wire [15:0] in_wt_data_int8_38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1560" *)
  wire [15:0] in_wt_data_int8_39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1561" *)
  wire [15:0] in_wt_data_int8_4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1562" *)
  wire [15:0] in_wt_data_int8_40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1563" *)
  wire [15:0] in_wt_data_int8_41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1564" *)
  wire [15:0] in_wt_data_int8_42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1565" *)
  wire [15:0] in_wt_data_int8_43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1566" *)
  wire [15:0] in_wt_data_int8_44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1567" *)
  wire [15:0] in_wt_data_int8_45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1568" *)
  wire [15:0] in_wt_data_int8_46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1569" *)
  wire [15:0] in_wt_data_int8_47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1570" *)
  wire [15:0] in_wt_data_int8_48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1571" *)
  wire [15:0] in_wt_data_int8_49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1572" *)
  wire [15:0] in_wt_data_int8_5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1573" *)
  wire [15:0] in_wt_data_int8_50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1574" *)
  wire [15:0] in_wt_data_int8_51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1575" *)
  wire [15:0] in_wt_data_int8_52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1576" *)
  wire [15:0] in_wt_data_int8_53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1577" *)
  wire [15:0] in_wt_data_int8_54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1578" *)
  wire [15:0] in_wt_data_int8_55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1579" *)
  wire [15:0] in_wt_data_int8_56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1580" *)
  wire [15:0] in_wt_data_int8_57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1581" *)
  wire [15:0] in_wt_data_int8_58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1582" *)
  wire [15:0] in_wt_data_int8_59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1583" *)
  wire [15:0] in_wt_data_int8_6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1584" *)
  wire [15:0] in_wt_data_int8_60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1585" *)
  wire [15:0] in_wt_data_int8_61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1586" *)
  wire [15:0] in_wt_data_int8_62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1587" *)
  wire [15:0] in_wt_data_int8_63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1588" *)
  wire [15:0] in_wt_data_int8_7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1589" *)
  wire [15:0] in_wt_data_int8_8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1590" *)
  wire [15:0] in_wt_data_int8_9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1591" *)
  wire [1023:0] in_wt_data_pack;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1592" *)
  wire [191:0] in_wt_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:674" *)
  input [127:0] in_wt_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1593" *)
  wire [127:0] in_wt_mask_int8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1594" *)
  wire [63:0] in_wt_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1595" *)
  wire [63:0] in_wt_norm;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:675" *)
  input in_wt_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:676" *)
  input [7:0] in_wt_sel;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:408" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:409" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:749" *)
  output [1023:0] wt0_actv_data;
  reg [1023:0] wt0_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:750" *)
  output [63:0] wt0_actv_nan;
  reg [63:0] wt0_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:751" *)
  output [127:0] wt0_actv_nz;
  reg [127:0] wt0_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:752" *)
  output [103:0] wt0_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1600" *)
  wire wt0_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1601" *)
  wire wt0_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1602" *)
  reg [1023:0] wt0_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:753" *)
  output [191:0] wt0_sd_exp;
  reg [191:0] wt0_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:754" *)
  output [63:0] wt0_sd_mask;
  reg [63:0] wt0_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1605" *)
  reg [63:0] wt0_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1606" *)
  reg [127:0] wt0_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:755" *)
  output wt0_sd_pvld;
  reg wt0_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1608" *)
  wire wt0_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:756" *)
  output [1023:0] wt1_actv_data;
  reg [1023:0] wt1_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:757" *)
  output [63:0] wt1_actv_nan;
  reg [63:0] wt1_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:758" *)
  output [127:0] wt1_actv_nz;
  reg [127:0] wt1_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:759" *)
  output [103:0] wt1_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1613" *)
  wire wt1_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1614" *)
  wire wt1_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1615" *)
  reg [1023:0] wt1_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:760" *)
  output [191:0] wt1_sd_exp;
  reg [191:0] wt1_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:761" *)
  output [63:0] wt1_sd_mask;
  reg [63:0] wt1_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1618" *)
  reg [63:0] wt1_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1619" *)
  reg [127:0] wt1_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:762" *)
  output wt1_sd_pvld;
  reg wt1_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1621" *)
  wire wt1_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:763" *)
  output [1023:0] wt2_actv_data;
  reg [1023:0] wt2_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:764" *)
  output [63:0] wt2_actv_nan;
  reg [63:0] wt2_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:765" *)
  output [127:0] wt2_actv_nz;
  reg [127:0] wt2_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:766" *)
  output [103:0] wt2_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1626" *)
  wire wt2_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1627" *)
  wire wt2_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1628" *)
  reg [1023:0] wt2_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:767" *)
  output [191:0] wt2_sd_exp;
  reg [191:0] wt2_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:768" *)
  output [63:0] wt2_sd_mask;
  reg [63:0] wt2_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1631" *)
  reg [63:0] wt2_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1632" *)
  reg [127:0] wt2_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:769" *)
  output wt2_sd_pvld;
  reg wt2_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1634" *)
  wire wt2_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:770" *)
  output [1023:0] wt3_actv_data;
  reg [1023:0] wt3_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:771" *)
  output [63:0] wt3_actv_nan;
  reg [63:0] wt3_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:772" *)
  output [127:0] wt3_actv_nz;
  reg [127:0] wt3_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:773" *)
  output [103:0] wt3_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1639" *)
  wire wt3_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1640" *)
  wire wt3_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1641" *)
  reg [1023:0] wt3_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:774" *)
  output [191:0] wt3_sd_exp;
  reg [191:0] wt3_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:775" *)
  output [63:0] wt3_sd_mask;
  reg [63:0] wt3_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1644" *)
  reg [63:0] wt3_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1645" *)
  reg [127:0] wt3_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:776" *)
  output wt3_sd_pvld;
  reg wt3_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1647" *)
  wire wt3_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:777" *)
  output [1023:0] wt4_actv_data;
  reg [1023:0] wt4_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:778" *)
  output [63:0] wt4_actv_nan;
  reg [63:0] wt4_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:779" *)
  output [127:0] wt4_actv_nz;
  reg [127:0] wt4_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:780" *)
  output [103:0] wt4_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1652" *)
  wire wt4_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1653" *)
  wire wt4_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1654" *)
  reg [1023:0] wt4_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:781" *)
  output [191:0] wt4_sd_exp;
  reg [191:0] wt4_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:782" *)
  output [63:0] wt4_sd_mask;
  reg [63:0] wt4_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1657" *)
  reg [63:0] wt4_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1658" *)
  reg [127:0] wt4_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:783" *)
  output wt4_sd_pvld;
  reg wt4_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1660" *)
  wire wt4_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:784" *)
  output [1023:0] wt5_actv_data;
  reg [1023:0] wt5_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:785" *)
  output [63:0] wt5_actv_nan;
  reg [63:0] wt5_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:786" *)
  output [127:0] wt5_actv_nz;
  reg [127:0] wt5_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:787" *)
  output [103:0] wt5_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1665" *)
  wire wt5_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1666" *)
  wire wt5_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1667" *)
  reg [1023:0] wt5_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:788" *)
  output [191:0] wt5_sd_exp;
  reg [191:0] wt5_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:789" *)
  output [63:0] wt5_sd_mask;
  reg [63:0] wt5_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1670" *)
  reg [63:0] wt5_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1671" *)
  reg [127:0] wt5_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:790" *)
  output wt5_sd_pvld;
  reg wt5_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1673" *)
  wire wt5_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:791" *)
  output [1023:0] wt6_actv_data;
  reg [1023:0] wt6_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:792" *)
  output [63:0] wt6_actv_nan;
  reg [63:0] wt6_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:793" *)
  output [127:0] wt6_actv_nz;
  reg [127:0] wt6_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:794" *)
  output [103:0] wt6_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1678" *)
  wire wt6_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1679" *)
  wire wt6_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1680" *)
  reg [1023:0] wt6_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:795" *)
  output [191:0] wt6_sd_exp;
  reg [191:0] wt6_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:796" *)
  output [63:0] wt6_sd_mask;
  reg [63:0] wt6_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1683" *)
  reg [63:0] wt6_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1684" *)
  reg [127:0] wt6_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:797" *)
  output wt6_sd_pvld;
  reg wt6_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1686" *)
  wire wt6_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:798" *)
  output [1023:0] wt7_actv_data;
  reg [1023:0] wt7_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:799" *)
  output [63:0] wt7_actv_nan;
  reg [63:0] wt7_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:800" *)
  output [127:0] wt7_actv_nz;
  reg [127:0] wt7_actv_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:801" *)
  output [103:0] wt7_actv_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1691" *)
  wire wt7_actv_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1692" *)
  wire wt7_actv_vld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1693" *)
  reg [1023:0] wt7_sd_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:802" *)
  output [191:0] wt7_sd_exp;
  reg [191:0] wt7_sd_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:803" *)
  output [63:0] wt7_sd_mask;
  reg [63:0] wt7_sd_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1696" *)
  reg [63:0] wt7_sd_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1697" *)
  reg [127:0] wt7_sd_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:804" *)
  output wt7_sd_pvld;
  reg wt7_sd_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1699" *)
  wire wt7_sd_pvld_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1700" *)
  wire wt_has_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1701" *)
  reg [1023:0] wt_pre_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1702" *)
  wire [1023:0] wt_pre_data_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1703" *)
  reg [191:0] wt_pre_exp;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1704" *)
  wire [191:0] wt_pre_exp_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1705" *)
  reg [63:0] wt_pre_mask;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1706" *)
  wire [63:0] wt_pre_mask_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1707" *)
  reg [63:0] wt_pre_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1708" *)
  reg [127:0] wt_pre_nz;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1709" *)
  wire [127:0] wt_pre_nz_w;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1710" *)
  reg [7:0] wt_pre_sel;
  assign _03419_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10000" *) _06409_;
  assign _03420_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10010" *) _06410_;
  assign _03421_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10020" *) _06411_;
  assign _03422_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10030" *) _06412_;
  assign _03423_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10040" *) _06413_;
  assign _03424_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10050" *) _06414_;
  assign _03425_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10060" *) _06415_;
  assign _03426_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10070" *) _06416_;
  assign _03427_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10080" *) _06417_;
  assign _03428_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10090" *) _06418_;
  assign _03429_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10100" *) _06419_;
  assign _03430_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10110" *) _06420_;
  assign _03431_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10120" *) _06421_;
  assign _03432_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10130" *) _06422_;
  assign _03433_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10140" *) _06423_;
  assign _03434_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10150" *) _06424_;
  assign _03435_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10160" *) _06425_;
  assign _03436_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10170" *) _06426_;
  assign _03437_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10180" *) _06427_;
  assign _03438_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10190" *) _06428_;
  assign _03439_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10200" *) _06429_;
  assign _03440_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10210" *) _06430_;
  assign _03441_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10220" *) _06431_;
  assign _03442_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10230" *) _06432_;
  assign _03443_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10240" *) _06433_;
  assign _03444_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10250" *) _06434_;
  assign _03445_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10260" *) _06435_;
  assign _03446_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10270" *) _06436_;
  assign _03447_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10280" *) _06437_;
  assign _03448_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10290" *) _06438_;
  assign _03449_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10300" *) _06439_;
  assign _03450_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10310" *) _06440_;
  assign _03451_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10320" *) _06441_;
  assign _03452_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10330" *) _06442_;
  assign _03453_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10340" *) _06443_;
  assign _03454_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10350" *) _06444_;
  assign _03455_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10360" *) _06445_;
  assign _03456_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10370" *) _06446_;
  assign _03457_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10380" *) _06447_;
  assign _03458_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10390" *) _06448_;
  assign _03459_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10400" *) _06449_;
  assign _03460_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10410" *) _06450_;
  assign _03461_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10420" *) _06451_;
  assign _03462_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10430" *) _06452_;
  assign _03463_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10440" *) _06453_;
  assign _03464_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10450" *) _06454_;
  assign _03465_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10460" *) _06455_;
  assign _03466_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10470" *) _06456_;
  assign _03467_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10480" *) _06457_;
  assign _03468_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10490" *) _06458_;
  assign _03469_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10500" *) _06459_;
  assign _03470_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10510" *) _06460_;
  assign _03471_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10520" *) _06461_;
  assign _03472_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10530" *) _06462_;
  assign _03473_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10540" *) _06463_;
  assign _03474_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10550" *) _06464_;
  assign _03475_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10560" *) _06465_;
  assign _03476_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10570" *) _06466_;
  assign _03477_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10580" *) _06467_;
  assign _03478_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10590" *) _06468_;
  assign _03479_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10600" *) _06469_;
  assign _03480_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10610" *) _06470_;
  assign _03481_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10620" *) _06471_;
  assign _03482_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10630" *) _06472_;
  assign _03483_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10640" *) _06473_;
  assign _03484_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10650" *) _06474_;
  assign _03485_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10686" *) cfg_is_fp16_d1[70];
  assign _03486_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10716" *) _06475_;
  assign _03487_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10726" *) _06476_;
  assign _03488_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10736" *) _06477_;
  assign _03489_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10746" *) _06478_;
  assign _03490_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10756" *) _06479_;
  assign _03491_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10766" *) _06480_;
  assign _03492_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10776" *) _06481_;
  assign _03493_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10786" *) _06482_;
  assign _03494_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10796" *) _06483_;
  assign _03495_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10806" *) _06484_;
  assign _03496_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10816" *) _06485_;
  assign _03497_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10826" *) _06486_;
  assign _03498_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10836" *) _06487_;
  assign _03499_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10846" *) _06488_;
  assign _03500_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10856" *) _06489_;
  assign _03501_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10866" *) _06490_;
  assign _03502_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10876" *) _06491_;
  assign _03503_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10886" *) _06492_;
  assign _03504_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10896" *) _06493_;
  assign _03505_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10906" *) _06494_;
  assign _03506_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10916" *) _06495_;
  assign _03507_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10926" *) _06496_;
  assign _03508_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10936" *) _06497_;
  assign _03509_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10946" *) _06498_;
  assign _03510_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10956" *) _06499_;
  assign _03511_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10966" *) _06500_;
  assign _03512_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10976" *) _06501_;
  assign _03513_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10986" *) _06502_;
  assign _03514_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10996" *) _06503_;
  assign _03515_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11006" *) _06504_;
  assign _03516_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11016" *) _06505_;
  assign _03517_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11026" *) _06506_;
  assign _03518_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11036" *) _06507_;
  assign _03519_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11046" *) _06508_;
  assign _03520_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11056" *) _06509_;
  assign _03521_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11066" *) _06510_;
  assign _03522_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11076" *) _06511_;
  assign _03523_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11086" *) _06512_;
  assign _03524_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11096" *) _06513_;
  assign _03525_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11106" *) _06514_;
  assign _03526_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11116" *) _06515_;
  assign _03527_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11126" *) _06516_;
  assign _03528_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11136" *) _06517_;
  assign _03529_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11146" *) _06518_;
  assign _03530_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11156" *) _06519_;
  assign _03531_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11166" *) _06520_;
  assign _03532_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11176" *) _06521_;
  assign _03533_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11186" *) _06522_;
  assign _03534_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11196" *) _06523_;
  assign _03535_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11206" *) _06524_;
  assign _03536_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11216" *) _06525_;
  assign _03537_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11226" *) _06526_;
  assign _03538_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11236" *) _06527_;
  assign _03539_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11246" *) _06528_;
  assign _03540_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11256" *) _06529_;
  assign _03541_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11266" *) _06530_;
  assign _03542_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11276" *) _06531_;
  assign _03543_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11286" *) _06532_;
  assign _03544_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11296" *) _06533_;
  assign _03545_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11306" *) _06534_;
  assign _03546_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11316" *) _06535_;
  assign _03547_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11326" *) _06536_;
  assign _03548_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11336" *) _06409_;
  assign _03549_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11346" *) _06410_;
  assign _03550_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11356" *) _06411_;
  assign _03551_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11366" *) _06412_;
  assign _03552_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11376" *) _06413_;
  assign _03553_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11386" *) _06414_;
  assign _03554_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11396" *) _06415_;
  assign _03555_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11406" *) _06416_;
  assign _03556_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11416" *) _06417_;
  assign _03557_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11426" *) _06418_;
  assign _03558_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11436" *) _06419_;
  assign _03559_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11446" *) _06420_;
  assign _03560_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11456" *) _06421_;
  assign _03561_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11466" *) _06422_;
  assign _03562_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11476" *) _06423_;
  assign _03563_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11486" *) _06424_;
  assign _03564_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11496" *) _06425_;
  assign _03565_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11506" *) _06426_;
  assign _03566_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11516" *) _06427_;
  assign _03567_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11526" *) _06428_;
  assign _03568_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11536" *) _06429_;
  assign _03569_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11546" *) _06430_;
  assign _03570_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11556" *) _06431_;
  assign _03571_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11566" *) _06432_;
  assign _03572_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11576" *) _06433_;
  assign _03573_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11586" *) _06434_;
  assign _03574_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11596" *) _06435_;
  assign _03575_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11606" *) _06436_;
  assign _03576_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11616" *) _06437_;
  assign _03577_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11626" *) _06438_;
  assign _03578_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11636" *) _06439_;
  assign _03579_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11646" *) _06440_;
  assign _03580_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11656" *) _06441_;
  assign _03581_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11666" *) _06442_;
  assign _03582_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11676" *) _06443_;
  assign _03583_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11686" *) _06444_;
  assign _03584_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11696" *) _06445_;
  assign _03585_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11706" *) _06446_;
  assign _03586_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11716" *) _06447_;
  assign _03587_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11726" *) _06448_;
  assign _03588_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11736" *) _06449_;
  assign _03589_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11746" *) _06450_;
  assign _03590_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11756" *) _06451_;
  assign _03591_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11766" *) _06452_;
  assign _03592_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11776" *) _06453_;
  assign _03593_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11786" *) _06454_;
  assign _03594_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11796" *) _06455_;
  assign _03595_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11806" *) _06456_;
  assign _03596_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11816" *) _06457_;
  assign _03597_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11826" *) _06458_;
  assign _03598_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11836" *) _06459_;
  assign _03599_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11846" *) _06460_;
  assign _03600_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11856" *) _06461_;
  assign _03601_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11866" *) _06462_;
  assign _03602_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11876" *) _06463_;
  assign _03603_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11886" *) _06464_;
  assign _03604_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11896" *) _06465_;
  assign _03605_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11906" *) _06466_;
  assign _03606_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11916" *) _06467_;
  assign _03607_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11926" *) _06468_;
  assign _03608_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11936" *) _06469_;
  assign _03609_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11946" *) _06470_;
  assign _03610_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11956" *) _06471_;
  assign _03611_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11966" *) _06472_;
  assign _03612_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11976" *) _06473_;
  assign _03613_ = wt_pre_sel[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11986" *) _06474_;
  assign _03614_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12022" *) cfg_is_fp16_d1[71];
  assign _03615_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12052" *) _06475_;
  assign _03616_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12062" *) _06476_;
  assign _03617_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12072" *) _06477_;
  assign _03618_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12082" *) _06478_;
  assign _03619_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12092" *) _06479_;
  assign _03620_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12102" *) _06480_;
  assign _03621_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12112" *) _06481_;
  assign _03622_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12122" *) _06482_;
  assign _03623_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12132" *) _06483_;
  assign _03624_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12142" *) _06484_;
  assign _03625_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12152" *) _06485_;
  assign _03626_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12162" *) _06486_;
  assign _03627_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12172" *) _06487_;
  assign _03628_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12182" *) _06488_;
  assign _03629_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12192" *) _06489_;
  assign _03630_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12202" *) _06490_;
  assign _03631_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12212" *) _06491_;
  assign _03632_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12222" *) _06492_;
  assign _03633_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12232" *) _06493_;
  assign _03634_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12242" *) _06494_;
  assign _03635_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12252" *) _06495_;
  assign _03636_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12262" *) _06496_;
  assign _03637_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12272" *) _06497_;
  assign _03638_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12282" *) _06498_;
  assign _03639_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12292" *) _06499_;
  assign _03640_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12302" *) _06500_;
  assign _03641_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12312" *) _06501_;
  assign _03642_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12322" *) _06502_;
  assign _03643_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12332" *) _06503_;
  assign _03644_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12342" *) _06504_;
  assign _03645_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12352" *) _06505_;
  assign _03646_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12362" *) _06506_;
  assign _03647_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12372" *) _06507_;
  assign _03648_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12382" *) _06508_;
  assign _03649_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12392" *) _06509_;
  assign _03650_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12402" *) _06510_;
  assign _03651_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12412" *) _06511_;
  assign _03652_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12422" *) _06512_;
  assign _03653_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12432" *) _06513_;
  assign _03654_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12442" *) _06514_;
  assign _03655_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12452" *) _06515_;
  assign _03656_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12462" *) _06516_;
  assign _03657_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12472" *) _06517_;
  assign _03658_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12482" *) _06518_;
  assign _03659_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12492" *) _06519_;
  assign _03660_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12502" *) _06520_;
  assign _03661_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12512" *) _06521_;
  assign _03662_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12522" *) _06522_;
  assign _03663_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12532" *) _06523_;
  assign _03664_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12542" *) _06524_;
  assign _03665_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12552" *) _06525_;
  assign _03666_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12562" *) _06526_;
  assign _03667_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12572" *) _06527_;
  assign _03668_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12582" *) _06528_;
  assign _03669_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12592" *) _06529_;
  assign _03670_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12602" *) _06530_;
  assign _03671_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12612" *) _06531_;
  assign _03672_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12622" *) _06532_;
  assign _03673_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12632" *) _06533_;
  assign _03674_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12642" *) _06534_;
  assign _03675_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12652" *) _06535_;
  assign _03676_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12662" *) _06536_;
  assign _03677_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12672" *) _06409_;
  assign _03678_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12682" *) _06410_;
  assign _03679_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12692" *) _06411_;
  assign _03680_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12702" *) _06412_;
  assign _03681_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12712" *) _06413_;
  assign _03682_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12722" *) _06414_;
  assign _03683_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12732" *) _06415_;
  assign _03684_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12742" *) _06416_;
  assign _03685_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12752" *) _06417_;
  assign _03686_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12762" *) _06418_;
  assign _03687_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12772" *) _06419_;
  assign _03688_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12782" *) _06420_;
  assign _03689_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12792" *) _06421_;
  assign _03690_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12802" *) _06422_;
  assign _03691_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12812" *) _06423_;
  assign _03692_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12822" *) _06424_;
  assign _03693_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12832" *) _06425_;
  assign _03694_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12842" *) _06426_;
  assign _03695_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12852" *) _06427_;
  assign _03696_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12862" *) _06428_;
  assign _03697_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12872" *) _06429_;
  assign _03698_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12882" *) _06430_;
  assign _03699_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12892" *) _06431_;
  assign _03700_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12902" *) _06432_;
  assign _03701_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12912" *) _06433_;
  assign _03702_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12922" *) _06434_;
  assign _03703_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12932" *) _06435_;
  assign _03704_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12942" *) _06436_;
  assign _03705_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12952" *) _06437_;
  assign _03706_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12962" *) _06438_;
  assign _03707_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12972" *) _06439_;
  assign _03708_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12982" *) _06440_;
  assign _03709_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12992" *) _06441_;
  assign _03710_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13002" *) _06442_;
  assign _03711_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13012" *) _06443_;
  assign _03712_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13022" *) _06444_;
  assign _03713_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13032" *) _06445_;
  assign _03714_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13042" *) _06446_;
  assign _03715_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13052" *) _06447_;
  assign _03716_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13062" *) _06448_;
  assign _03717_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13072" *) _06449_;
  assign _03718_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13082" *) _06450_;
  assign _03719_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13092" *) _06451_;
  assign _03720_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13102" *) _06452_;
  assign _03721_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13112" *) _06453_;
  assign _03722_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13122" *) _06454_;
  assign _03723_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13132" *) _06455_;
  assign _03724_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13142" *) _06456_;
  assign _03725_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13152" *) _06457_;
  assign _03726_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13162" *) _06458_;
  assign _03727_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13172" *) _06459_;
  assign _03728_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13182" *) _06460_;
  assign _03729_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13192" *) _06461_;
  assign _03730_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13202" *) _06462_;
  assign _03731_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13212" *) _06463_;
  assign _03732_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13222" *) _06464_;
  assign _03733_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13232" *) _06465_;
  assign _03734_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13242" *) _06466_;
  assign _03735_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13252" *) _06467_;
  assign _03736_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13262" *) _06468_;
  assign _03737_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13272" *) _06469_;
  assign _03738_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13282" *) _06470_;
  assign _03739_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13292" *) _06471_;
  assign _03740_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13302" *) _06472_;
  assign _03741_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13312" *) _06473_;
  assign _03742_ = wt_pre_sel[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13322" *) _06474_;
  assign _03743_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13358" *) cfg_is_fp16_d1[72];
  assign _03744_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13388" *) _06475_;
  assign _03745_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13398" *) _06476_;
  assign _03746_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13408" *) _06477_;
  assign _03747_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13418" *) _06478_;
  assign _03748_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13428" *) _06479_;
  assign _03749_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13438" *) _06480_;
  assign _03750_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13448" *) _06481_;
  assign _03751_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13458" *) _06482_;
  assign _03752_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13468" *) _06483_;
  assign _03753_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13478" *) _06484_;
  assign _03754_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13488" *) _06485_;
  assign _03755_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13498" *) _06486_;
  assign _03756_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13508" *) _06487_;
  assign _03757_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13518" *) _06488_;
  assign _03758_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13528" *) _06489_;
  assign _03759_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13538" *) _06490_;
  assign _03760_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13548" *) _06491_;
  assign _03761_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13558" *) _06492_;
  assign _03762_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13568" *) _06493_;
  assign _03763_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13578" *) _06494_;
  assign _03764_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13588" *) _06495_;
  assign _03765_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13598" *) _06496_;
  assign _03766_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13608" *) _06497_;
  assign _03767_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13618" *) _06498_;
  assign _03768_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13628" *) _06499_;
  assign _03769_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13638" *) _06500_;
  assign _03770_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13648" *) _06501_;
  assign _03771_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13658" *) _06502_;
  assign _03772_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13668" *) _06503_;
  assign _03773_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13678" *) _06504_;
  assign _03774_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13688" *) _06505_;
  assign _03775_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13698" *) _06506_;
  assign _03776_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13708" *) _06507_;
  assign _03777_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13718" *) _06508_;
  assign _03778_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13728" *) _06509_;
  assign _03779_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13738" *) _06510_;
  assign _03780_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13748" *) _06511_;
  assign _03781_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13758" *) _06512_;
  assign _03782_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13768" *) _06513_;
  assign _03783_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13778" *) _06514_;
  assign _03784_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13788" *) _06515_;
  assign _03785_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13798" *) _06516_;
  assign _03786_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13808" *) _06517_;
  assign _03787_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13818" *) _06518_;
  assign _03788_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13828" *) _06519_;
  assign _03789_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13838" *) _06520_;
  assign _03790_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13848" *) _06521_;
  assign _03791_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13858" *) _06522_;
  assign _03792_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13868" *) _06523_;
  assign _03793_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13878" *) _06524_;
  assign _03794_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13888" *) _06525_;
  assign _03795_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13898" *) _06526_;
  assign _03796_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13908" *) _06527_;
  assign _03797_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13918" *) _06528_;
  assign _03798_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13928" *) _06529_;
  assign _03799_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13938" *) _06530_;
  assign _03800_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13948" *) _06531_;
  assign _03801_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13958" *) _06532_;
  assign _03802_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13968" *) _06533_;
  assign _03803_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13978" *) _06534_;
  assign _03804_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13988" *) _06535_;
  assign _03805_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13998" *) _06536_;
  assign _03806_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14008" *) _06409_;
  assign _03807_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14018" *) _06410_;
  assign _03808_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14028" *) _06411_;
  assign _03809_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14038" *) _06412_;
  assign _03810_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14048" *) _06413_;
  assign _03811_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14058" *) _06414_;
  assign _03812_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14068" *) _06415_;
  assign _03813_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14078" *) _06416_;
  assign _03814_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14088" *) _06417_;
  assign _03815_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14098" *) _06418_;
  assign _03816_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14108" *) _06419_;
  assign _03817_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14118" *) _06420_;
  assign _03818_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14128" *) _06421_;
  assign _03819_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14138" *) _06422_;
  assign _03820_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14148" *) _06423_;
  assign _03821_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14158" *) _06424_;
  assign _03822_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14168" *) _06425_;
  assign _03823_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14178" *) _06426_;
  assign _03824_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14188" *) _06427_;
  assign _03825_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14198" *) _06428_;
  assign _03826_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14208" *) _06429_;
  assign _03827_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14218" *) _06430_;
  assign _03828_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14228" *) _06431_;
  assign _03829_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14238" *) _06432_;
  assign _03830_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14248" *) _06433_;
  assign _03831_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14258" *) _06434_;
  assign _03832_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14268" *) _06435_;
  assign _03833_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14278" *) _06436_;
  assign _03834_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14288" *) _06437_;
  assign _03835_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14298" *) _06438_;
  assign _03836_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14308" *) _06439_;
  assign _03837_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14318" *) _06440_;
  assign _03838_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14328" *) _06441_;
  assign _03839_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14338" *) _06442_;
  assign _03840_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14348" *) _06443_;
  assign _03841_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14358" *) _06444_;
  assign _03842_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14368" *) _06445_;
  assign _03843_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14378" *) _06446_;
  assign _03844_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14388" *) _06447_;
  assign _03845_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14398" *) _06448_;
  assign _03846_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14408" *) _06449_;
  assign _03847_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14418" *) _06450_;
  assign _03848_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14428" *) _06451_;
  assign _03849_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14438" *) _06452_;
  assign _03850_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14448" *) _06453_;
  assign _03851_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14458" *) _06454_;
  assign _03852_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14468" *) _06455_;
  assign _03853_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14478" *) _06456_;
  assign _03854_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14488" *) _06457_;
  assign _03855_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14498" *) _06458_;
  assign _03856_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14508" *) _06459_;
  assign _03857_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14518" *) _06460_;
  assign _03858_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14528" *) _06461_;
  assign _03859_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14538" *) _06462_;
  assign _03860_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14548" *) _06463_;
  assign _03861_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14558" *) _06464_;
  assign _03862_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14568" *) _06465_;
  assign _03863_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14578" *) _06466_;
  assign _03864_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14588" *) _06467_;
  assign _03865_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14598" *) _06468_;
  assign _03866_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14608" *) _06469_;
  assign _03867_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14618" *) _06470_;
  assign _03868_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14628" *) _06471_;
  assign _03869_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14638" *) _06472_;
  assign _03870_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14648" *) _06473_;
  assign _03871_ = wt_pre_sel[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14658" *) _06474_;
  assign _03872_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14694" *) cfg_is_fp16_d1[73];
  assign _03873_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14724" *) _06475_;
  assign _03874_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14734" *) _06476_;
  assign _03875_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14744" *) _06477_;
  assign _03876_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14754" *) _06478_;
  assign _03877_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14764" *) _06479_;
  assign _03878_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14774" *) _06480_;
  assign _03879_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14784" *) _06481_;
  assign _03880_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14794" *) _06482_;
  assign _03881_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14804" *) _06483_;
  assign _03882_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14814" *) _06484_;
  assign _03883_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14824" *) _06485_;
  assign _03884_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14834" *) _06486_;
  assign _03885_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14844" *) _06487_;
  assign _03886_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14854" *) _06488_;
  assign _03887_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14864" *) _06489_;
  assign _03888_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14874" *) _06490_;
  assign _03889_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14884" *) _06491_;
  assign _03890_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14894" *) _06492_;
  assign _03891_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14904" *) _06493_;
  assign _03892_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14914" *) _06494_;
  assign _03893_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14924" *) _06495_;
  assign _03894_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14934" *) _06496_;
  assign _03895_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14944" *) _06497_;
  assign _03896_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14954" *) _06498_;
  assign _03897_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14964" *) _06499_;
  assign _03898_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14974" *) _06500_;
  assign _03899_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14984" *) _06501_;
  assign _03900_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14994" *) _06502_;
  assign _03901_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15004" *) _06503_;
  assign _03902_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15014" *) _06504_;
  assign _03903_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15024" *) _06505_;
  assign _03904_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15034" *) _06506_;
  assign _03905_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15044" *) _06507_;
  assign _03906_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15054" *) _06508_;
  assign _03907_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15064" *) _06509_;
  assign _03908_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15074" *) _06510_;
  assign _03909_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15084" *) _06511_;
  assign _03910_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15094" *) _06512_;
  assign _03911_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15104" *) _06513_;
  assign _03912_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15114" *) _06514_;
  assign _03913_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15124" *) _06515_;
  assign _03914_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15134" *) _06516_;
  assign _03915_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15144" *) _06517_;
  assign _03916_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15154" *) _06518_;
  assign _03917_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15164" *) _06519_;
  assign _03918_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15174" *) _06520_;
  assign _03919_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15184" *) _06521_;
  assign _03920_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15194" *) _06522_;
  assign _03921_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15204" *) _06523_;
  assign _03922_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15214" *) _06524_;
  assign _03923_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15224" *) _06525_;
  assign _03924_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15234" *) _06526_;
  assign _03925_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15244" *) _06527_;
  assign _03926_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15254" *) _06528_;
  assign _03927_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15264" *) _06529_;
  assign _03928_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15274" *) _06530_;
  assign _03929_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15284" *) _06531_;
  assign _03930_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15294" *) _06532_;
  assign _03931_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15304" *) _06533_;
  assign _03932_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15314" *) _06534_;
  assign _03933_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15324" *) _06535_;
  assign _03934_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15334" *) _06536_;
  assign _03935_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15344" *) _06409_;
  assign _03936_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15354" *) _06410_;
  assign _03937_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15364" *) _06411_;
  assign _03938_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15374" *) _06412_;
  assign _03939_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15384" *) _06413_;
  assign _03940_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15394" *) _06414_;
  assign _03941_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15404" *) _06415_;
  assign _03942_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15414" *) _06416_;
  assign _03943_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15424" *) _06417_;
  assign _03944_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15434" *) _06418_;
  assign _03945_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15444" *) _06419_;
  assign _03946_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15454" *) _06420_;
  assign _03947_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15464" *) _06421_;
  assign _03948_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15474" *) _06422_;
  assign _03949_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15484" *) _06423_;
  assign _03950_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15494" *) _06424_;
  assign _03951_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15504" *) _06425_;
  assign _03952_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15514" *) _06426_;
  assign _03953_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15524" *) _06427_;
  assign _03954_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15534" *) _06428_;
  assign _03955_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15544" *) _06429_;
  assign _03956_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15554" *) _06430_;
  assign _03957_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15564" *) _06431_;
  assign _03958_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15574" *) _06432_;
  assign _03959_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15584" *) _06433_;
  assign _03960_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15594" *) _06434_;
  assign _03961_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15604" *) _06435_;
  assign _03962_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15614" *) _06436_;
  assign _03963_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15624" *) _06437_;
  assign _03964_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15634" *) _06438_;
  assign _03965_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15644" *) _06439_;
  assign _03966_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15654" *) _06440_;
  assign _03967_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15664" *) _06441_;
  assign _03968_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15674" *) _06442_;
  assign _03969_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15684" *) _06443_;
  assign _03970_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15694" *) _06444_;
  assign _03971_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15704" *) _06445_;
  assign _03972_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15714" *) _06446_;
  assign _03973_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15724" *) _06447_;
  assign _03974_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15734" *) _06448_;
  assign _03975_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15744" *) _06449_;
  assign _03976_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15754" *) _06450_;
  assign _03977_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15764" *) _06451_;
  assign _03978_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15774" *) _06452_;
  assign _03979_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15784" *) _06453_;
  assign _03980_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15794" *) _06454_;
  assign _03981_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15804" *) _06455_;
  assign _03982_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15814" *) _06456_;
  assign _03983_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15824" *) _06457_;
  assign _03984_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15834" *) _06458_;
  assign _03985_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15844" *) _06459_;
  assign _03986_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15854" *) _06460_;
  assign _03987_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15864" *) _06461_;
  assign _03988_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15874" *) _06462_;
  assign _03989_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15884" *) _06463_;
  assign _03990_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15894" *) _06464_;
  assign _03991_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15904" *) _06465_;
  assign _03992_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15914" *) _06466_;
  assign _03993_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15924" *) _06467_;
  assign _03994_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15934" *) _06468_;
  assign _03995_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15944" *) _06469_;
  assign _03996_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15954" *) _06470_;
  assign _03997_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15964" *) _06471_;
  assign _03998_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15974" *) _06472_;
  assign _03999_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15984" *) _06473_;
  assign _04000_ = wt_pre_sel[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15994" *) _06474_;
  assign _04001_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16028" *) wt0_actv_pvld_w;
  assign _04002_ = _04001_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16038" *) cfg_is_fp16_d1[74];
  assign _04003_ = { _06537_, _06537_, _06537_, _06537_, _06537_, _06537_, _06537_, _06537_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16049" *) wt0_sd_data[7:0];
  assign _04004_ = { _06538_, _06538_, _06538_, _06538_, _06538_, _06538_, _06538_, _06538_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16059" *) wt0_sd_data[15:8];
  assign _04005_ = { _06539_, _06539_, _06539_, _06539_, _06539_, _06539_, _06539_, _06539_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16069" *) wt0_sd_data[23:16];
  assign _04006_ = { _06540_, _06540_, _06540_, _06540_, _06540_, _06540_, _06540_, _06540_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16079" *) wt0_sd_data[31:24];
  assign _04007_ = { _06541_, _06541_, _06541_, _06541_, _06541_, _06541_, _06541_, _06541_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16089" *) wt0_sd_data[39:32];
  assign _04008_ = { _06542_, _06542_, _06542_, _06542_, _06542_, _06542_, _06542_, _06542_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16099" *) wt0_sd_data[47:40];
  assign _04009_ = { _06543_, _06543_, _06543_, _06543_, _06543_, _06543_, _06543_, _06543_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16109" *) wt0_sd_data[55:48];
  assign _04010_ = { _06544_, _06544_, _06544_, _06544_, _06544_, _06544_, _06544_, _06544_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16119" *) wt0_sd_data[63:56];
  assign _04011_ = { _06545_, _06545_, _06545_, _06545_, _06545_, _06545_, _06545_, _06545_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16129" *) wt0_sd_data[71:64];
  assign _04012_ = { _06546_, _06546_, _06546_, _06546_, _06546_, _06546_, _06546_, _06546_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16139" *) wt0_sd_data[79:72];
  assign _04013_ = { _06547_, _06547_, _06547_, _06547_, _06547_, _06547_, _06547_, _06547_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16149" *) wt0_sd_data[87:80];
  assign _04014_ = { _06548_, _06548_, _06548_, _06548_, _06548_, _06548_, _06548_, _06548_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16159" *) wt0_sd_data[95:88];
  assign _04015_ = { _06549_, _06549_, _06549_, _06549_, _06549_, _06549_, _06549_, _06549_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16169" *) wt0_sd_data[103:96];
  assign _04016_ = { _06550_, _06550_, _06550_, _06550_, _06550_, _06550_, _06550_, _06550_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16179" *) wt0_sd_data[111:104];
  assign _04017_ = { _06551_, _06551_, _06551_, _06551_, _06551_, _06551_, _06551_, _06551_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16189" *) wt0_sd_data[119:112];
  assign _04018_ = { _06552_, _06552_, _06552_, _06552_, _06552_, _06552_, _06552_, _06552_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16199" *) wt0_sd_data[127:120];
  assign _04019_ = { _06553_, _06553_, _06553_, _06553_, _06553_, _06553_, _06553_, _06553_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16209" *) wt0_sd_data[135:128];
  assign _04020_ = { _06554_, _06554_, _06554_, _06554_, _06554_, _06554_, _06554_, _06554_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16219" *) wt0_sd_data[143:136];
  assign _04021_ = { _06555_, _06555_, _06555_, _06555_, _06555_, _06555_, _06555_, _06555_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16229" *) wt0_sd_data[151:144];
  assign _04022_ = { _06556_, _06556_, _06556_, _06556_, _06556_, _06556_, _06556_, _06556_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16239" *) wt0_sd_data[159:152];
  assign _04023_ = { _06557_, _06557_, _06557_, _06557_, _06557_, _06557_, _06557_, _06557_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16249" *) wt0_sd_data[167:160];
  assign _04024_ = { _06558_, _06558_, _06558_, _06558_, _06558_, _06558_, _06558_, _06558_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16259" *) wt0_sd_data[175:168];
  assign _04025_ = { _06559_, _06559_, _06559_, _06559_, _06559_, _06559_, _06559_, _06559_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16269" *) wt0_sd_data[183:176];
  assign _04026_ = { _06560_, _06560_, _06560_, _06560_, _06560_, _06560_, _06560_, _06560_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16279" *) wt0_sd_data[191:184];
  assign _04027_ = { _06561_, _06561_, _06561_, _06561_, _06561_, _06561_, _06561_, _06561_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16289" *) wt0_sd_data[199:192];
  assign _04028_ = { _06562_, _06562_, _06562_, _06562_, _06562_, _06562_, _06562_, _06562_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16299" *) wt0_sd_data[207:200];
  assign _04029_ = { _06563_, _06563_, _06563_, _06563_, _06563_, _06563_, _06563_, _06563_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16309" *) wt0_sd_data[215:208];
  assign _04030_ = { _06564_, _06564_, _06564_, _06564_, _06564_, _06564_, _06564_, _06564_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16319" *) wt0_sd_data[223:216];
  assign _04031_ = { _06565_, _06565_, _06565_, _06565_, _06565_, _06565_, _06565_, _06565_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16329" *) wt0_sd_data[231:224];
  assign _04032_ = { _06566_, _06566_, _06566_, _06566_, _06566_, _06566_, _06566_, _06566_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16339" *) wt0_sd_data[239:232];
  assign _04033_ = { _06567_, _06567_, _06567_, _06567_, _06567_, _06567_, _06567_, _06567_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16349" *) wt0_sd_data[247:240];
  assign _04034_ = { _06568_, _06568_, _06568_, _06568_, _06568_, _06568_, _06568_, _06568_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16359" *) wt0_sd_data[255:248];
  assign _04035_ = { _06569_, _06569_, _06569_, _06569_, _06569_, _06569_, _06569_, _06569_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16369" *) wt0_sd_data[263:256];
  assign _04036_ = { _06570_, _06570_, _06570_, _06570_, _06570_, _06570_, _06570_, _06570_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16379" *) wt0_sd_data[271:264];
  assign _04037_ = { _06571_, _06571_, _06571_, _06571_, _06571_, _06571_, _06571_, _06571_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16389" *) wt0_sd_data[279:272];
  assign _04038_ = { _06572_, _06572_, _06572_, _06572_, _06572_, _06572_, _06572_, _06572_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16399" *) wt0_sd_data[287:280];
  assign _04039_ = { _06573_, _06573_, _06573_, _06573_, _06573_, _06573_, _06573_, _06573_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16409" *) wt0_sd_data[295:288];
  assign _04040_ = { _06574_, _06574_, _06574_, _06574_, _06574_, _06574_, _06574_, _06574_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16419" *) wt0_sd_data[303:296];
  assign _04041_ = { _06575_, _06575_, _06575_, _06575_, _06575_, _06575_, _06575_, _06575_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16429" *) wt0_sd_data[311:304];
  assign _04042_ = { _06576_, _06576_, _06576_, _06576_, _06576_, _06576_, _06576_, _06576_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16439" *) wt0_sd_data[319:312];
  assign _04043_ = { _06577_, _06577_, _06577_, _06577_, _06577_, _06577_, _06577_, _06577_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16449" *) wt0_sd_data[327:320];
  assign _04044_ = { _06578_, _06578_, _06578_, _06578_, _06578_, _06578_, _06578_, _06578_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16459" *) wt0_sd_data[335:328];
  assign _04045_ = { _06579_, _06579_, _06579_, _06579_, _06579_, _06579_, _06579_, _06579_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16469" *) wt0_sd_data[343:336];
  assign _04046_ = { _06580_, _06580_, _06580_, _06580_, _06580_, _06580_, _06580_, _06580_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16479" *) wt0_sd_data[351:344];
  assign _04047_ = { _06581_, _06581_, _06581_, _06581_, _06581_, _06581_, _06581_, _06581_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16489" *) wt0_sd_data[359:352];
  assign _04048_ = { _06582_, _06582_, _06582_, _06582_, _06582_, _06582_, _06582_, _06582_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16499" *) wt0_sd_data[367:360];
  assign _04049_ = { _06583_, _06583_, _06583_, _06583_, _06583_, _06583_, _06583_, _06583_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16509" *) wt0_sd_data[375:368];
  assign _04050_ = { _06584_, _06584_, _06584_, _06584_, _06584_, _06584_, _06584_, _06584_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16519" *) wt0_sd_data[383:376];
  assign _04051_ = { _06585_, _06585_, _06585_, _06585_, _06585_, _06585_, _06585_, _06585_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16529" *) wt0_sd_data[391:384];
  assign _04052_ = { _06586_, _06586_, _06586_, _06586_, _06586_, _06586_, _06586_, _06586_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16539" *) wt0_sd_data[399:392];
  assign _04053_ = { _06587_, _06587_, _06587_, _06587_, _06587_, _06587_, _06587_, _06587_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16549" *) wt0_sd_data[407:400];
  assign _04054_ = { _06588_, _06588_, _06588_, _06588_, _06588_, _06588_, _06588_, _06588_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16559" *) wt0_sd_data[415:408];
  assign _04055_ = { _06589_, _06589_, _06589_, _06589_, _06589_, _06589_, _06589_, _06589_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16569" *) wt0_sd_data[423:416];
  assign _04056_ = { _06590_, _06590_, _06590_, _06590_, _06590_, _06590_, _06590_, _06590_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16579" *) wt0_sd_data[431:424];
  assign _04057_ = { _06591_, _06591_, _06591_, _06591_, _06591_, _06591_, _06591_, _06591_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16589" *) wt0_sd_data[439:432];
  assign _04058_ = { _06592_, _06592_, _06592_, _06592_, _06592_, _06592_, _06592_, _06592_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16599" *) wt0_sd_data[447:440];
  assign _04059_ = { _06593_, _06593_, _06593_, _06593_, _06593_, _06593_, _06593_, _06593_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16609" *) wt0_sd_data[455:448];
  assign _04060_ = { _06594_, _06594_, _06594_, _06594_, _06594_, _06594_, _06594_, _06594_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16619" *) wt0_sd_data[463:456];
  assign _04061_ = { _06595_, _06595_, _06595_, _06595_, _06595_, _06595_, _06595_, _06595_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16629" *) wt0_sd_data[471:464];
  assign _04062_ = { _06596_, _06596_, _06596_, _06596_, _06596_, _06596_, _06596_, _06596_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16639" *) wt0_sd_data[479:472];
  assign _04063_ = { _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16649" *) wt0_sd_data[487:480];
  assign _04064_ = { _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16659" *) wt0_sd_data[495:488];
  assign _04065_ = { _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16669" *) wt0_sd_data[503:496];
  assign _04066_ = { _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16679" *) wt0_sd_data[511:504];
  assign _04067_ = { _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16689" *) wt0_sd_data[519:512];
  assign _04068_ = { _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16699" *) wt0_sd_data[527:520];
  assign _04069_ = { _06603_, _06603_, _06603_, _06603_, _06603_, _06603_, _06603_, _06603_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16709" *) wt0_sd_data[535:528];
  assign _04070_ = { _06604_, _06604_, _06604_, _06604_, _06604_, _06604_, _06604_, _06604_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16719" *) wt0_sd_data[543:536];
  assign _04071_ = { _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16729" *) wt0_sd_data[551:544];
  assign _04072_ = { _06606_, _06606_, _06606_, _06606_, _06606_, _06606_, _06606_, _06606_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16739" *) wt0_sd_data[559:552];
  assign _04073_ = { _06607_, _06607_, _06607_, _06607_, _06607_, _06607_, _06607_, _06607_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16749" *) wt0_sd_data[567:560];
  assign _04074_ = { _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16759" *) wt0_sd_data[575:568];
  assign _04075_ = { _06609_, _06609_, _06609_, _06609_, _06609_, _06609_, _06609_, _06609_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16769" *) wt0_sd_data[583:576];
  assign _04076_ = { _06610_, _06610_, _06610_, _06610_, _06610_, _06610_, _06610_, _06610_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16779" *) wt0_sd_data[591:584];
  assign _04077_ = { _06611_, _06611_, _06611_, _06611_, _06611_, _06611_, _06611_, _06611_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16789" *) wt0_sd_data[599:592];
  assign _04078_ = { _06612_, _06612_, _06612_, _06612_, _06612_, _06612_, _06612_, _06612_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16799" *) wt0_sd_data[607:600];
  assign _04079_ = { _06613_, _06613_, _06613_, _06613_, _06613_, _06613_, _06613_, _06613_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16809" *) wt0_sd_data[615:608];
  assign _04080_ = { _06614_, _06614_, _06614_, _06614_, _06614_, _06614_, _06614_, _06614_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16819" *) wt0_sd_data[623:616];
  assign _04081_ = { _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16829" *) wt0_sd_data[631:624];
  assign _04082_ = { _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16839" *) wt0_sd_data[639:632];
  assign _04083_ = { _06617_, _06617_, _06617_, _06617_, _06617_, _06617_, _06617_, _06617_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16849" *) wt0_sd_data[647:640];
  assign _04084_ = { _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16859" *) wt0_sd_data[655:648];
  assign _04085_ = { _06619_, _06619_, _06619_, _06619_, _06619_, _06619_, _06619_, _06619_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16869" *) wt0_sd_data[663:656];
  assign _04086_ = { _06620_, _06620_, _06620_, _06620_, _06620_, _06620_, _06620_, _06620_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16879" *) wt0_sd_data[671:664];
  assign _04087_ = { _06621_, _06621_, _06621_, _06621_, _06621_, _06621_, _06621_, _06621_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16889" *) wt0_sd_data[679:672];
  assign _04088_ = { _06622_, _06622_, _06622_, _06622_, _06622_, _06622_, _06622_, _06622_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16899" *) wt0_sd_data[687:680];
  assign _04089_ = { _06623_, _06623_, _06623_, _06623_, _06623_, _06623_, _06623_, _06623_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16909" *) wt0_sd_data[695:688];
  assign _04090_ = { _06624_, _06624_, _06624_, _06624_, _06624_, _06624_, _06624_, _06624_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16919" *) wt0_sd_data[703:696];
  assign _04091_ = { _06625_, _06625_, _06625_, _06625_, _06625_, _06625_, _06625_, _06625_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16929" *) wt0_sd_data[711:704];
  assign _04092_ = { _06626_, _06626_, _06626_, _06626_, _06626_, _06626_, _06626_, _06626_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16939" *) wt0_sd_data[719:712];
  assign _04093_ = { _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16949" *) wt0_sd_data[727:720];
  assign _04094_ = { _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16959" *) wt0_sd_data[735:728];
  assign _04095_ = { _06629_, _06629_, _06629_, _06629_, _06629_, _06629_, _06629_, _06629_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16969" *) wt0_sd_data[743:736];
  assign _04096_ = { _06630_, _06630_, _06630_, _06630_, _06630_, _06630_, _06630_, _06630_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16979" *) wt0_sd_data[751:744];
  assign _04097_ = { _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16989" *) wt0_sd_data[759:752];
  assign _04098_ = { _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16999" *) wt0_sd_data[767:760];
  assign _04099_ = { _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17009" *) wt0_sd_data[775:768];
  assign _04100_ = { _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17019" *) wt0_sd_data[783:776];
  assign _04101_ = { _06635_, _06635_, _06635_, _06635_, _06635_, _06635_, _06635_, _06635_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17029" *) wt0_sd_data[791:784];
  assign _04102_ = { _06636_, _06636_, _06636_, _06636_, _06636_, _06636_, _06636_, _06636_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17039" *) wt0_sd_data[799:792];
  assign _04103_ = { _06637_, _06637_, _06637_, _06637_, _06637_, _06637_, _06637_, _06637_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17049" *) wt0_sd_data[807:800];
  assign _04104_ = { _06638_, _06638_, _06638_, _06638_, _06638_, _06638_, _06638_, _06638_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17059" *) wt0_sd_data[815:808];
  assign _04105_ = { _06639_, _06639_, _06639_, _06639_, _06639_, _06639_, _06639_, _06639_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17069" *) wt0_sd_data[823:816];
  assign _04106_ = { _06640_, _06640_, _06640_, _06640_, _06640_, _06640_, _06640_, _06640_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17079" *) wt0_sd_data[831:824];
  assign _04107_ = { _06641_, _06641_, _06641_, _06641_, _06641_, _06641_, _06641_, _06641_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17089" *) wt0_sd_data[839:832];
  assign _04108_ = { _06642_, _06642_, _06642_, _06642_, _06642_, _06642_, _06642_, _06642_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17099" *) wt0_sd_data[847:840];
  assign _04109_ = { _06643_, _06643_, _06643_, _06643_, _06643_, _06643_, _06643_, _06643_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17109" *) wt0_sd_data[855:848];
  assign _04110_ = { _06644_, _06644_, _06644_, _06644_, _06644_, _06644_, _06644_, _06644_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17119" *) wt0_sd_data[863:856];
  assign _04111_ = { _06645_, _06645_, _06645_, _06645_, _06645_, _06645_, _06645_, _06645_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17129" *) wt0_sd_data[871:864];
  assign _04112_ = { _06646_, _06646_, _06646_, _06646_, _06646_, _06646_, _06646_, _06646_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17139" *) wt0_sd_data[879:872];
  assign _04113_ = { _06647_, _06647_, _06647_, _06647_, _06647_, _06647_, _06647_, _06647_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17149" *) wt0_sd_data[887:880];
  assign _04114_ = { _06648_, _06648_, _06648_, _06648_, _06648_, _06648_, _06648_, _06648_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17159" *) wt0_sd_data[895:888];
  assign _04115_ = { _06649_, _06649_, _06649_, _06649_, _06649_, _06649_, _06649_, _06649_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17169" *) wt0_sd_data[903:896];
  assign _04116_ = { _06650_, _06650_, _06650_, _06650_, _06650_, _06650_, _06650_, _06650_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17179" *) wt0_sd_data[911:904];
  assign _04117_ = { _06651_, _06651_, _06651_, _06651_, _06651_, _06651_, _06651_, _06651_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17189" *) wt0_sd_data[919:912];
  assign _04118_ = { _06652_, _06652_, _06652_, _06652_, _06652_, _06652_, _06652_, _06652_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17199" *) wt0_sd_data[927:920];
  assign _04119_ = { _06653_, _06653_, _06653_, _06653_, _06653_, _06653_, _06653_, _06653_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17209" *) wt0_sd_data[935:928];
  assign _04120_ = { _06654_, _06654_, _06654_, _06654_, _06654_, _06654_, _06654_, _06654_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17219" *) wt0_sd_data[943:936];
  assign _04121_ = { _06655_, _06655_, _06655_, _06655_, _06655_, _06655_, _06655_, _06655_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17229" *) wt0_sd_data[951:944];
  assign _04122_ = { _06656_, _06656_, _06656_, _06656_, _06656_, _06656_, _06656_, _06656_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17239" *) wt0_sd_data[959:952];
  assign _04123_ = { _06657_, _06657_, _06657_, _06657_, _06657_, _06657_, _06657_, _06657_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17249" *) wt0_sd_data[967:960];
  assign _04124_ = { _06658_, _06658_, _06658_, _06658_, _06658_, _06658_, _06658_, _06658_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17259" *) wt0_sd_data[975:968];
  assign _04125_ = { _06659_, _06659_, _06659_, _06659_, _06659_, _06659_, _06659_, _06659_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17269" *) wt0_sd_data[983:976];
  assign _04126_ = { _06660_, _06660_, _06660_, _06660_, _06660_, _06660_, _06660_, _06660_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17279" *) wt0_sd_data[991:984];
  assign _04127_ = { _06661_, _06661_, _06661_, _06661_, _06661_, _06661_, _06661_, _06661_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17289" *) wt0_sd_data[999:992];
  assign _04128_ = { _06662_, _06662_, _06662_, _06662_, _06662_, _06662_, _06662_, _06662_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17299" *) wt0_sd_data[1007:1000];
  assign _04129_ = { _06663_, _06663_, _06663_, _06663_, _06663_, _06663_, _06663_, _06663_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17309" *) wt0_sd_data[1015:1008];
  assign _04130_ = { _06664_, _06664_, _06664_, _06664_, _06664_, _06664_, _06664_, _06664_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17319" *) wt0_sd_data[1023:1016];
  assign _04131_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17352" *) wt1_actv_pvld_w;
  assign _04132_ = _04131_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17362" *) cfg_is_fp16_d1[75];
  assign _04133_ = { _06665_, _06665_, _06665_, _06665_, _06665_, _06665_, _06665_, _06665_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17373" *) wt1_sd_data[7:0];
  assign _04134_ = { _06666_, _06666_, _06666_, _06666_, _06666_, _06666_, _06666_, _06666_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17383" *) wt1_sd_data[15:8];
  assign _04135_ = { _06667_, _06667_, _06667_, _06667_, _06667_, _06667_, _06667_, _06667_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17393" *) wt1_sd_data[23:16];
  assign _04136_ = { _06668_, _06668_, _06668_, _06668_, _06668_, _06668_, _06668_, _06668_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17403" *) wt1_sd_data[31:24];
  assign _04137_ = { _06669_, _06669_, _06669_, _06669_, _06669_, _06669_, _06669_, _06669_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17413" *) wt1_sd_data[39:32];
  assign _04138_ = { _06670_, _06670_, _06670_, _06670_, _06670_, _06670_, _06670_, _06670_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17423" *) wt1_sd_data[47:40];
  assign _04139_ = { _06671_, _06671_, _06671_, _06671_, _06671_, _06671_, _06671_, _06671_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17433" *) wt1_sd_data[55:48];
  assign _04140_ = { _06672_, _06672_, _06672_, _06672_, _06672_, _06672_, _06672_, _06672_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17443" *) wt1_sd_data[63:56];
  assign _04141_ = { _06673_, _06673_, _06673_, _06673_, _06673_, _06673_, _06673_, _06673_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17453" *) wt1_sd_data[71:64];
  assign _04142_ = { _06674_, _06674_, _06674_, _06674_, _06674_, _06674_, _06674_, _06674_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17463" *) wt1_sd_data[79:72];
  assign _04143_ = { _06675_, _06675_, _06675_, _06675_, _06675_, _06675_, _06675_, _06675_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17473" *) wt1_sd_data[87:80];
  assign _04144_ = { _06676_, _06676_, _06676_, _06676_, _06676_, _06676_, _06676_, _06676_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17483" *) wt1_sd_data[95:88];
  assign _04145_ = { _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17493" *) wt1_sd_data[103:96];
  assign _04146_ = { _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17503" *) wt1_sd_data[111:104];
  assign _04147_ = { _06679_, _06679_, _06679_, _06679_, _06679_, _06679_, _06679_, _06679_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17513" *) wt1_sd_data[119:112];
  assign _04148_ = { _06680_, _06680_, _06680_, _06680_, _06680_, _06680_, _06680_, _06680_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17523" *) wt1_sd_data[127:120];
  assign _04149_ = { _06681_, _06681_, _06681_, _06681_, _06681_, _06681_, _06681_, _06681_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17533" *) wt1_sd_data[135:128];
  assign _04150_ = { _06682_, _06682_, _06682_, _06682_, _06682_, _06682_, _06682_, _06682_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17543" *) wt1_sd_data[143:136];
  assign _04151_ = { _06683_, _06683_, _06683_, _06683_, _06683_, _06683_, _06683_, _06683_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17553" *) wt1_sd_data[151:144];
  assign _04152_ = { _06684_, _06684_, _06684_, _06684_, _06684_, _06684_, _06684_, _06684_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17563" *) wt1_sd_data[159:152];
  assign _04153_ = { _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17573" *) wt1_sd_data[167:160];
  assign _04154_ = { _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17583" *) wt1_sd_data[175:168];
  assign _04155_ = { _06687_, _06687_, _06687_, _06687_, _06687_, _06687_, _06687_, _06687_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17593" *) wt1_sd_data[183:176];
  assign _04156_ = { _06688_, _06688_, _06688_, _06688_, _06688_, _06688_, _06688_, _06688_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17603" *) wt1_sd_data[191:184];
  assign _04157_ = { _06689_, _06689_, _06689_, _06689_, _06689_, _06689_, _06689_, _06689_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17613" *) wt1_sd_data[199:192];
  assign _04158_ = { _06690_, _06690_, _06690_, _06690_, _06690_, _06690_, _06690_, _06690_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17623" *) wt1_sd_data[207:200];
  assign _04159_ = { _06691_, _06691_, _06691_, _06691_, _06691_, _06691_, _06691_, _06691_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17633" *) wt1_sd_data[215:208];
  assign _04160_ = { _06692_, _06692_, _06692_, _06692_, _06692_, _06692_, _06692_, _06692_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17643" *) wt1_sd_data[223:216];
  assign _04161_ = { _06693_, _06693_, _06693_, _06693_, _06693_, _06693_, _06693_, _06693_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17653" *) wt1_sd_data[231:224];
  assign _04162_ = { _06694_, _06694_, _06694_, _06694_, _06694_, _06694_, _06694_, _06694_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17663" *) wt1_sd_data[239:232];
  assign _04163_ = { _06695_, _06695_, _06695_, _06695_, _06695_, _06695_, _06695_, _06695_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17673" *) wt1_sd_data[247:240];
  assign _04164_ = { _06696_, _06696_, _06696_, _06696_, _06696_, _06696_, _06696_, _06696_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17683" *) wt1_sd_data[255:248];
  assign _04165_ = { _06697_, _06697_, _06697_, _06697_, _06697_, _06697_, _06697_, _06697_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17693" *) wt1_sd_data[263:256];
  assign _04166_ = { _06698_, _06698_, _06698_, _06698_, _06698_, _06698_, _06698_, _06698_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17703" *) wt1_sd_data[271:264];
  assign _04167_ = { _06699_, _06699_, _06699_, _06699_, _06699_, _06699_, _06699_, _06699_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17713" *) wt1_sd_data[279:272];
  assign _04168_ = { _06700_, _06700_, _06700_, _06700_, _06700_, _06700_, _06700_, _06700_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17723" *) wt1_sd_data[287:280];
  assign _04169_ = { _06701_, _06701_, _06701_, _06701_, _06701_, _06701_, _06701_, _06701_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17733" *) wt1_sd_data[295:288];
  assign _04170_ = { _06702_, _06702_, _06702_, _06702_, _06702_, _06702_, _06702_, _06702_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17743" *) wt1_sd_data[303:296];
  assign _04171_ = { _06703_, _06703_, _06703_, _06703_, _06703_, _06703_, _06703_, _06703_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17753" *) wt1_sd_data[311:304];
  assign _04172_ = { _06704_, _06704_, _06704_, _06704_, _06704_, _06704_, _06704_, _06704_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17763" *) wt1_sd_data[319:312];
  assign _04173_ = { _06705_, _06705_, _06705_, _06705_, _06705_, _06705_, _06705_, _06705_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17773" *) wt1_sd_data[327:320];
  assign _04174_ = { _06706_, _06706_, _06706_, _06706_, _06706_, _06706_, _06706_, _06706_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17783" *) wt1_sd_data[335:328];
  assign _04175_ = { _06707_, _06707_, _06707_, _06707_, _06707_, _06707_, _06707_, _06707_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17793" *) wt1_sd_data[343:336];
  assign _04176_ = { _06708_, _06708_, _06708_, _06708_, _06708_, _06708_, _06708_, _06708_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17803" *) wt1_sd_data[351:344];
  assign _04177_ = { _06709_, _06709_, _06709_, _06709_, _06709_, _06709_, _06709_, _06709_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17813" *) wt1_sd_data[359:352];
  assign _04178_ = { _06710_, _06710_, _06710_, _06710_, _06710_, _06710_, _06710_, _06710_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17823" *) wt1_sd_data[367:360];
  assign _04179_ = { _06711_, _06711_, _06711_, _06711_, _06711_, _06711_, _06711_, _06711_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17833" *) wt1_sd_data[375:368];
  assign _04180_ = { _06712_, _06712_, _06712_, _06712_, _06712_, _06712_, _06712_, _06712_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17843" *) wt1_sd_data[383:376];
  assign _04181_ = { _06713_, _06713_, _06713_, _06713_, _06713_, _06713_, _06713_, _06713_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17853" *) wt1_sd_data[391:384];
  assign _04182_ = { _06714_, _06714_, _06714_, _06714_, _06714_, _06714_, _06714_, _06714_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17863" *) wt1_sd_data[399:392];
  assign _04183_ = { _06715_, _06715_, _06715_, _06715_, _06715_, _06715_, _06715_, _06715_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17873" *) wt1_sd_data[407:400];
  assign _04184_ = { _06716_, _06716_, _06716_, _06716_, _06716_, _06716_, _06716_, _06716_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17883" *) wt1_sd_data[415:408];
  assign _04185_ = { _06717_, _06717_, _06717_, _06717_, _06717_, _06717_, _06717_, _06717_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17893" *) wt1_sd_data[423:416];
  assign _04186_ = { _06718_, _06718_, _06718_, _06718_, _06718_, _06718_, _06718_, _06718_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17903" *) wt1_sd_data[431:424];
  assign _04187_ = { _06719_, _06719_, _06719_, _06719_, _06719_, _06719_, _06719_, _06719_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17913" *) wt1_sd_data[439:432];
  assign _04188_ = { _06720_, _06720_, _06720_, _06720_, _06720_, _06720_, _06720_, _06720_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17923" *) wt1_sd_data[447:440];
  assign _04189_ = { _06721_, _06721_, _06721_, _06721_, _06721_, _06721_, _06721_, _06721_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17933" *) wt1_sd_data[455:448];
  assign _04190_ = { _06722_, _06722_, _06722_, _06722_, _06722_, _06722_, _06722_, _06722_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17943" *) wt1_sd_data[463:456];
  assign _04191_ = { _06723_, _06723_, _06723_, _06723_, _06723_, _06723_, _06723_, _06723_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17953" *) wt1_sd_data[471:464];
  assign _04192_ = { _06724_, _06724_, _06724_, _06724_, _06724_, _06724_, _06724_, _06724_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17963" *) wt1_sd_data[479:472];
  assign _04193_ = { _06725_, _06725_, _06725_, _06725_, _06725_, _06725_, _06725_, _06725_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17973" *) wt1_sd_data[487:480];
  assign _04194_ = { _06726_, _06726_, _06726_, _06726_, _06726_, _06726_, _06726_, _06726_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17983" *) wt1_sd_data[495:488];
  assign _04195_ = { _06727_, _06727_, _06727_, _06727_, _06727_, _06727_, _06727_, _06727_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17993" *) wt1_sd_data[503:496];
  assign _04196_ = { _06728_, _06728_, _06728_, _06728_, _06728_, _06728_, _06728_, _06728_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18003" *) wt1_sd_data[511:504];
  assign _04197_ = { _06729_, _06729_, _06729_, _06729_, _06729_, _06729_, _06729_, _06729_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18013" *) wt1_sd_data[519:512];
  assign _04198_ = { _06730_, _06730_, _06730_, _06730_, _06730_, _06730_, _06730_, _06730_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18023" *) wt1_sd_data[527:520];
  assign _04199_ = { _06731_, _06731_, _06731_, _06731_, _06731_, _06731_, _06731_, _06731_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18033" *) wt1_sd_data[535:528];
  assign _04200_ = { _06732_, _06732_, _06732_, _06732_, _06732_, _06732_, _06732_, _06732_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18043" *) wt1_sd_data[543:536];
  assign _04201_ = { _06733_, _06733_, _06733_, _06733_, _06733_, _06733_, _06733_, _06733_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18053" *) wt1_sd_data[551:544];
  assign _04202_ = { _06734_, _06734_, _06734_, _06734_, _06734_, _06734_, _06734_, _06734_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18063" *) wt1_sd_data[559:552];
  assign _04203_ = { _06735_, _06735_, _06735_, _06735_, _06735_, _06735_, _06735_, _06735_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18073" *) wt1_sd_data[567:560];
  assign _04204_ = { _06736_, _06736_, _06736_, _06736_, _06736_, _06736_, _06736_, _06736_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18083" *) wt1_sd_data[575:568];
  assign _04205_ = { _06737_, _06737_, _06737_, _06737_, _06737_, _06737_, _06737_, _06737_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18093" *) wt1_sd_data[583:576];
  assign _04206_ = { _06738_, _06738_, _06738_, _06738_, _06738_, _06738_, _06738_, _06738_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18103" *) wt1_sd_data[591:584];
  assign _04207_ = { _06739_, _06739_, _06739_, _06739_, _06739_, _06739_, _06739_, _06739_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18113" *) wt1_sd_data[599:592];
  assign _04208_ = { _06740_, _06740_, _06740_, _06740_, _06740_, _06740_, _06740_, _06740_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18123" *) wt1_sd_data[607:600];
  assign _04209_ = { _06741_, _06741_, _06741_, _06741_, _06741_, _06741_, _06741_, _06741_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18133" *) wt1_sd_data[615:608];
  assign _04210_ = { _06742_, _06742_, _06742_, _06742_, _06742_, _06742_, _06742_, _06742_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18143" *) wt1_sd_data[623:616];
  assign _04211_ = { _06743_, _06743_, _06743_, _06743_, _06743_, _06743_, _06743_, _06743_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18153" *) wt1_sd_data[631:624];
  assign _04212_ = { _06744_, _06744_, _06744_, _06744_, _06744_, _06744_, _06744_, _06744_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18163" *) wt1_sd_data[639:632];
  assign _04213_ = { _06745_, _06745_, _06745_, _06745_, _06745_, _06745_, _06745_, _06745_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18173" *) wt1_sd_data[647:640];
  assign _04214_ = { _06746_, _06746_, _06746_, _06746_, _06746_, _06746_, _06746_, _06746_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18183" *) wt1_sd_data[655:648];
  assign _04215_ = { _06747_, _06747_, _06747_, _06747_, _06747_, _06747_, _06747_, _06747_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18193" *) wt1_sd_data[663:656];
  assign _04216_ = { _06748_, _06748_, _06748_, _06748_, _06748_, _06748_, _06748_, _06748_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18203" *) wt1_sd_data[671:664];
  assign _04217_ = { _06749_, _06749_, _06749_, _06749_, _06749_, _06749_, _06749_, _06749_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18213" *) wt1_sd_data[679:672];
  assign _04218_ = { _06750_, _06750_, _06750_, _06750_, _06750_, _06750_, _06750_, _06750_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18223" *) wt1_sd_data[687:680];
  assign _04219_ = { _06751_, _06751_, _06751_, _06751_, _06751_, _06751_, _06751_, _06751_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18233" *) wt1_sd_data[695:688];
  assign _04220_ = { _06752_, _06752_, _06752_, _06752_, _06752_, _06752_, _06752_, _06752_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18243" *) wt1_sd_data[703:696];
  assign _04221_ = { _06753_, _06753_, _06753_, _06753_, _06753_, _06753_, _06753_, _06753_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18253" *) wt1_sd_data[711:704];
  assign _04222_ = { _06754_, _06754_, _06754_, _06754_, _06754_, _06754_, _06754_, _06754_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18263" *) wt1_sd_data[719:712];
  assign _04223_ = { _06755_, _06755_, _06755_, _06755_, _06755_, _06755_, _06755_, _06755_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18273" *) wt1_sd_data[727:720];
  assign _04224_ = { _06756_, _06756_, _06756_, _06756_, _06756_, _06756_, _06756_, _06756_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18283" *) wt1_sd_data[735:728];
  assign _04225_ = { _06757_, _06757_, _06757_, _06757_, _06757_, _06757_, _06757_, _06757_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18293" *) wt1_sd_data[743:736];
  assign _04226_ = { _06758_, _06758_, _06758_, _06758_, _06758_, _06758_, _06758_, _06758_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18303" *) wt1_sd_data[751:744];
  assign _04227_ = { _06759_, _06759_, _06759_, _06759_, _06759_, _06759_, _06759_, _06759_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18313" *) wt1_sd_data[759:752];
  assign _04228_ = { _06760_, _06760_, _06760_, _06760_, _06760_, _06760_, _06760_, _06760_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18323" *) wt1_sd_data[767:760];
  assign _04229_ = { _06761_, _06761_, _06761_, _06761_, _06761_, _06761_, _06761_, _06761_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18333" *) wt1_sd_data[775:768];
  assign _04230_ = { _06762_, _06762_, _06762_, _06762_, _06762_, _06762_, _06762_, _06762_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18343" *) wt1_sd_data[783:776];
  assign _04231_ = { _06763_, _06763_, _06763_, _06763_, _06763_, _06763_, _06763_, _06763_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18353" *) wt1_sd_data[791:784];
  assign _04232_ = { _06764_, _06764_, _06764_, _06764_, _06764_, _06764_, _06764_, _06764_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18363" *) wt1_sd_data[799:792];
  assign _04233_ = { _06765_, _06765_, _06765_, _06765_, _06765_, _06765_, _06765_, _06765_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18373" *) wt1_sd_data[807:800];
  assign _04234_ = { _06766_, _06766_, _06766_, _06766_, _06766_, _06766_, _06766_, _06766_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18383" *) wt1_sd_data[815:808];
  assign _04235_ = { _06767_, _06767_, _06767_, _06767_, _06767_, _06767_, _06767_, _06767_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18393" *) wt1_sd_data[823:816];
  assign _04236_ = { _06768_, _06768_, _06768_, _06768_, _06768_, _06768_, _06768_, _06768_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18403" *) wt1_sd_data[831:824];
  assign _04237_ = { _06769_, _06769_, _06769_, _06769_, _06769_, _06769_, _06769_, _06769_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18413" *) wt1_sd_data[839:832];
  assign _04238_ = { _06770_, _06770_, _06770_, _06770_, _06770_, _06770_, _06770_, _06770_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18423" *) wt1_sd_data[847:840];
  assign _04239_ = { _06771_, _06771_, _06771_, _06771_, _06771_, _06771_, _06771_, _06771_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18433" *) wt1_sd_data[855:848];
  assign _04240_ = { _06772_, _06772_, _06772_, _06772_, _06772_, _06772_, _06772_, _06772_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18443" *) wt1_sd_data[863:856];
  assign _04241_ = { _06773_, _06773_, _06773_, _06773_, _06773_, _06773_, _06773_, _06773_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18453" *) wt1_sd_data[871:864];
  assign _04242_ = { _06774_, _06774_, _06774_, _06774_, _06774_, _06774_, _06774_, _06774_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18463" *) wt1_sd_data[879:872];
  assign _04243_ = { _06775_, _06775_, _06775_, _06775_, _06775_, _06775_, _06775_, _06775_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18473" *) wt1_sd_data[887:880];
  assign _04244_ = { _06776_, _06776_, _06776_, _06776_, _06776_, _06776_, _06776_, _06776_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18483" *) wt1_sd_data[895:888];
  assign _04245_ = { _06777_, _06777_, _06777_, _06777_, _06777_, _06777_, _06777_, _06777_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18493" *) wt1_sd_data[903:896];
  assign _04246_ = { _06778_, _06778_, _06778_, _06778_, _06778_, _06778_, _06778_, _06778_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18503" *) wt1_sd_data[911:904];
  assign _04247_ = { _06779_, _06779_, _06779_, _06779_, _06779_, _06779_, _06779_, _06779_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18513" *) wt1_sd_data[919:912];
  assign _04248_ = { _06780_, _06780_, _06780_, _06780_, _06780_, _06780_, _06780_, _06780_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18523" *) wt1_sd_data[927:920];
  assign _04249_ = { _06781_, _06781_, _06781_, _06781_, _06781_, _06781_, _06781_, _06781_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18533" *) wt1_sd_data[935:928];
  assign _04250_ = { _06782_, _06782_, _06782_, _06782_, _06782_, _06782_, _06782_, _06782_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18543" *) wt1_sd_data[943:936];
  assign _04251_ = { _06783_, _06783_, _06783_, _06783_, _06783_, _06783_, _06783_, _06783_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18553" *) wt1_sd_data[951:944];
  assign _04252_ = { _06784_, _06784_, _06784_, _06784_, _06784_, _06784_, _06784_, _06784_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18563" *) wt1_sd_data[959:952];
  assign _04253_ = { _06785_, _06785_, _06785_, _06785_, _06785_, _06785_, _06785_, _06785_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18573" *) wt1_sd_data[967:960];
  assign _04254_ = { _06786_, _06786_, _06786_, _06786_, _06786_, _06786_, _06786_, _06786_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18583" *) wt1_sd_data[975:968];
  assign _04255_ = { _06787_, _06787_, _06787_, _06787_, _06787_, _06787_, _06787_, _06787_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18593" *) wt1_sd_data[983:976];
  assign _04256_ = { _06788_, _06788_, _06788_, _06788_, _06788_, _06788_, _06788_, _06788_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18603" *) wt1_sd_data[991:984];
  assign _04257_ = { _06789_, _06789_, _06789_, _06789_, _06789_, _06789_, _06789_, _06789_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18613" *) wt1_sd_data[999:992];
  assign _04258_ = { _06790_, _06790_, _06790_, _06790_, _06790_, _06790_, _06790_, _06790_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18623" *) wt1_sd_data[1007:1000];
  assign _04259_ = { _06791_, _06791_, _06791_, _06791_, _06791_, _06791_, _06791_, _06791_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18633" *) wt1_sd_data[1015:1008];
  assign _04260_ = { _06792_, _06792_, _06792_, _06792_, _06792_, _06792_, _06792_, _06792_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18643" *) wt1_sd_data[1023:1016];
  assign _04261_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18676" *) wt2_actv_pvld_w;
  assign _04262_ = _04261_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18686" *) cfg_is_fp16_d1[76];
  assign _04263_ = { _06793_, _06793_, _06793_, _06793_, _06793_, _06793_, _06793_, _06793_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18697" *) wt2_sd_data[7:0];
  assign _04264_ = { _06794_, _06794_, _06794_, _06794_, _06794_, _06794_, _06794_, _06794_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18707" *) wt2_sd_data[15:8];
  assign _04265_ = { _06795_, _06795_, _06795_, _06795_, _06795_, _06795_, _06795_, _06795_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18717" *) wt2_sd_data[23:16];
  assign _04266_ = { _06796_, _06796_, _06796_, _06796_, _06796_, _06796_, _06796_, _06796_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18727" *) wt2_sd_data[31:24];
  assign _04267_ = { _06797_, _06797_, _06797_, _06797_, _06797_, _06797_, _06797_, _06797_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18737" *) wt2_sd_data[39:32];
  assign _04268_ = { _06798_, _06798_, _06798_, _06798_, _06798_, _06798_, _06798_, _06798_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18747" *) wt2_sd_data[47:40];
  assign _04269_ = { _06799_, _06799_, _06799_, _06799_, _06799_, _06799_, _06799_, _06799_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18757" *) wt2_sd_data[55:48];
  assign _04270_ = { _06800_, _06800_, _06800_, _06800_, _06800_, _06800_, _06800_, _06800_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18767" *) wt2_sd_data[63:56];
  assign _04271_ = { _06801_, _06801_, _06801_, _06801_, _06801_, _06801_, _06801_, _06801_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18777" *) wt2_sd_data[71:64];
  assign _04272_ = { _06802_, _06802_, _06802_, _06802_, _06802_, _06802_, _06802_, _06802_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18787" *) wt2_sd_data[79:72];
  assign _04273_ = { _06803_, _06803_, _06803_, _06803_, _06803_, _06803_, _06803_, _06803_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18797" *) wt2_sd_data[87:80];
  assign _04274_ = { _06804_, _06804_, _06804_, _06804_, _06804_, _06804_, _06804_, _06804_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18807" *) wt2_sd_data[95:88];
  assign _04275_ = { _06805_, _06805_, _06805_, _06805_, _06805_, _06805_, _06805_, _06805_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18817" *) wt2_sd_data[103:96];
  assign _04276_ = { _06806_, _06806_, _06806_, _06806_, _06806_, _06806_, _06806_, _06806_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18827" *) wt2_sd_data[111:104];
  assign _04277_ = { _06807_, _06807_, _06807_, _06807_, _06807_, _06807_, _06807_, _06807_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18837" *) wt2_sd_data[119:112];
  assign _04278_ = { _06808_, _06808_, _06808_, _06808_, _06808_, _06808_, _06808_, _06808_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18847" *) wt2_sd_data[127:120];
  assign _04279_ = { _06809_, _06809_, _06809_, _06809_, _06809_, _06809_, _06809_, _06809_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18857" *) wt2_sd_data[135:128];
  assign _04280_ = { _06810_, _06810_, _06810_, _06810_, _06810_, _06810_, _06810_, _06810_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18867" *) wt2_sd_data[143:136];
  assign _04281_ = { _06811_, _06811_, _06811_, _06811_, _06811_, _06811_, _06811_, _06811_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18877" *) wt2_sd_data[151:144];
  assign _04282_ = { _06812_, _06812_, _06812_, _06812_, _06812_, _06812_, _06812_, _06812_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18887" *) wt2_sd_data[159:152];
  assign _04283_ = { _06813_, _06813_, _06813_, _06813_, _06813_, _06813_, _06813_, _06813_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18897" *) wt2_sd_data[167:160];
  assign _04284_ = { _06814_, _06814_, _06814_, _06814_, _06814_, _06814_, _06814_, _06814_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18907" *) wt2_sd_data[175:168];
  assign _04285_ = { _06815_, _06815_, _06815_, _06815_, _06815_, _06815_, _06815_, _06815_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18917" *) wt2_sd_data[183:176];
  assign _04286_ = { _06816_, _06816_, _06816_, _06816_, _06816_, _06816_, _06816_, _06816_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18927" *) wt2_sd_data[191:184];
  assign _04287_ = { _06817_, _06817_, _06817_, _06817_, _06817_, _06817_, _06817_, _06817_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18937" *) wt2_sd_data[199:192];
  assign _04288_ = { _06818_, _06818_, _06818_, _06818_, _06818_, _06818_, _06818_, _06818_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18947" *) wt2_sd_data[207:200];
  assign _04289_ = { _06819_, _06819_, _06819_, _06819_, _06819_, _06819_, _06819_, _06819_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18957" *) wt2_sd_data[215:208];
  assign _04290_ = { _06820_, _06820_, _06820_, _06820_, _06820_, _06820_, _06820_, _06820_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18967" *) wt2_sd_data[223:216];
  assign _04291_ = { _06821_, _06821_, _06821_, _06821_, _06821_, _06821_, _06821_, _06821_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18977" *) wt2_sd_data[231:224];
  assign _04292_ = { _06822_, _06822_, _06822_, _06822_, _06822_, _06822_, _06822_, _06822_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18987" *) wt2_sd_data[239:232];
  assign _04293_ = { _06823_, _06823_, _06823_, _06823_, _06823_, _06823_, _06823_, _06823_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18997" *) wt2_sd_data[247:240];
  assign _04294_ = { _06824_, _06824_, _06824_, _06824_, _06824_, _06824_, _06824_, _06824_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19007" *) wt2_sd_data[255:248];
  assign _04295_ = { _06825_, _06825_, _06825_, _06825_, _06825_, _06825_, _06825_, _06825_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19017" *) wt2_sd_data[263:256];
  assign _04296_ = { _06826_, _06826_, _06826_, _06826_, _06826_, _06826_, _06826_, _06826_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19027" *) wt2_sd_data[271:264];
  assign _04297_ = { _06827_, _06827_, _06827_, _06827_, _06827_, _06827_, _06827_, _06827_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19037" *) wt2_sd_data[279:272];
  assign _04298_ = { _06828_, _06828_, _06828_, _06828_, _06828_, _06828_, _06828_, _06828_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19047" *) wt2_sd_data[287:280];
  assign _04299_ = { _06829_, _06829_, _06829_, _06829_, _06829_, _06829_, _06829_, _06829_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19057" *) wt2_sd_data[295:288];
  assign _04300_ = { _06830_, _06830_, _06830_, _06830_, _06830_, _06830_, _06830_, _06830_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19067" *) wt2_sd_data[303:296];
  assign _04301_ = { _06831_, _06831_, _06831_, _06831_, _06831_, _06831_, _06831_, _06831_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19077" *) wt2_sd_data[311:304];
  assign _04302_ = { _06832_, _06832_, _06832_, _06832_, _06832_, _06832_, _06832_, _06832_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19087" *) wt2_sd_data[319:312];
  assign _04303_ = { _06833_, _06833_, _06833_, _06833_, _06833_, _06833_, _06833_, _06833_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19097" *) wt2_sd_data[327:320];
  assign _04304_ = { _06834_, _06834_, _06834_, _06834_, _06834_, _06834_, _06834_, _06834_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19107" *) wt2_sd_data[335:328];
  assign _04305_ = { _06835_, _06835_, _06835_, _06835_, _06835_, _06835_, _06835_, _06835_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19117" *) wt2_sd_data[343:336];
  assign _04306_ = { _06836_, _06836_, _06836_, _06836_, _06836_, _06836_, _06836_, _06836_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19127" *) wt2_sd_data[351:344];
  assign _04307_ = { _06837_, _06837_, _06837_, _06837_, _06837_, _06837_, _06837_, _06837_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19137" *) wt2_sd_data[359:352];
  assign _04308_ = { _06838_, _06838_, _06838_, _06838_, _06838_, _06838_, _06838_, _06838_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19147" *) wt2_sd_data[367:360];
  assign _04309_ = { _06839_, _06839_, _06839_, _06839_, _06839_, _06839_, _06839_, _06839_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19157" *) wt2_sd_data[375:368];
  assign _04310_ = { _06840_, _06840_, _06840_, _06840_, _06840_, _06840_, _06840_, _06840_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19167" *) wt2_sd_data[383:376];
  assign _04311_ = { _06841_, _06841_, _06841_, _06841_, _06841_, _06841_, _06841_, _06841_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19177" *) wt2_sd_data[391:384];
  assign _04312_ = { _06842_, _06842_, _06842_, _06842_, _06842_, _06842_, _06842_, _06842_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19187" *) wt2_sd_data[399:392];
  assign _04313_ = { _06843_, _06843_, _06843_, _06843_, _06843_, _06843_, _06843_, _06843_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19197" *) wt2_sd_data[407:400];
  assign _04314_ = { _06844_, _06844_, _06844_, _06844_, _06844_, _06844_, _06844_, _06844_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19207" *) wt2_sd_data[415:408];
  assign _04315_ = { _06845_, _06845_, _06845_, _06845_, _06845_, _06845_, _06845_, _06845_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19217" *) wt2_sd_data[423:416];
  assign _04316_ = { _06846_, _06846_, _06846_, _06846_, _06846_, _06846_, _06846_, _06846_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19227" *) wt2_sd_data[431:424];
  assign _04317_ = { _06847_, _06847_, _06847_, _06847_, _06847_, _06847_, _06847_, _06847_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19237" *) wt2_sd_data[439:432];
  assign _04318_ = { _06848_, _06848_, _06848_, _06848_, _06848_, _06848_, _06848_, _06848_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19247" *) wt2_sd_data[447:440];
  assign _04319_ = { _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19257" *) wt2_sd_data[455:448];
  assign _04320_ = { _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19267" *) wt2_sd_data[463:456];
  assign _04321_ = { _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19277" *) wt2_sd_data[471:464];
  assign _04322_ = { _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19287" *) wt2_sd_data[479:472];
  assign _04323_ = { _06853_, _06853_, _06853_, _06853_, _06853_, _06853_, _06853_, _06853_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19297" *) wt2_sd_data[487:480];
  assign _04324_ = { _06854_, _06854_, _06854_, _06854_, _06854_, _06854_, _06854_, _06854_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19307" *) wt2_sd_data[495:488];
  assign _04325_ = { _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19317" *) wt2_sd_data[503:496];
  assign _04326_ = { _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19327" *) wt2_sd_data[511:504];
  assign _04327_ = { _06857_, _06857_, _06857_, _06857_, _06857_, _06857_, _06857_, _06857_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19337" *) wt2_sd_data[519:512];
  assign _04328_ = { _06858_, _06858_, _06858_, _06858_, _06858_, _06858_, _06858_, _06858_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19347" *) wt2_sd_data[527:520];
  assign _04329_ = { _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19357" *) wt2_sd_data[535:528];
  assign _04330_ = { _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19367" *) wt2_sd_data[543:536];
  assign _04331_ = { _06861_, _06861_, _06861_, _06861_, _06861_, _06861_, _06861_, _06861_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19377" *) wt2_sd_data[551:544];
  assign _04332_ = { _06862_, _06862_, _06862_, _06862_, _06862_, _06862_, _06862_, _06862_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19387" *) wt2_sd_data[559:552];
  assign _04333_ = { _06863_, _06863_, _06863_, _06863_, _06863_, _06863_, _06863_, _06863_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19397" *) wt2_sd_data[567:560];
  assign _04334_ = { _06864_, _06864_, _06864_, _06864_, _06864_, _06864_, _06864_, _06864_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19407" *) wt2_sd_data[575:568];
  assign _04335_ = { _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19417" *) wt2_sd_data[583:576];
  assign _04336_ = { _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19427" *) wt2_sd_data[591:584];
  assign _04337_ = { _06867_, _06867_, _06867_, _06867_, _06867_, _06867_, _06867_, _06867_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19437" *) wt2_sd_data[599:592];
  assign _04338_ = { _06868_, _06868_, _06868_, _06868_, _06868_, _06868_, _06868_, _06868_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19447" *) wt2_sd_data[607:600];
  assign _04339_ = { _06869_, _06869_, _06869_, _06869_, _06869_, _06869_, _06869_, _06869_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19457" *) wt2_sd_data[615:608];
  assign _04340_ = { _06870_, _06870_, _06870_, _06870_, _06870_, _06870_, _06870_, _06870_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19467" *) wt2_sd_data[623:616];
  assign _04341_ = { _06871_, _06871_, _06871_, _06871_, _06871_, _06871_, _06871_, _06871_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19477" *) wt2_sd_data[631:624];
  assign _04342_ = { _06872_, _06872_, _06872_, _06872_, _06872_, _06872_, _06872_, _06872_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19487" *) wt2_sd_data[639:632];
  assign _04343_ = { _06873_, _06873_, _06873_, _06873_, _06873_, _06873_, _06873_, _06873_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19497" *) wt2_sd_data[647:640];
  assign _04344_ = { _06874_, _06874_, _06874_, _06874_, _06874_, _06874_, _06874_, _06874_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19507" *) wt2_sd_data[655:648];
  assign _04345_ = { _06875_, _06875_, _06875_, _06875_, _06875_, _06875_, _06875_, _06875_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19517" *) wt2_sd_data[663:656];
  assign _04346_ = { _06876_, _06876_, _06876_, _06876_, _06876_, _06876_, _06876_, _06876_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19527" *) wt2_sd_data[671:664];
  assign _04347_ = { _06877_, _06877_, _06877_, _06877_, _06877_, _06877_, _06877_, _06877_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19537" *) wt2_sd_data[679:672];
  assign _04348_ = { _06878_, _06878_, _06878_, _06878_, _06878_, _06878_, _06878_, _06878_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19547" *) wt2_sd_data[687:680];
  assign _04349_ = { _06879_, _06879_, _06879_, _06879_, _06879_, _06879_, _06879_, _06879_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19557" *) wt2_sd_data[695:688];
  assign _04350_ = { _06880_, _06880_, _06880_, _06880_, _06880_, _06880_, _06880_, _06880_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19567" *) wt2_sd_data[703:696];
  assign _04351_ = { _06881_, _06881_, _06881_, _06881_, _06881_, _06881_, _06881_, _06881_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19577" *) wt2_sd_data[711:704];
  assign _04352_ = { _06882_, _06882_, _06882_, _06882_, _06882_, _06882_, _06882_, _06882_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19587" *) wt2_sd_data[719:712];
  assign _04353_ = { _06883_, _06883_, _06883_, _06883_, _06883_, _06883_, _06883_, _06883_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19597" *) wt2_sd_data[727:720];
  assign _04354_ = { _06884_, _06884_, _06884_, _06884_, _06884_, _06884_, _06884_, _06884_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19607" *) wt2_sd_data[735:728];
  assign _04355_ = { _06885_, _06885_, _06885_, _06885_, _06885_, _06885_, _06885_, _06885_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19617" *) wt2_sd_data[743:736];
  assign _04356_ = { _06886_, _06886_, _06886_, _06886_, _06886_, _06886_, _06886_, _06886_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19627" *) wt2_sd_data[751:744];
  assign _04357_ = { _06887_, _06887_, _06887_, _06887_, _06887_, _06887_, _06887_, _06887_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19637" *) wt2_sd_data[759:752];
  assign _04358_ = { _06888_, _06888_, _06888_, _06888_, _06888_, _06888_, _06888_, _06888_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19647" *) wt2_sd_data[767:760];
  assign _04359_ = { _06889_, _06889_, _06889_, _06889_, _06889_, _06889_, _06889_, _06889_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19657" *) wt2_sd_data[775:768];
  assign _04360_ = { _06890_, _06890_, _06890_, _06890_, _06890_, _06890_, _06890_, _06890_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19667" *) wt2_sd_data[783:776];
  assign _04361_ = { _06891_, _06891_, _06891_, _06891_, _06891_, _06891_, _06891_, _06891_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19677" *) wt2_sd_data[791:784];
  assign _04362_ = { _06892_, _06892_, _06892_, _06892_, _06892_, _06892_, _06892_, _06892_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19687" *) wt2_sd_data[799:792];
  assign _04363_ = { _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19697" *) wt2_sd_data[807:800];
  assign _04364_ = { _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19707" *) wt2_sd_data[815:808];
  assign _04365_ = { _06895_, _06895_, _06895_, _06895_, _06895_, _06895_, _06895_, _06895_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19717" *) wt2_sd_data[823:816];
  assign _04366_ = { _06896_, _06896_, _06896_, _06896_, _06896_, _06896_, _06896_, _06896_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19727" *) wt2_sd_data[831:824];
  assign _04367_ = { _06897_, _06897_, _06897_, _06897_, _06897_, _06897_, _06897_, _06897_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19737" *) wt2_sd_data[839:832];
  assign _04368_ = { _06898_, _06898_, _06898_, _06898_, _06898_, _06898_, _06898_, _06898_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19747" *) wt2_sd_data[847:840];
  assign _04369_ = { _06899_, _06899_, _06899_, _06899_, _06899_, _06899_, _06899_, _06899_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19757" *) wt2_sd_data[855:848];
  assign _04370_ = { _06900_, _06900_, _06900_, _06900_, _06900_, _06900_, _06900_, _06900_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19767" *) wt2_sd_data[863:856];
  assign _04371_ = { _06901_, _06901_, _06901_, _06901_, _06901_, _06901_, _06901_, _06901_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19777" *) wt2_sd_data[871:864];
  assign _04372_ = { _06902_, _06902_, _06902_, _06902_, _06902_, _06902_, _06902_, _06902_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19787" *) wt2_sd_data[879:872];
  assign _04373_ = { _06903_, _06903_, _06903_, _06903_, _06903_, _06903_, _06903_, _06903_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19797" *) wt2_sd_data[887:880];
  assign _04374_ = { _06904_, _06904_, _06904_, _06904_, _06904_, _06904_, _06904_, _06904_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19807" *) wt2_sd_data[895:888];
  assign _04375_ = { _06905_, _06905_, _06905_, _06905_, _06905_, _06905_, _06905_, _06905_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19817" *) wt2_sd_data[903:896];
  assign _04376_ = { _06906_, _06906_, _06906_, _06906_, _06906_, _06906_, _06906_, _06906_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19827" *) wt2_sd_data[911:904];
  assign _04377_ = { _06907_, _06907_, _06907_, _06907_, _06907_, _06907_, _06907_, _06907_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19837" *) wt2_sd_data[919:912];
  assign _04378_ = { _06908_, _06908_, _06908_, _06908_, _06908_, _06908_, _06908_, _06908_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19847" *) wt2_sd_data[927:920];
  assign _04379_ = { _06909_, _06909_, _06909_, _06909_, _06909_, _06909_, _06909_, _06909_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19857" *) wt2_sd_data[935:928];
  assign _04380_ = { _06910_, _06910_, _06910_, _06910_, _06910_, _06910_, _06910_, _06910_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19867" *) wt2_sd_data[943:936];
  assign _04381_ = { _06911_, _06911_, _06911_, _06911_, _06911_, _06911_, _06911_, _06911_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19877" *) wt2_sd_data[951:944];
  assign _04382_ = { _06912_, _06912_, _06912_, _06912_, _06912_, _06912_, _06912_, _06912_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19887" *) wt2_sd_data[959:952];
  assign _04383_ = { _06913_, _06913_, _06913_, _06913_, _06913_, _06913_, _06913_, _06913_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19897" *) wt2_sd_data[967:960];
  assign _04384_ = { _06914_, _06914_, _06914_, _06914_, _06914_, _06914_, _06914_, _06914_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19907" *) wt2_sd_data[975:968];
  assign _04385_ = { _06915_, _06915_, _06915_, _06915_, _06915_, _06915_, _06915_, _06915_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19917" *) wt2_sd_data[983:976];
  assign _04386_ = { _06916_, _06916_, _06916_, _06916_, _06916_, _06916_, _06916_, _06916_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19927" *) wt2_sd_data[991:984];
  assign _04387_ = { _06917_, _06917_, _06917_, _06917_, _06917_, _06917_, _06917_, _06917_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19937" *) wt2_sd_data[999:992];
  assign _04388_ = { _06918_, _06918_, _06918_, _06918_, _06918_, _06918_, _06918_, _06918_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19947" *) wt2_sd_data[1007:1000];
  assign _04389_ = { _06919_, _06919_, _06919_, _06919_, _06919_, _06919_, _06919_, _06919_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19957" *) wt2_sd_data[1015:1008];
  assign _04390_ = { _06920_, _06920_, _06920_, _06920_, _06920_, _06920_, _06920_, _06920_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19967" *) wt2_sd_data[1023:1016];
  assign _04391_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20000" *) wt3_actv_pvld_w;
  assign _04392_ = _04391_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20010" *) cfg_is_fp16_d1[77];
  assign _04393_ = { _06921_, _06921_, _06921_, _06921_, _06921_, _06921_, _06921_, _06921_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20021" *) wt3_sd_data[7:0];
  assign _04394_ = { _06922_, _06922_, _06922_, _06922_, _06922_, _06922_, _06922_, _06922_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20031" *) wt3_sd_data[15:8];
  assign _04395_ = { _06923_, _06923_, _06923_, _06923_, _06923_, _06923_, _06923_, _06923_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20041" *) wt3_sd_data[23:16];
  assign _04396_ = { _06924_, _06924_, _06924_, _06924_, _06924_, _06924_, _06924_, _06924_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20051" *) wt3_sd_data[31:24];
  assign _04397_ = { _06925_, _06925_, _06925_, _06925_, _06925_, _06925_, _06925_, _06925_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20061" *) wt3_sd_data[39:32];
  assign _04398_ = { _06926_, _06926_, _06926_, _06926_, _06926_, _06926_, _06926_, _06926_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20071" *) wt3_sd_data[47:40];
  assign _04399_ = { _06927_, _06927_, _06927_, _06927_, _06927_, _06927_, _06927_, _06927_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20081" *) wt3_sd_data[55:48];
  assign _04400_ = { _06928_, _06928_, _06928_, _06928_, _06928_, _06928_, _06928_, _06928_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20091" *) wt3_sd_data[63:56];
  assign _04401_ = { _06929_, _06929_, _06929_, _06929_, _06929_, _06929_, _06929_, _06929_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20101" *) wt3_sd_data[71:64];
  assign _04402_ = { _06930_, _06930_, _06930_, _06930_, _06930_, _06930_, _06930_, _06930_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20111" *) wt3_sd_data[79:72];
  assign _04403_ = { _06931_, _06931_, _06931_, _06931_, _06931_, _06931_, _06931_, _06931_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20121" *) wt3_sd_data[87:80];
  assign _04404_ = { _06932_, _06932_, _06932_, _06932_, _06932_, _06932_, _06932_, _06932_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20131" *) wt3_sd_data[95:88];
  assign _04405_ = { _06933_, _06933_, _06933_, _06933_, _06933_, _06933_, _06933_, _06933_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20141" *) wt3_sd_data[103:96];
  assign _04406_ = { _06934_, _06934_, _06934_, _06934_, _06934_, _06934_, _06934_, _06934_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20151" *) wt3_sd_data[111:104];
  assign _04407_ = { _06935_, _06935_, _06935_, _06935_, _06935_, _06935_, _06935_, _06935_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20161" *) wt3_sd_data[119:112];
  assign _04408_ = { _06936_, _06936_, _06936_, _06936_, _06936_, _06936_, _06936_, _06936_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20171" *) wt3_sd_data[127:120];
  assign _04409_ = { _06937_, _06937_, _06937_, _06937_, _06937_, _06937_, _06937_, _06937_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20181" *) wt3_sd_data[135:128];
  assign _04410_ = { _06938_, _06938_, _06938_, _06938_, _06938_, _06938_, _06938_, _06938_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20191" *) wt3_sd_data[143:136];
  assign _04411_ = { _06939_, _06939_, _06939_, _06939_, _06939_, _06939_, _06939_, _06939_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20201" *) wt3_sd_data[151:144];
  assign _04412_ = { _06940_, _06940_, _06940_, _06940_, _06940_, _06940_, _06940_, _06940_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20211" *) wt3_sd_data[159:152];
  assign _04413_ = { _06941_, _06941_, _06941_, _06941_, _06941_, _06941_, _06941_, _06941_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20221" *) wt3_sd_data[167:160];
  assign _04414_ = { _06942_, _06942_, _06942_, _06942_, _06942_, _06942_, _06942_, _06942_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20231" *) wt3_sd_data[175:168];
  assign _04415_ = { _06943_, _06943_, _06943_, _06943_, _06943_, _06943_, _06943_, _06943_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20241" *) wt3_sd_data[183:176];
  assign _04416_ = { _06944_, _06944_, _06944_, _06944_, _06944_, _06944_, _06944_, _06944_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20251" *) wt3_sd_data[191:184];
  assign _04417_ = { _06945_, _06945_, _06945_, _06945_, _06945_, _06945_, _06945_, _06945_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20261" *) wt3_sd_data[199:192];
  assign _04418_ = { _06946_, _06946_, _06946_, _06946_, _06946_, _06946_, _06946_, _06946_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20271" *) wt3_sd_data[207:200];
  assign _04419_ = { _06947_, _06947_, _06947_, _06947_, _06947_, _06947_, _06947_, _06947_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20281" *) wt3_sd_data[215:208];
  assign _04420_ = { _06948_, _06948_, _06948_, _06948_, _06948_, _06948_, _06948_, _06948_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20291" *) wt3_sd_data[223:216];
  assign _04421_ = { _06949_, _06949_, _06949_, _06949_, _06949_, _06949_, _06949_, _06949_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20301" *) wt3_sd_data[231:224];
  assign _04422_ = { _06950_, _06950_, _06950_, _06950_, _06950_, _06950_, _06950_, _06950_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20311" *) wt3_sd_data[239:232];
  assign _04423_ = { _06951_, _06951_, _06951_, _06951_, _06951_, _06951_, _06951_, _06951_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20321" *) wt3_sd_data[247:240];
  assign _04424_ = { _06952_, _06952_, _06952_, _06952_, _06952_, _06952_, _06952_, _06952_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20331" *) wt3_sd_data[255:248];
  assign _04425_ = { _06953_, _06953_, _06953_, _06953_, _06953_, _06953_, _06953_, _06953_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20341" *) wt3_sd_data[263:256];
  assign _04426_ = { _06954_, _06954_, _06954_, _06954_, _06954_, _06954_, _06954_, _06954_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20351" *) wt3_sd_data[271:264];
  assign _04427_ = { _06955_, _06955_, _06955_, _06955_, _06955_, _06955_, _06955_, _06955_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20361" *) wt3_sd_data[279:272];
  assign _04428_ = { _06956_, _06956_, _06956_, _06956_, _06956_, _06956_, _06956_, _06956_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20371" *) wt3_sd_data[287:280];
  assign _04429_ = { _06957_, _06957_, _06957_, _06957_, _06957_, _06957_, _06957_, _06957_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20381" *) wt3_sd_data[295:288];
  assign _04430_ = { _06958_, _06958_, _06958_, _06958_, _06958_, _06958_, _06958_, _06958_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20391" *) wt3_sd_data[303:296];
  assign _04431_ = { _06959_, _06959_, _06959_, _06959_, _06959_, _06959_, _06959_, _06959_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20401" *) wt3_sd_data[311:304];
  assign _04432_ = { _06960_, _06960_, _06960_, _06960_, _06960_, _06960_, _06960_, _06960_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20411" *) wt3_sd_data[319:312];
  assign _04433_ = { _06961_, _06961_, _06961_, _06961_, _06961_, _06961_, _06961_, _06961_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20421" *) wt3_sd_data[327:320];
  assign _04434_ = { _06962_, _06962_, _06962_, _06962_, _06962_, _06962_, _06962_, _06962_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20431" *) wt3_sd_data[335:328];
  assign _04435_ = { _06963_, _06963_, _06963_, _06963_, _06963_, _06963_, _06963_, _06963_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20441" *) wt3_sd_data[343:336];
  assign _04436_ = { _06964_, _06964_, _06964_, _06964_, _06964_, _06964_, _06964_, _06964_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20451" *) wt3_sd_data[351:344];
  assign _04437_ = { _06965_, _06965_, _06965_, _06965_, _06965_, _06965_, _06965_, _06965_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20461" *) wt3_sd_data[359:352];
  assign _04438_ = { _06966_, _06966_, _06966_, _06966_, _06966_, _06966_, _06966_, _06966_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20471" *) wt3_sd_data[367:360];
  assign _04439_ = { _06967_, _06967_, _06967_, _06967_, _06967_, _06967_, _06967_, _06967_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20481" *) wt3_sd_data[375:368];
  assign _04440_ = { _06968_, _06968_, _06968_, _06968_, _06968_, _06968_, _06968_, _06968_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20491" *) wt3_sd_data[383:376];
  assign _04441_ = { _06969_, _06969_, _06969_, _06969_, _06969_, _06969_, _06969_, _06969_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20501" *) wt3_sd_data[391:384];
  assign _04442_ = { _06970_, _06970_, _06970_, _06970_, _06970_, _06970_, _06970_, _06970_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20511" *) wt3_sd_data[399:392];
  assign _04443_ = { _06971_, _06971_, _06971_, _06971_, _06971_, _06971_, _06971_, _06971_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20521" *) wt3_sd_data[407:400];
  assign _04444_ = { _06972_, _06972_, _06972_, _06972_, _06972_, _06972_, _06972_, _06972_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20531" *) wt3_sd_data[415:408];
  assign _04445_ = { _06973_, _06973_, _06973_, _06973_, _06973_, _06973_, _06973_, _06973_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20541" *) wt3_sd_data[423:416];
  assign _04446_ = { _06974_, _06974_, _06974_, _06974_, _06974_, _06974_, _06974_, _06974_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20551" *) wt3_sd_data[431:424];
  assign _04447_ = { _06975_, _06975_, _06975_, _06975_, _06975_, _06975_, _06975_, _06975_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20561" *) wt3_sd_data[439:432];
  assign _04448_ = { _06976_, _06976_, _06976_, _06976_, _06976_, _06976_, _06976_, _06976_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20571" *) wt3_sd_data[447:440];
  assign _04449_ = { _06977_, _06977_, _06977_, _06977_, _06977_, _06977_, _06977_, _06977_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20581" *) wt3_sd_data[455:448];
  assign _04450_ = { _06978_, _06978_, _06978_, _06978_, _06978_, _06978_, _06978_, _06978_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20591" *) wt3_sd_data[463:456];
  assign _04451_ = { _06979_, _06979_, _06979_, _06979_, _06979_, _06979_, _06979_, _06979_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20601" *) wt3_sd_data[471:464];
  assign _04452_ = { _06980_, _06980_, _06980_, _06980_, _06980_, _06980_, _06980_, _06980_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20611" *) wt3_sd_data[479:472];
  assign _04453_ = { _06981_, _06981_, _06981_, _06981_, _06981_, _06981_, _06981_, _06981_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20621" *) wt3_sd_data[487:480];
  assign _04454_ = { _06982_, _06982_, _06982_, _06982_, _06982_, _06982_, _06982_, _06982_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20631" *) wt3_sd_data[495:488];
  assign _04455_ = { _06983_, _06983_, _06983_, _06983_, _06983_, _06983_, _06983_, _06983_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20641" *) wt3_sd_data[503:496];
  assign _04456_ = { _06984_, _06984_, _06984_, _06984_, _06984_, _06984_, _06984_, _06984_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20651" *) wt3_sd_data[511:504];
  assign _04457_ = { _06985_, _06985_, _06985_, _06985_, _06985_, _06985_, _06985_, _06985_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20661" *) wt3_sd_data[519:512];
  assign _04458_ = { _06986_, _06986_, _06986_, _06986_, _06986_, _06986_, _06986_, _06986_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20671" *) wt3_sd_data[527:520];
  assign _04459_ = { _06987_, _06987_, _06987_, _06987_, _06987_, _06987_, _06987_, _06987_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20681" *) wt3_sd_data[535:528];
  assign _04460_ = { _06988_, _06988_, _06988_, _06988_, _06988_, _06988_, _06988_, _06988_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20691" *) wt3_sd_data[543:536];
  assign _04461_ = { _06989_, _06989_, _06989_, _06989_, _06989_, _06989_, _06989_, _06989_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20701" *) wt3_sd_data[551:544];
  assign _04462_ = { _06990_, _06990_, _06990_, _06990_, _06990_, _06990_, _06990_, _06990_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20711" *) wt3_sd_data[559:552];
  assign _04463_ = { _06991_, _06991_, _06991_, _06991_, _06991_, _06991_, _06991_, _06991_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20721" *) wt3_sd_data[567:560];
  assign _04464_ = { _06992_, _06992_, _06992_, _06992_, _06992_, _06992_, _06992_, _06992_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20731" *) wt3_sd_data[575:568];
  assign _04465_ = { _06993_, _06993_, _06993_, _06993_, _06993_, _06993_, _06993_, _06993_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20741" *) wt3_sd_data[583:576];
  assign _04466_ = { _06994_, _06994_, _06994_, _06994_, _06994_, _06994_, _06994_, _06994_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20751" *) wt3_sd_data[591:584];
  assign _04467_ = { _06995_, _06995_, _06995_, _06995_, _06995_, _06995_, _06995_, _06995_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20761" *) wt3_sd_data[599:592];
  assign _04468_ = { _06996_, _06996_, _06996_, _06996_, _06996_, _06996_, _06996_, _06996_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20771" *) wt3_sd_data[607:600];
  assign _04469_ = { _06997_, _06997_, _06997_, _06997_, _06997_, _06997_, _06997_, _06997_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20781" *) wt3_sd_data[615:608];
  assign _04470_ = { _06998_, _06998_, _06998_, _06998_, _06998_, _06998_, _06998_, _06998_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20791" *) wt3_sd_data[623:616];
  assign _04471_ = { _06999_, _06999_, _06999_, _06999_, _06999_, _06999_, _06999_, _06999_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20801" *) wt3_sd_data[631:624];
  assign _04472_ = { _07000_, _07000_, _07000_, _07000_, _07000_, _07000_, _07000_, _07000_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20811" *) wt3_sd_data[639:632];
  assign _04473_ = { _07001_, _07001_, _07001_, _07001_, _07001_, _07001_, _07001_, _07001_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20821" *) wt3_sd_data[647:640];
  assign _04474_ = { _07002_, _07002_, _07002_, _07002_, _07002_, _07002_, _07002_, _07002_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20831" *) wt3_sd_data[655:648];
  assign _04475_ = { _07003_, _07003_, _07003_, _07003_, _07003_, _07003_, _07003_, _07003_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20841" *) wt3_sd_data[663:656];
  assign _04476_ = { _07004_, _07004_, _07004_, _07004_, _07004_, _07004_, _07004_, _07004_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20851" *) wt3_sd_data[671:664];
  assign _04477_ = { _07005_, _07005_, _07005_, _07005_, _07005_, _07005_, _07005_, _07005_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20861" *) wt3_sd_data[679:672];
  assign _04478_ = { _07006_, _07006_, _07006_, _07006_, _07006_, _07006_, _07006_, _07006_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20871" *) wt3_sd_data[687:680];
  assign _04479_ = { _07007_, _07007_, _07007_, _07007_, _07007_, _07007_, _07007_, _07007_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20881" *) wt3_sd_data[695:688];
  assign _04480_ = { _07008_, _07008_, _07008_, _07008_, _07008_, _07008_, _07008_, _07008_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20891" *) wt3_sd_data[703:696];
  assign _04481_ = { _07009_, _07009_, _07009_, _07009_, _07009_, _07009_, _07009_, _07009_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20901" *) wt3_sd_data[711:704];
  assign _04482_ = { _07010_, _07010_, _07010_, _07010_, _07010_, _07010_, _07010_, _07010_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20911" *) wt3_sd_data[719:712];
  assign _04483_ = { _07011_, _07011_, _07011_, _07011_, _07011_, _07011_, _07011_, _07011_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20921" *) wt3_sd_data[727:720];
  assign _04484_ = { _07012_, _07012_, _07012_, _07012_, _07012_, _07012_, _07012_, _07012_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20931" *) wt3_sd_data[735:728];
  assign _04485_ = { _07013_, _07013_, _07013_, _07013_, _07013_, _07013_, _07013_, _07013_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20941" *) wt3_sd_data[743:736];
  assign _04486_ = { _07014_, _07014_, _07014_, _07014_, _07014_, _07014_, _07014_, _07014_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20951" *) wt3_sd_data[751:744];
  assign _04487_ = { _07015_, _07015_, _07015_, _07015_, _07015_, _07015_, _07015_, _07015_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20961" *) wt3_sd_data[759:752];
  assign _04488_ = { _07016_, _07016_, _07016_, _07016_, _07016_, _07016_, _07016_, _07016_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20971" *) wt3_sd_data[767:760];
  assign _04489_ = { _07017_, _07017_, _07017_, _07017_, _07017_, _07017_, _07017_, _07017_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20981" *) wt3_sd_data[775:768];
  assign _04490_ = { _07018_, _07018_, _07018_, _07018_, _07018_, _07018_, _07018_, _07018_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20991" *) wt3_sd_data[783:776];
  assign _04491_ = { _07019_, _07019_, _07019_, _07019_, _07019_, _07019_, _07019_, _07019_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21001" *) wt3_sd_data[791:784];
  assign _04492_ = { _07020_, _07020_, _07020_, _07020_, _07020_, _07020_, _07020_, _07020_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21011" *) wt3_sd_data[799:792];
  assign _04493_ = { _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21021" *) wt3_sd_data[807:800];
  assign _04494_ = { _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21031" *) wt3_sd_data[815:808];
  assign _04495_ = { _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21041" *) wt3_sd_data[823:816];
  assign _04496_ = { _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21051" *) wt3_sd_data[831:824];
  assign _04497_ = { _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21061" *) wt3_sd_data[839:832];
  assign _04498_ = { _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21071" *) wt3_sd_data[847:840];
  assign _04499_ = { _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21081" *) wt3_sd_data[855:848];
  assign _04500_ = { _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21091" *) wt3_sd_data[863:856];
  assign _04501_ = { _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21101" *) wt3_sd_data[871:864];
  assign _04502_ = { _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21111" *) wt3_sd_data[879:872];
  assign _04503_ = { _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21121" *) wt3_sd_data[887:880];
  assign _04504_ = { _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21131" *) wt3_sd_data[895:888];
  assign _04505_ = { _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21141" *) wt3_sd_data[903:896];
  assign _04506_ = { _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21151" *) wt3_sd_data[911:904];
  assign _04507_ = { _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21161" *) wt3_sd_data[919:912];
  assign _04508_ = { _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21171" *) wt3_sd_data[927:920];
  assign _04509_ = { _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21181" *) wt3_sd_data[935:928];
  assign _04510_ = { _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21191" *) wt3_sd_data[943:936];
  assign _04511_ = { _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21201" *) wt3_sd_data[951:944];
  assign _04512_ = { _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21211" *) wt3_sd_data[959:952];
  assign _04513_ = { _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21221" *) wt3_sd_data[967:960];
  assign _04514_ = { _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21231" *) wt3_sd_data[975:968];
  assign _04515_ = { _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21241" *) wt3_sd_data[983:976];
  assign _04516_ = { _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21251" *) wt3_sd_data[991:984];
  assign _04517_ = { _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21261" *) wt3_sd_data[999:992];
  assign _04518_ = { _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21271" *) wt3_sd_data[1007:1000];
  assign _04519_ = { _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21281" *) wt3_sd_data[1015:1008];
  assign _04520_ = { _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21291" *) wt3_sd_data[1023:1016];
  assign _04521_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21324" *) wt4_actv_pvld_w;
  assign _04522_ = _04521_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21334" *) cfg_is_fp16_d1[78];
  assign _04523_ = { _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21345" *) wt4_sd_data[7:0];
  assign _04524_ = { _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21355" *) wt4_sd_data[15:8];
  assign _04525_ = { _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21365" *) wt4_sd_data[23:16];
  assign _04526_ = { _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21375" *) wt4_sd_data[31:24];
  assign _04527_ = { _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21385" *) wt4_sd_data[39:32];
  assign _04528_ = { _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21395" *) wt4_sd_data[47:40];
  assign _04529_ = { _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21405" *) wt4_sd_data[55:48];
  assign _04530_ = { _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21415" *) wt4_sd_data[63:56];
  assign _04531_ = { _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21425" *) wt4_sd_data[71:64];
  assign _04532_ = { _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21435" *) wt4_sd_data[79:72];
  assign _04533_ = { _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21445" *) wt4_sd_data[87:80];
  assign _04534_ = { _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21455" *) wt4_sd_data[95:88];
  assign _04535_ = { _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21465" *) wt4_sd_data[103:96];
  assign _04536_ = { _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21475" *) wt4_sd_data[111:104];
  assign _04537_ = { _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21485" *) wt4_sd_data[119:112];
  assign _04538_ = { _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21495" *) wt4_sd_data[127:120];
  assign _04539_ = { _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21505" *) wt4_sd_data[135:128];
  assign _04540_ = { _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21515" *) wt4_sd_data[143:136];
  assign _04541_ = { _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21525" *) wt4_sd_data[151:144];
  assign _04542_ = { _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21535" *) wt4_sd_data[159:152];
  assign _04543_ = { _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21545" *) wt4_sd_data[167:160];
  assign _04544_ = { _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21555" *) wt4_sd_data[175:168];
  assign _04545_ = { _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21565" *) wt4_sd_data[183:176];
  assign _04546_ = { _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21575" *) wt4_sd_data[191:184];
  assign _04547_ = { _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21585" *) wt4_sd_data[199:192];
  assign _04548_ = { _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21595" *) wt4_sd_data[207:200];
  assign _04549_ = { _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21605" *) wt4_sd_data[215:208];
  assign _04550_ = { _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21615" *) wt4_sd_data[223:216];
  assign _04551_ = { _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21625" *) wt4_sd_data[231:224];
  assign _04552_ = { _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21635" *) wt4_sd_data[239:232];
  assign _04553_ = { _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21645" *) wt4_sd_data[247:240];
  assign _04554_ = { _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21655" *) wt4_sd_data[255:248];
  assign _04555_ = { _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21665" *) wt4_sd_data[263:256];
  assign _04556_ = { _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21675" *) wt4_sd_data[271:264];
  assign _04557_ = { _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21685" *) wt4_sd_data[279:272];
  assign _04558_ = { _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21695" *) wt4_sd_data[287:280];
  assign _04559_ = { _07085_, _07085_, _07085_, _07085_, _07085_, _07085_, _07085_, _07085_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21705" *) wt4_sd_data[295:288];
  assign _04560_ = { _07086_, _07086_, _07086_, _07086_, _07086_, _07086_, _07086_, _07086_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21715" *) wt4_sd_data[303:296];
  assign in_wt_data_int16_63 = { cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2172" *) { in_wt_data127, in_wt_data126 };
  assign _04561_ = { _07087_, _07087_, _07087_, _07087_, _07087_, _07087_, _07087_, _07087_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21725" *) wt4_sd_data[311:304];
  assign in_wt_data_int16_62 = { cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2173" *) { in_wt_data125, in_wt_data124 };
  assign _04562_ = { _07088_, _07088_, _07088_, _07088_, _07088_, _07088_, _07088_, _07088_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21735" *) wt4_sd_data[319:312];
  assign in_wt_data_int16_61 = { cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2174" *) { in_wt_data123, in_wt_data122 };
  assign _04563_ = { _07089_, _07089_, _07089_, _07089_, _07089_, _07089_, _07089_, _07089_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21745" *) wt4_sd_data[327:320];
  assign in_wt_data_int16_60 = { cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2175" *) { in_wt_data121, in_wt_data120 };
  assign _04564_ = { _07090_, _07090_, _07090_, _07090_, _07090_, _07090_, _07090_, _07090_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21755" *) wt4_sd_data[335:328];
  assign in_wt_data_int16_59 = { cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2176" *) { in_wt_data119, in_wt_data118 };
  assign _04565_ = { _07091_, _07091_, _07091_, _07091_, _07091_, _07091_, _07091_, _07091_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21765" *) wt4_sd_data[343:336];
  assign in_wt_data_int16_58 = { cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2177" *) { in_wt_data117, in_wt_data116 };
  assign _04566_ = { _07092_, _07092_, _07092_, _07092_, _07092_, _07092_, _07092_, _07092_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21775" *) wt4_sd_data[351:344];
  assign in_wt_data_int16_57 = { cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2178" *) { in_wt_data115, in_wt_data114 };
  assign _04567_ = { _07093_, _07093_, _07093_, _07093_, _07093_, _07093_, _07093_, _07093_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21785" *) wt4_sd_data[359:352];
  assign in_wt_data_int16_56 = { cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2179" *) { in_wt_data113, in_wt_data112 };
  assign _04568_ = { _07094_, _07094_, _07094_, _07094_, _07094_, _07094_, _07094_, _07094_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21795" *) wt4_sd_data[367:360];
  assign in_wt_data_int16_55 = { cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2180" *) { in_wt_data111, in_wt_data110 };
  assign _04569_ = { _07095_, _07095_, _07095_, _07095_, _07095_, _07095_, _07095_, _07095_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21805" *) wt4_sd_data[375:368];
  assign in_wt_data_int16_54 = { cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2181" *) { in_wt_data109, in_wt_data108 };
  assign _04570_ = { _07096_, _07096_, _07096_, _07096_, _07096_, _07096_, _07096_, _07096_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21815" *) wt4_sd_data[383:376];
  assign in_wt_data_int16_53 = { cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2182" *) { in_wt_data107, in_wt_data106 };
  assign _04571_ = { _07097_, _07097_, _07097_, _07097_, _07097_, _07097_, _07097_, _07097_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21825" *) wt4_sd_data[391:384];
  assign in_wt_data_int16_52 = { cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2183" *) { in_wt_data105, in_wt_data104 };
  assign _04572_ = { _07098_, _07098_, _07098_, _07098_, _07098_, _07098_, _07098_, _07098_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21835" *) wt4_sd_data[399:392];
  assign in_wt_data_int16_51 = { cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2184" *) { in_wt_data103, in_wt_data102 };
  assign _04573_ = { _07099_, _07099_, _07099_, _07099_, _07099_, _07099_, _07099_, _07099_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21845" *) wt4_sd_data[407:400];
  assign in_wt_data_int16_50 = { cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2185" *) { in_wt_data101, in_wt_data100 };
  assign _04574_ = { _07100_, _07100_, _07100_, _07100_, _07100_, _07100_, _07100_, _07100_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21855" *) wt4_sd_data[415:408];
  assign in_wt_data_int16_49 = { cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2186" *) { in_wt_data99, in_wt_data98 };
  assign _04575_ = { _07101_, _07101_, _07101_, _07101_, _07101_, _07101_, _07101_, _07101_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21865" *) wt4_sd_data[423:416];
  assign in_wt_data_int16_48 = { cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2187" *) { in_wt_data97, in_wt_data96 };
  assign _04576_ = { _07102_, _07102_, _07102_, _07102_, _07102_, _07102_, _07102_, _07102_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21875" *) wt4_sd_data[431:424];
  assign in_wt_data_int16_47 = { cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2188" *) { in_wt_data95, in_wt_data94 };
  assign _04577_ = { _07103_, _07103_, _07103_, _07103_, _07103_, _07103_, _07103_, _07103_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21885" *) wt4_sd_data[439:432];
  assign in_wt_data_int16_46 = { cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2189" *) { in_wt_data93, in_wt_data92 };
  assign _04578_ = { _07104_, _07104_, _07104_, _07104_, _07104_, _07104_, _07104_, _07104_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21895" *) wt4_sd_data[447:440];
  assign in_wt_data_int16_45 = { cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2190" *) { in_wt_data91, in_wt_data90 };
  assign _04579_ = { _07105_, _07105_, _07105_, _07105_, _07105_, _07105_, _07105_, _07105_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21905" *) wt4_sd_data[455:448];
  assign in_wt_data_int16_44 = { cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2191" *) { in_wt_data89, in_wt_data88 };
  assign _04580_ = { _07106_, _07106_, _07106_, _07106_, _07106_, _07106_, _07106_, _07106_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21915" *) wt4_sd_data[463:456];
  assign in_wt_data_int16_43 = { cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2192" *) { in_wt_data87, in_wt_data86 };
  assign _04581_ = { _07107_, _07107_, _07107_, _07107_, _07107_, _07107_, _07107_, _07107_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21925" *) wt4_sd_data[471:464];
  assign in_wt_data_int16_42 = { cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2193" *) { in_wt_data85, in_wt_data84 };
  assign _04582_ = { _07108_, _07108_, _07108_, _07108_, _07108_, _07108_, _07108_, _07108_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21935" *) wt4_sd_data[479:472];
  assign in_wt_data_int16_41 = { cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2194" *) { in_wt_data83, in_wt_data82 };
  assign _04583_ = { _07109_, _07109_, _07109_, _07109_, _07109_, _07109_, _07109_, _07109_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21945" *) wt4_sd_data[487:480];
  assign in_wt_data_int16_40 = { cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2195" *) { in_wt_data81, in_wt_data80 };
  assign _04584_ = { _07110_, _07110_, _07110_, _07110_, _07110_, _07110_, _07110_, _07110_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21955" *) wt4_sd_data[495:488];
  assign in_wt_data_int16_39 = { cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2196" *) { in_wt_data79, in_wt_data78 };
  assign _04585_ = { _07111_, _07111_, _07111_, _07111_, _07111_, _07111_, _07111_, _07111_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21965" *) wt4_sd_data[503:496];
  assign in_wt_data_int16_38 = { cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2197" *) { in_wt_data77, in_wt_data76 };
  assign _04586_ = { _07112_, _07112_, _07112_, _07112_, _07112_, _07112_, _07112_, _07112_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21975" *) wt4_sd_data[511:504];
  assign in_wt_data_int16_37 = { cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2198" *) { in_wt_data75, in_wt_data74 };
  assign _04587_ = { _07113_, _07113_, _07113_, _07113_, _07113_, _07113_, _07113_, _07113_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21985" *) wt4_sd_data[519:512];
  assign in_wt_data_int16_36 = { cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2199" *) { in_wt_data73, in_wt_data72 };
  assign _04588_ = { _07114_, _07114_, _07114_, _07114_, _07114_, _07114_, _07114_, _07114_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21995" *) wt4_sd_data[527:520];
  assign in_wt_data_int16_35 = { cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2200" *) { in_wt_data71, in_wt_data70 };
  assign _04589_ = { _07115_, _07115_, _07115_, _07115_, _07115_, _07115_, _07115_, _07115_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22005" *) wt4_sd_data[535:528];
  assign in_wt_data_int16_34 = { cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2201" *) { in_wt_data69, in_wt_data68 };
  assign _04590_ = { _07116_, _07116_, _07116_, _07116_, _07116_, _07116_, _07116_, _07116_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22015" *) wt4_sd_data[543:536];
  assign in_wt_data_int16_33 = { cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2202" *) { in_wt_data67, in_wt_data66 };
  assign _04591_ = { _07117_, _07117_, _07117_, _07117_, _07117_, _07117_, _07117_, _07117_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22025" *) wt4_sd_data[551:544];
  assign in_wt_data_int16_32 = { cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2203" *) { in_wt_data65, in_wt_data64 };
  assign _04592_ = { _07118_, _07118_, _07118_, _07118_, _07118_, _07118_, _07118_, _07118_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22035" *) wt4_sd_data[559:552];
  assign in_wt_data_int16_31 = { cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2204" *) { in_wt_data63, in_wt_data62 };
  assign _04593_ = { _07119_, _07119_, _07119_, _07119_, _07119_, _07119_, _07119_, _07119_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22045" *) wt4_sd_data[567:560];
  assign in_wt_data_int16_30 = { cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2205" *) { in_wt_data61, in_wt_data60 };
  assign _04594_ = { _07120_, _07120_, _07120_, _07120_, _07120_, _07120_, _07120_, _07120_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22055" *) wt4_sd_data[575:568];
  assign in_wt_data_int16_29 = { cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2206" *) { in_wt_data59, in_wt_data58 };
  assign _04595_ = { _07121_, _07121_, _07121_, _07121_, _07121_, _07121_, _07121_, _07121_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22065" *) wt4_sd_data[583:576];
  assign in_wt_data_int16_28 = { cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2207" *) { in_wt_data57, in_wt_data56 };
  assign _04596_ = { _07122_, _07122_, _07122_, _07122_, _07122_, _07122_, _07122_, _07122_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22075" *) wt4_sd_data[591:584];
  assign in_wt_data_int16_27 = { cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2208" *) { in_wt_data55, in_wt_data54 };
  assign _04597_ = { _07123_, _07123_, _07123_, _07123_, _07123_, _07123_, _07123_, _07123_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22085" *) wt4_sd_data[599:592];
  assign in_wt_data_int16_26 = { cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2209" *) { in_wt_data53, in_wt_data52 };
  assign _04598_ = { _07124_, _07124_, _07124_, _07124_, _07124_, _07124_, _07124_, _07124_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22095" *) wt4_sd_data[607:600];
  assign in_wt_data_int16_25 = { cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2210" *) { in_wt_data51, in_wt_data50 };
  assign _04599_ = { _07125_, _07125_, _07125_, _07125_, _07125_, _07125_, _07125_, _07125_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22105" *) wt4_sd_data[615:608];
  assign in_wt_data_int16_24 = { cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2211" *) { in_wt_data49, in_wt_data48 };
  assign _04600_ = { _07126_, _07126_, _07126_, _07126_, _07126_, _07126_, _07126_, _07126_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22115" *) wt4_sd_data[623:616];
  assign in_wt_data_int16_23 = { cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2212" *) { in_wt_data47, in_wt_data46 };
  assign _04601_ = { _07127_, _07127_, _07127_, _07127_, _07127_, _07127_, _07127_, _07127_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22125" *) wt4_sd_data[631:624];
  assign in_wt_data_int16_22 = { cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2213" *) { in_wt_data45, in_wt_data44 };
  assign _04602_ = { _07128_, _07128_, _07128_, _07128_, _07128_, _07128_, _07128_, _07128_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22135" *) wt4_sd_data[639:632];
  assign in_wt_data_int16_21 = { cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2214" *) { in_wt_data43, in_wt_data42 };
  assign _04603_ = { _07129_, _07129_, _07129_, _07129_, _07129_, _07129_, _07129_, _07129_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22145" *) wt4_sd_data[647:640];
  assign in_wt_data_int16_20 = { cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2215" *) { in_wt_data41, in_wt_data40 };
  assign _04604_ = { _07130_, _07130_, _07130_, _07130_, _07130_, _07130_, _07130_, _07130_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22155" *) wt4_sd_data[655:648];
  assign in_wt_data_int16_19 = { cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2216" *) { in_wt_data39, in_wt_data38 };
  assign _04605_ = { _07131_, _07131_, _07131_, _07131_, _07131_, _07131_, _07131_, _07131_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22165" *) wt4_sd_data[663:656];
  assign in_wt_data_int16_18 = { cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2217" *) { in_wt_data37, in_wt_data36 };
  assign _04606_ = { _07132_, _07132_, _07132_, _07132_, _07132_, _07132_, _07132_, _07132_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22175" *) wt4_sd_data[671:664];
  assign in_wt_data_int16_17 = { cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2218" *) { in_wt_data35, in_wt_data34 };
  assign _04607_ = { _07133_, _07133_, _07133_, _07133_, _07133_, _07133_, _07133_, _07133_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22185" *) wt4_sd_data[679:672];
  assign in_wt_data_int16_16 = { cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2219" *) { in_wt_data33, in_wt_data32 };
  assign _04608_ = { _07134_, _07134_, _07134_, _07134_, _07134_, _07134_, _07134_, _07134_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22195" *) wt4_sd_data[687:680];
  assign in_wt_data_int16_15 = { cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2220" *) { in_wt_data31, in_wt_data30 };
  assign _04609_ = { _07135_, _07135_, _07135_, _07135_, _07135_, _07135_, _07135_, _07135_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22205" *) wt4_sd_data[695:688];
  assign in_wt_data_int16_14 = { cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2221" *) { in_wt_data29, in_wt_data28 };
  assign _04610_ = { _07136_, _07136_, _07136_, _07136_, _07136_, _07136_, _07136_, _07136_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22215" *) wt4_sd_data[703:696];
  assign in_wt_data_int16_13 = { cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2222" *) { in_wt_data27, in_wt_data26 };
  assign _04611_ = { _07137_, _07137_, _07137_, _07137_, _07137_, _07137_, _07137_, _07137_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22225" *) wt4_sd_data[711:704];
  assign in_wt_data_int16_12 = { cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2223" *) { in_wt_data25, in_wt_data24 };
  assign _04612_ = { _07138_, _07138_, _07138_, _07138_, _07138_, _07138_, _07138_, _07138_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22235" *) wt4_sd_data[719:712];
  assign in_wt_data_int16_11 = { cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2224" *) { in_wt_data23, in_wt_data22 };
  assign _04613_ = { _07139_, _07139_, _07139_, _07139_, _07139_, _07139_, _07139_, _07139_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22245" *) wt4_sd_data[727:720];
  assign in_wt_data_int16_10 = { cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2225" *) { in_wt_data21, in_wt_data20 };
  assign _04614_ = { _07140_, _07140_, _07140_, _07140_, _07140_, _07140_, _07140_, _07140_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22255" *) wt4_sd_data[735:728];
  assign in_wt_data_int16_9 = { cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2226" *) { in_wt_data19, in_wt_data18 };
  assign _04615_ = { _07141_, _07141_, _07141_, _07141_, _07141_, _07141_, _07141_, _07141_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22265" *) wt4_sd_data[743:736];
  assign in_wt_data_int16_8 = { cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2227" *) { in_wt_data17, in_wt_data16 };
  assign _04616_ = { _07142_, _07142_, _07142_, _07142_, _07142_, _07142_, _07142_, _07142_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22275" *) wt4_sd_data[751:744];
  assign in_wt_data_int16_7 = { cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2228" *) { in_wt_data15, in_wt_data14 };
  assign _04617_ = { _07143_, _07143_, _07143_, _07143_, _07143_, _07143_, _07143_, _07143_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22285" *) wt4_sd_data[759:752];
  assign in_wt_data_int16_6 = { cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2229" *) { in_wt_data13, in_wt_data12 };
  assign _04618_ = { _07144_, _07144_, _07144_, _07144_, _07144_, _07144_, _07144_, _07144_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22295" *) wt4_sd_data[767:760];
  assign in_wt_data_int16_5 = { cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2230" *) { in_wt_data11, in_wt_data10 };
  assign _04619_ = { _07145_, _07145_, _07145_, _07145_, _07145_, _07145_, _07145_, _07145_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22305" *) wt4_sd_data[775:768];
  assign in_wt_data_int16_4 = { cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2231" *) { in_wt_data9, in_wt_data8 };
  assign _04620_ = { _07146_, _07146_, _07146_, _07146_, _07146_, _07146_, _07146_, _07146_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22315" *) wt4_sd_data[783:776];
  assign in_wt_data_int16_3 = { cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2232" *) { in_wt_data7, in_wt_data6 };
  assign _04621_ = { _07147_, _07147_, _07147_, _07147_, _07147_, _07147_, _07147_, _07147_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22325" *) wt4_sd_data[791:784];
  assign in_wt_data_int16_2 = { cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2233" *) { in_wt_data5, in_wt_data4 };
  assign _04622_ = { _07148_, _07148_, _07148_, _07148_, _07148_, _07148_, _07148_, _07148_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22335" *) wt4_sd_data[799:792];
  assign in_wt_data_int16_1 = { cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2234" *) { in_wt_data3, in_wt_data2 };
  assign _04623_ = { _07149_, _07149_, _07149_, _07149_, _07149_, _07149_, _07149_, _07149_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22345" *) wt4_sd_data[807:800];
  assign in_wt_data_int16_0 = { cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2235" *) { in_wt_data1, in_wt_data0 };
  assign _04624_ = { _07150_, _07150_, _07150_, _07150_, _07150_, _07150_, _07150_, _07150_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22355" *) wt4_sd_data[815:808];
  assign _04625_ = { _07151_, _07151_, _07151_, _07151_, _07151_, _07151_, _07151_, _07151_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22365" *) wt4_sd_data[823:816];
  assign _04626_ = { _07152_, _07152_, _07152_, _07152_, _07152_, _07152_, _07152_, _07152_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22375" *) wt4_sd_data[831:824];
  assign _04627_ = { _07153_, _07153_, _07153_, _07153_, _07153_, _07153_, _07153_, _07153_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22385" *) wt4_sd_data[839:832];
  assign _04628_ = { _07154_, _07154_, _07154_, _07154_, _07154_, _07154_, _07154_, _07154_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22395" *) wt4_sd_data[847:840];
  assign _04629_ = { _07155_, _07155_, _07155_, _07155_, _07155_, _07155_, _07155_, _07155_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22405" *) wt4_sd_data[855:848];
  assign _04630_ = { _07156_, _07156_, _07156_, _07156_, _07156_, _07156_, _07156_, _07156_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22415" *) wt4_sd_data[863:856];
  assign _04631_ = { _07157_, _07157_, _07157_, _07157_, _07157_, _07157_, _07157_, _07157_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22425" *) wt4_sd_data[871:864];
  assign _04632_ = { _07158_, _07158_, _07158_, _07158_, _07158_, _07158_, _07158_, _07158_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22435" *) wt4_sd_data[879:872];
  assign _04633_ = { _07159_, _07159_, _07159_, _07159_, _07159_, _07159_, _07159_, _07159_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22445" *) wt4_sd_data[887:880];
  assign _04634_ = { _07160_, _07160_, _07160_, _07160_, _07160_, _07160_, _07160_, _07160_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22455" *) wt4_sd_data[895:888];
  assign _04635_ = { _07161_, _07161_, _07161_, _07161_, _07161_, _07161_, _07161_, _07161_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22465" *) wt4_sd_data[903:896];
  assign _04636_ = { _07162_, _07162_, _07162_, _07162_, _07162_, _07162_, _07162_, _07162_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22475" *) wt4_sd_data[911:904];
  assign _04637_ = { _07163_, _07163_, _07163_, _07163_, _07163_, _07163_, _07163_, _07163_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22485" *) wt4_sd_data[919:912];
  assign _04638_ = { _07164_, _07164_, _07164_, _07164_, _07164_, _07164_, _07164_, _07164_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22495" *) wt4_sd_data[927:920];
  assign _04639_ = { _07165_, _07165_, _07165_, _07165_, _07165_, _07165_, _07165_, _07165_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22505" *) wt4_sd_data[935:928];
  assign _04640_ = { _07166_, _07166_, _07166_, _07166_, _07166_, _07166_, _07166_, _07166_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22515" *) wt4_sd_data[943:936];
  assign _04641_ = { _07167_, _07167_, _07167_, _07167_, _07167_, _07167_, _07167_, _07167_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22525" *) wt4_sd_data[951:944];
  assign _04642_ = { _07168_, _07168_, _07168_, _07168_, _07168_, _07168_, _07168_, _07168_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22535" *) wt4_sd_data[959:952];
  assign _04643_ = { _07169_, _07169_, _07169_, _07169_, _07169_, _07169_, _07169_, _07169_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22545" *) wt4_sd_data[967:960];
  assign _04644_ = { _07170_, _07170_, _07170_, _07170_, _07170_, _07170_, _07170_, _07170_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22555" *) wt4_sd_data[975:968];
  assign _04645_ = { _07171_, _07171_, _07171_, _07171_, _07171_, _07171_, _07171_, _07171_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22565" *) wt4_sd_data[983:976];
  assign _04646_ = { _07172_, _07172_, _07172_, _07172_, _07172_, _07172_, _07172_, _07172_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22575" *) wt4_sd_data[991:984];
  assign _04647_ = { _07173_, _07173_, _07173_, _07173_, _07173_, _07173_, _07173_, _07173_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22585" *) wt4_sd_data[999:992];
  assign _04648_ = { _07174_, _07174_, _07174_, _07174_, _07174_, _07174_, _07174_, _07174_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22595" *) wt4_sd_data[1007:1000];
  assign _04649_ = { _07175_, _07175_, _07175_, _07175_, _07175_, _07175_, _07175_, _07175_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22605" *) wt4_sd_data[1015:1008];
  assign _04650_ = { _07176_, _07176_, _07176_, _07176_, _07176_, _07176_, _07176_, _07176_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22615" *) wt4_sd_data[1023:1016];
  assign _04651_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22648" *) wt5_actv_pvld_w;
  assign _04652_ = _04651_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22658" *) cfg_is_fp16_d1[79];
  assign _04653_ = { _07177_, _07177_, _07177_, _07177_, _07177_, _07177_, _07177_, _07177_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22669" *) wt5_sd_data[7:0];
  assign _04654_ = { _07178_, _07178_, _07178_, _07178_, _07178_, _07178_, _07178_, _07178_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22679" *) wt5_sd_data[15:8];
  assign _04655_ = { _07179_, _07179_, _07179_, _07179_, _07179_, _07179_, _07179_, _07179_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22689" *) wt5_sd_data[23:16];
  assign _04656_ = { _07180_, _07180_, _07180_, _07180_, _07180_, _07180_, _07180_, _07180_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22699" *) wt5_sd_data[31:24];
  assign _04657_ = { _07181_, _07181_, _07181_, _07181_, _07181_, _07181_, _07181_, _07181_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22709" *) wt5_sd_data[39:32];
  assign _04658_ = { _07182_, _07182_, _07182_, _07182_, _07182_, _07182_, _07182_, _07182_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22719" *) wt5_sd_data[47:40];
  assign _04659_ = { _07183_, _07183_, _07183_, _07183_, _07183_, _07183_, _07183_, _07183_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22729" *) wt5_sd_data[55:48];
  assign _04660_ = { _07184_, _07184_, _07184_, _07184_, _07184_, _07184_, _07184_, _07184_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22739" *) wt5_sd_data[63:56];
  assign _04661_ = { _07185_, _07185_, _07185_, _07185_, _07185_, _07185_, _07185_, _07185_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22749" *) wt5_sd_data[71:64];
  assign _04662_ = { _07186_, _07186_, _07186_, _07186_, _07186_, _07186_, _07186_, _07186_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22759" *) wt5_sd_data[79:72];
  assign _04663_ = { _07187_, _07187_, _07187_, _07187_, _07187_, _07187_, _07187_, _07187_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22769" *) wt5_sd_data[87:80];
  assign _04664_ = { _07188_, _07188_, _07188_, _07188_, _07188_, _07188_, _07188_, _07188_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22779" *) wt5_sd_data[95:88];
  assign _04665_ = { _07189_, _07189_, _07189_, _07189_, _07189_, _07189_, _07189_, _07189_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22789" *) wt5_sd_data[103:96];
  assign _04666_ = { _07190_, _07190_, _07190_, _07190_, _07190_, _07190_, _07190_, _07190_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22799" *) wt5_sd_data[111:104];
  assign _04667_ = { _07191_, _07191_, _07191_, _07191_, _07191_, _07191_, _07191_, _07191_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22809" *) wt5_sd_data[119:112];
  assign _04668_ = { _07192_, _07192_, _07192_, _07192_, _07192_, _07192_, _07192_, _07192_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22819" *) wt5_sd_data[127:120];
  assign _04669_ = { _07193_, _07193_, _07193_, _07193_, _07193_, _07193_, _07193_, _07193_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22829" *) wt5_sd_data[135:128];
  assign _04670_ = { _07194_, _07194_, _07194_, _07194_, _07194_, _07194_, _07194_, _07194_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22839" *) wt5_sd_data[143:136];
  assign _04671_ = { _07195_, _07195_, _07195_, _07195_, _07195_, _07195_, _07195_, _07195_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22849" *) wt5_sd_data[151:144];
  assign _04672_ = { _07196_, _07196_, _07196_, _07196_, _07196_, _07196_, _07196_, _07196_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22859" *) wt5_sd_data[159:152];
  assign _04673_ = { _07197_, _07197_, _07197_, _07197_, _07197_, _07197_, _07197_, _07197_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22869" *) wt5_sd_data[167:160];
  assign _04674_ = { _07198_, _07198_, _07198_, _07198_, _07198_, _07198_, _07198_, _07198_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22879" *) wt5_sd_data[175:168];
  assign _04675_ = { _07199_, _07199_, _07199_, _07199_, _07199_, _07199_, _07199_, _07199_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22889" *) wt5_sd_data[183:176];
  assign _04676_ = { _07200_, _07200_, _07200_, _07200_, _07200_, _07200_, _07200_, _07200_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22899" *) wt5_sd_data[191:184];
  assign _04677_ = { _07201_, _07201_, _07201_, _07201_, _07201_, _07201_, _07201_, _07201_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22909" *) wt5_sd_data[199:192];
  assign _04678_ = { _07202_, _07202_, _07202_, _07202_, _07202_, _07202_, _07202_, _07202_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22919" *) wt5_sd_data[207:200];
  assign _04679_ = { _07203_, _07203_, _07203_, _07203_, _07203_, _07203_, _07203_, _07203_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22929" *) wt5_sd_data[215:208];
  assign _04680_ = { _07204_, _07204_, _07204_, _07204_, _07204_, _07204_, _07204_, _07204_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22939" *) wt5_sd_data[223:216];
  assign _04681_ = { _07205_, _07205_, _07205_, _07205_, _07205_, _07205_, _07205_, _07205_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22949" *) wt5_sd_data[231:224];
  assign _04682_ = { _07206_, _07206_, _07206_, _07206_, _07206_, _07206_, _07206_, _07206_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22959" *) wt5_sd_data[239:232];
  assign _04683_ = { _07207_, _07207_, _07207_, _07207_, _07207_, _07207_, _07207_, _07207_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22969" *) wt5_sd_data[247:240];
  assign _04684_ = { _07208_, _07208_, _07208_, _07208_, _07208_, _07208_, _07208_, _07208_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22979" *) wt5_sd_data[255:248];
  assign _04685_ = { _07209_, _07209_, _07209_, _07209_, _07209_, _07209_, _07209_, _07209_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22989" *) wt5_sd_data[263:256];
  assign _04686_ = { _07210_, _07210_, _07210_, _07210_, _07210_, _07210_, _07210_, _07210_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22999" *) wt5_sd_data[271:264];
  assign _04687_ = { _07211_, _07211_, _07211_, _07211_, _07211_, _07211_, _07211_, _07211_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23009" *) wt5_sd_data[279:272];
  assign _04688_ = { _07212_, _07212_, _07212_, _07212_, _07212_, _07212_, _07212_, _07212_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23019" *) wt5_sd_data[287:280];
  assign _04689_ = { _07213_, _07213_, _07213_, _07213_, _07213_, _07213_, _07213_, _07213_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23029" *) wt5_sd_data[295:288];
  assign _04690_ = { _07214_, _07214_, _07214_, _07214_, _07214_, _07214_, _07214_, _07214_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23039" *) wt5_sd_data[303:296];
  assign _04691_ = { _07215_, _07215_, _07215_, _07215_, _07215_, _07215_, _07215_, _07215_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23049" *) wt5_sd_data[311:304];
  assign _04692_ = { _07216_, _07216_, _07216_, _07216_, _07216_, _07216_, _07216_, _07216_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23059" *) wt5_sd_data[319:312];
  assign _04693_ = { _07217_, _07217_, _07217_, _07217_, _07217_, _07217_, _07217_, _07217_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23069" *) wt5_sd_data[327:320];
  assign _04694_ = { _07218_, _07218_, _07218_, _07218_, _07218_, _07218_, _07218_, _07218_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23079" *) wt5_sd_data[335:328];
  assign _04695_ = { _07219_, _07219_, _07219_, _07219_, _07219_, _07219_, _07219_, _07219_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23089" *) wt5_sd_data[343:336];
  assign _04696_ = { _07220_, _07220_, _07220_, _07220_, _07220_, _07220_, _07220_, _07220_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23099" *) wt5_sd_data[351:344];
  assign _04697_ = { _07221_, _07221_, _07221_, _07221_, _07221_, _07221_, _07221_, _07221_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23109" *) wt5_sd_data[359:352];
  assign _04698_ = { _07222_, _07222_, _07222_, _07222_, _07222_, _07222_, _07222_, _07222_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23119" *) wt5_sd_data[367:360];
  assign _04699_ = { _07223_, _07223_, _07223_, _07223_, _07223_, _07223_, _07223_, _07223_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23129" *) wt5_sd_data[375:368];
  assign _04700_ = { _07224_, _07224_, _07224_, _07224_, _07224_, _07224_, _07224_, _07224_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23139" *) wt5_sd_data[383:376];
  assign _04701_ = { _07225_, _07225_, _07225_, _07225_, _07225_, _07225_, _07225_, _07225_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23149" *) wt5_sd_data[391:384];
  assign _04702_ = { _07226_, _07226_, _07226_, _07226_, _07226_, _07226_, _07226_, _07226_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23159" *) wt5_sd_data[399:392];
  assign _04703_ = { _07227_, _07227_, _07227_, _07227_, _07227_, _07227_, _07227_, _07227_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23169" *) wt5_sd_data[407:400];
  assign _04704_ = { _07228_, _07228_, _07228_, _07228_, _07228_, _07228_, _07228_, _07228_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23179" *) wt5_sd_data[415:408];
  assign _04705_ = { _07229_, _07229_, _07229_, _07229_, _07229_, _07229_, _07229_, _07229_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23189" *) wt5_sd_data[423:416];
  assign _04706_ = { _07230_, _07230_, _07230_, _07230_, _07230_, _07230_, _07230_, _07230_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23199" *) wt5_sd_data[431:424];
  assign _04707_ = { _07231_, _07231_, _07231_, _07231_, _07231_, _07231_, _07231_, _07231_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23209" *) wt5_sd_data[439:432];
  assign _04708_ = { _07232_, _07232_, _07232_, _07232_, _07232_, _07232_, _07232_, _07232_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23219" *) wt5_sd_data[447:440];
  assign _04709_ = { _07233_, _07233_, _07233_, _07233_, _07233_, _07233_, _07233_, _07233_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23229" *) wt5_sd_data[455:448];
  assign _04710_ = { _07234_, _07234_, _07234_, _07234_, _07234_, _07234_, _07234_, _07234_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23239" *) wt5_sd_data[463:456];
  assign _04711_ = { _07235_, _07235_, _07235_, _07235_, _07235_, _07235_, _07235_, _07235_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23249" *) wt5_sd_data[471:464];
  assign _04712_ = { _07236_, _07236_, _07236_, _07236_, _07236_, _07236_, _07236_, _07236_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23259" *) wt5_sd_data[479:472];
  assign _04713_ = { _07237_, _07237_, _07237_, _07237_, _07237_, _07237_, _07237_, _07237_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23269" *) wt5_sd_data[487:480];
  assign _04714_ = { _07238_, _07238_, _07238_, _07238_, _07238_, _07238_, _07238_, _07238_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23279" *) wt5_sd_data[495:488];
  assign _04715_ = { _07239_, _07239_, _07239_, _07239_, _07239_, _07239_, _07239_, _07239_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23289" *) wt5_sd_data[503:496];
  assign _04716_ = { _07240_, _07240_, _07240_, _07240_, _07240_, _07240_, _07240_, _07240_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23299" *) wt5_sd_data[511:504];
  assign _04717_ = { _07241_, _07241_, _07241_, _07241_, _07241_, _07241_, _07241_, _07241_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23309" *) wt5_sd_data[519:512];
  assign _04718_ = { _07242_, _07242_, _07242_, _07242_, _07242_, _07242_, _07242_, _07242_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23319" *) wt5_sd_data[527:520];
  assign _04719_ = { _07243_, _07243_, _07243_, _07243_, _07243_, _07243_, _07243_, _07243_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23329" *) wt5_sd_data[535:528];
  assign _04720_ = { _07244_, _07244_, _07244_, _07244_, _07244_, _07244_, _07244_, _07244_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23339" *) wt5_sd_data[543:536];
  assign _04721_ = { _07245_, _07245_, _07245_, _07245_, _07245_, _07245_, _07245_, _07245_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23349" *) wt5_sd_data[551:544];
  assign _04722_ = { _07246_, _07246_, _07246_, _07246_, _07246_, _07246_, _07246_, _07246_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23359" *) wt5_sd_data[559:552];
  assign _04723_ = { _07247_, _07247_, _07247_, _07247_, _07247_, _07247_, _07247_, _07247_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23369" *) wt5_sd_data[567:560];
  assign _04724_ = { _07248_, _07248_, _07248_, _07248_, _07248_, _07248_, _07248_, _07248_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23379" *) wt5_sd_data[575:568];
  assign _04725_ = { _07249_, _07249_, _07249_, _07249_, _07249_, _07249_, _07249_, _07249_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23389" *) wt5_sd_data[583:576];
  assign _04726_ = { _07250_, _07250_, _07250_, _07250_, _07250_, _07250_, _07250_, _07250_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23399" *) wt5_sd_data[591:584];
  assign _04727_ = { _07251_, _07251_, _07251_, _07251_, _07251_, _07251_, _07251_, _07251_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23409" *) wt5_sd_data[599:592];
  assign _04728_ = { _07252_, _07252_, _07252_, _07252_, _07252_, _07252_, _07252_, _07252_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23419" *) wt5_sd_data[607:600];
  assign _04729_ = { _07253_, _07253_, _07253_, _07253_, _07253_, _07253_, _07253_, _07253_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23429" *) wt5_sd_data[615:608];
  assign _04730_ = { _07254_, _07254_, _07254_, _07254_, _07254_, _07254_, _07254_, _07254_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23439" *) wt5_sd_data[623:616];
  assign _04731_ = { _07255_, _07255_, _07255_, _07255_, _07255_, _07255_, _07255_, _07255_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23449" *) wt5_sd_data[631:624];
  assign _04732_ = { _07256_, _07256_, _07256_, _07256_, _07256_, _07256_, _07256_, _07256_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23459" *) wt5_sd_data[639:632];
  assign _04733_ = { _07257_, _07257_, _07257_, _07257_, _07257_, _07257_, _07257_, _07257_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23469" *) wt5_sd_data[647:640];
  assign _04734_ = { _07258_, _07258_, _07258_, _07258_, _07258_, _07258_, _07258_, _07258_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23479" *) wt5_sd_data[655:648];
  assign _04735_ = { _07259_, _07259_, _07259_, _07259_, _07259_, _07259_, _07259_, _07259_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23489" *) wt5_sd_data[663:656];
  assign _04736_ = { _07260_, _07260_, _07260_, _07260_, _07260_, _07260_, _07260_, _07260_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23499" *) wt5_sd_data[671:664];
  assign _04737_ = { _07261_, _07261_, _07261_, _07261_, _07261_, _07261_, _07261_, _07261_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23509" *) wt5_sd_data[679:672];
  assign _04738_ = { _07262_, _07262_, _07262_, _07262_, _07262_, _07262_, _07262_, _07262_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23519" *) wt5_sd_data[687:680];
  assign _04739_ = { _07263_, _07263_, _07263_, _07263_, _07263_, _07263_, _07263_, _07263_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23529" *) wt5_sd_data[695:688];
  assign _04740_ = { _07264_, _07264_, _07264_, _07264_, _07264_, _07264_, _07264_, _07264_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23539" *) wt5_sd_data[703:696];
  assign _04741_ = { _07265_, _07265_, _07265_, _07265_, _07265_, _07265_, _07265_, _07265_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23549" *) wt5_sd_data[711:704];
  assign _04742_ = { _07266_, _07266_, _07266_, _07266_, _07266_, _07266_, _07266_, _07266_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23559" *) wt5_sd_data[719:712];
  assign _04743_ = { _07267_, _07267_, _07267_, _07267_, _07267_, _07267_, _07267_, _07267_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23569" *) wt5_sd_data[727:720];
  assign _04744_ = { _07268_, _07268_, _07268_, _07268_, _07268_, _07268_, _07268_, _07268_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23579" *) wt5_sd_data[735:728];
  assign _04745_ = { _07269_, _07269_, _07269_, _07269_, _07269_, _07269_, _07269_, _07269_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23589" *) wt5_sd_data[743:736];
  assign _04746_ = { _07270_, _07270_, _07270_, _07270_, _07270_, _07270_, _07270_, _07270_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23599" *) wt5_sd_data[751:744];
  assign _04747_ = { _07271_, _07271_, _07271_, _07271_, _07271_, _07271_, _07271_, _07271_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23609" *) wt5_sd_data[759:752];
  assign _04748_ = { _07272_, _07272_, _07272_, _07272_, _07272_, _07272_, _07272_, _07272_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23619" *) wt5_sd_data[767:760];
  assign _04749_ = { _07273_, _07273_, _07273_, _07273_, _07273_, _07273_, _07273_, _07273_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23629" *) wt5_sd_data[775:768];
  assign _04750_ = { _07274_, _07274_, _07274_, _07274_, _07274_, _07274_, _07274_, _07274_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23639" *) wt5_sd_data[783:776];
  assign _04751_ = { _07275_, _07275_, _07275_, _07275_, _07275_, _07275_, _07275_, _07275_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23649" *) wt5_sd_data[791:784];
  assign _04752_ = { _07276_, _07276_, _07276_, _07276_, _07276_, _07276_, _07276_, _07276_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23659" *) wt5_sd_data[799:792];
  assign _04753_ = { _07277_, _07277_, _07277_, _07277_, _07277_, _07277_, _07277_, _07277_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23669" *) wt5_sd_data[807:800];
  assign _04754_ = { _07278_, _07278_, _07278_, _07278_, _07278_, _07278_, _07278_, _07278_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23679" *) wt5_sd_data[815:808];
  assign _04755_ = { _07279_, _07279_, _07279_, _07279_, _07279_, _07279_, _07279_, _07279_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23689" *) wt5_sd_data[823:816];
  assign _04756_ = { _07280_, _07280_, _07280_, _07280_, _07280_, _07280_, _07280_, _07280_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23699" *) wt5_sd_data[831:824];
  assign _04757_ = { _07281_, _07281_, _07281_, _07281_, _07281_, _07281_, _07281_, _07281_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23709" *) wt5_sd_data[839:832];
  assign _04758_ = { _07282_, _07282_, _07282_, _07282_, _07282_, _07282_, _07282_, _07282_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23719" *) wt5_sd_data[847:840];
  assign _04759_ = { _07283_, _07283_, _07283_, _07283_, _07283_, _07283_, _07283_, _07283_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23729" *) wt5_sd_data[855:848];
  assign _04760_ = { _07284_, _07284_, _07284_, _07284_, _07284_, _07284_, _07284_, _07284_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23739" *) wt5_sd_data[863:856];
  assign _04761_ = { _07285_, _07285_, _07285_, _07285_, _07285_, _07285_, _07285_, _07285_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23749" *) wt5_sd_data[871:864];
  assign _04762_ = { _07286_, _07286_, _07286_, _07286_, _07286_, _07286_, _07286_, _07286_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23759" *) wt5_sd_data[879:872];
  assign _04763_ = { _07287_, _07287_, _07287_, _07287_, _07287_, _07287_, _07287_, _07287_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23769" *) wt5_sd_data[887:880];
  assign _04764_ = { _07288_, _07288_, _07288_, _07288_, _07288_, _07288_, _07288_, _07288_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23779" *) wt5_sd_data[895:888];
  assign _04765_ = { _07289_, _07289_, _07289_, _07289_, _07289_, _07289_, _07289_, _07289_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23789" *) wt5_sd_data[903:896];
  assign _04766_ = { _07290_, _07290_, _07290_, _07290_, _07290_, _07290_, _07290_, _07290_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23799" *) wt5_sd_data[911:904];
  assign _04767_ = { _07291_, _07291_, _07291_, _07291_, _07291_, _07291_, _07291_, _07291_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23809" *) wt5_sd_data[919:912];
  assign _04768_ = { _07292_, _07292_, _07292_, _07292_, _07292_, _07292_, _07292_, _07292_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23819" *) wt5_sd_data[927:920];
  assign _04769_ = { _07293_, _07293_, _07293_, _07293_, _07293_, _07293_, _07293_, _07293_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23829" *) wt5_sd_data[935:928];
  assign _04770_ = { _07294_, _07294_, _07294_, _07294_, _07294_, _07294_, _07294_, _07294_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23839" *) wt5_sd_data[943:936];
  assign _04771_ = { _07295_, _07295_, _07295_, _07295_, _07295_, _07295_, _07295_, _07295_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23849" *) wt5_sd_data[951:944];
  assign _04772_ = { _07296_, _07296_, _07296_, _07296_, _07296_, _07296_, _07296_, _07296_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23859" *) wt5_sd_data[959:952];
  assign _04773_ = { _07297_, _07297_, _07297_, _07297_, _07297_, _07297_, _07297_, _07297_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23869" *) wt5_sd_data[967:960];
  assign _04774_ = { _07298_, _07298_, _07298_, _07298_, _07298_, _07298_, _07298_, _07298_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23879" *) wt5_sd_data[975:968];
  assign _04775_ = { _07299_, _07299_, _07299_, _07299_, _07299_, _07299_, _07299_, _07299_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23889" *) wt5_sd_data[983:976];
  assign _04776_ = { _07300_, _07300_, _07300_, _07300_, _07300_, _07300_, _07300_, _07300_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23899" *) wt5_sd_data[991:984];
  assign _04777_ = { _07301_, _07301_, _07301_, _07301_, _07301_, _07301_, _07301_, _07301_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23909" *) wt5_sd_data[999:992];
  assign _04778_ = { _07302_, _07302_, _07302_, _07302_, _07302_, _07302_, _07302_, _07302_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23919" *) wt5_sd_data[1007:1000];
  assign _04779_ = { _07303_, _07303_, _07303_, _07303_, _07303_, _07303_, _07303_, _07303_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23929" *) wt5_sd_data[1015:1008];
  assign _04780_ = { _07304_, _07304_, _07304_, _07304_, _07304_, _07304_, _07304_, _07304_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23939" *) wt5_sd_data[1023:1016];
  assign _04781_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23972" *) wt6_actv_pvld_w;
  assign _04782_ = _04781_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23982" *) cfg_is_fp16_d1[80];
  assign _04783_ = { _07305_, _07305_, _07305_, _07305_, _07305_, _07305_, _07305_, _07305_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23993" *) wt6_sd_data[7:0];
  assign _04784_ = { _07306_, _07306_, _07306_, _07306_, _07306_, _07306_, _07306_, _07306_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24003" *) wt6_sd_data[15:8];
  assign _04785_ = { _07307_, _07307_, _07307_, _07307_, _07307_, _07307_, _07307_, _07307_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24013" *) wt6_sd_data[23:16];
  assign _04786_ = { _07308_, _07308_, _07308_, _07308_, _07308_, _07308_, _07308_, _07308_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24023" *) wt6_sd_data[31:24];
  assign _04787_ = { _07309_, _07309_, _07309_, _07309_, _07309_, _07309_, _07309_, _07309_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24033" *) wt6_sd_data[39:32];
  assign _04788_ = { _07310_, _07310_, _07310_, _07310_, _07310_, _07310_, _07310_, _07310_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24043" *) wt6_sd_data[47:40];
  assign _04789_ = { _07311_, _07311_, _07311_, _07311_, _07311_, _07311_, _07311_, _07311_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24053" *) wt6_sd_data[55:48];
  assign _04790_ = { _07312_, _07312_, _07312_, _07312_, _07312_, _07312_, _07312_, _07312_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24063" *) wt6_sd_data[63:56];
  assign _04791_ = { _07313_, _07313_, _07313_, _07313_, _07313_, _07313_, _07313_, _07313_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24073" *) wt6_sd_data[71:64];
  assign _04792_ = { _07314_, _07314_, _07314_, _07314_, _07314_, _07314_, _07314_, _07314_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24083" *) wt6_sd_data[79:72];
  assign _04793_ = { _07315_, _07315_, _07315_, _07315_, _07315_, _07315_, _07315_, _07315_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24093" *) wt6_sd_data[87:80];
  assign _04794_ = { _07316_, _07316_, _07316_, _07316_, _07316_, _07316_, _07316_, _07316_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24103" *) wt6_sd_data[95:88];
  assign _04795_ = { _07317_, _07317_, _07317_, _07317_, _07317_, _07317_, _07317_, _07317_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24113" *) wt6_sd_data[103:96];
  assign _04796_ = { _07318_, _07318_, _07318_, _07318_, _07318_, _07318_, _07318_, _07318_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24123" *) wt6_sd_data[111:104];
  assign _04797_ = { _07319_, _07319_, _07319_, _07319_, _07319_, _07319_, _07319_, _07319_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24133" *) wt6_sd_data[119:112];
  assign _04798_ = { _07320_, _07320_, _07320_, _07320_, _07320_, _07320_, _07320_, _07320_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24143" *) wt6_sd_data[127:120];
  assign _04799_ = { _07321_, _07321_, _07321_, _07321_, _07321_, _07321_, _07321_, _07321_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24153" *) wt6_sd_data[135:128];
  assign _04800_ = { _07322_, _07322_, _07322_, _07322_, _07322_, _07322_, _07322_, _07322_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24163" *) wt6_sd_data[143:136];
  assign _04801_ = { _07323_, _07323_, _07323_, _07323_, _07323_, _07323_, _07323_, _07323_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24173" *) wt6_sd_data[151:144];
  assign _04802_ = { _07324_, _07324_, _07324_, _07324_, _07324_, _07324_, _07324_, _07324_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24183" *) wt6_sd_data[159:152];
  assign _04803_ = { _07325_, _07325_, _07325_, _07325_, _07325_, _07325_, _07325_, _07325_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24193" *) wt6_sd_data[167:160];
  assign _04804_ = { _07326_, _07326_, _07326_, _07326_, _07326_, _07326_, _07326_, _07326_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24203" *) wt6_sd_data[175:168];
  assign _04805_ = { _07327_, _07327_, _07327_, _07327_, _07327_, _07327_, _07327_, _07327_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24213" *) wt6_sd_data[183:176];
  assign _04806_ = { _07328_, _07328_, _07328_, _07328_, _07328_, _07328_, _07328_, _07328_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24223" *) wt6_sd_data[191:184];
  assign _04807_ = { _07329_, _07329_, _07329_, _07329_, _07329_, _07329_, _07329_, _07329_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24233" *) wt6_sd_data[199:192];
  assign _04808_ = { _07330_, _07330_, _07330_, _07330_, _07330_, _07330_, _07330_, _07330_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24243" *) wt6_sd_data[207:200];
  assign _04809_ = { _07331_, _07331_, _07331_, _07331_, _07331_, _07331_, _07331_, _07331_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24253" *) wt6_sd_data[215:208];
  assign _04810_ = { _07332_, _07332_, _07332_, _07332_, _07332_, _07332_, _07332_, _07332_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24263" *) wt6_sd_data[223:216];
  assign _04811_ = { _07333_, _07333_, _07333_, _07333_, _07333_, _07333_, _07333_, _07333_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24273" *) wt6_sd_data[231:224];
  assign _04812_ = { _07334_, _07334_, _07334_, _07334_, _07334_, _07334_, _07334_, _07334_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24283" *) wt6_sd_data[239:232];
  assign _04813_ = { _07335_, _07335_, _07335_, _07335_, _07335_, _07335_, _07335_, _07335_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24293" *) wt6_sd_data[247:240];
  assign _04814_ = { _07336_, _07336_, _07336_, _07336_, _07336_, _07336_, _07336_, _07336_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24303" *) wt6_sd_data[255:248];
  assign _04815_ = { _07337_, _07337_, _07337_, _07337_, _07337_, _07337_, _07337_, _07337_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24313" *) wt6_sd_data[263:256];
  assign _04816_ = { _07338_, _07338_, _07338_, _07338_, _07338_, _07338_, _07338_, _07338_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24323" *) wt6_sd_data[271:264];
  assign _04817_ = { _07339_, _07339_, _07339_, _07339_, _07339_, _07339_, _07339_, _07339_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24333" *) wt6_sd_data[279:272];
  assign _04818_ = { _07340_, _07340_, _07340_, _07340_, _07340_, _07340_, _07340_, _07340_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24343" *) wt6_sd_data[287:280];
  assign _04819_ = { _07341_, _07341_, _07341_, _07341_, _07341_, _07341_, _07341_, _07341_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24353" *) wt6_sd_data[295:288];
  assign _04820_ = { _07342_, _07342_, _07342_, _07342_, _07342_, _07342_, _07342_, _07342_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24363" *) wt6_sd_data[303:296];
  assign in_wt_data_int8_63 = { cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2437" *) { in_wt_data127, in_wt_data63 };
  assign _04821_ = { _07343_, _07343_, _07343_, _07343_, _07343_, _07343_, _07343_, _07343_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24373" *) wt6_sd_data[311:304];
  assign in_wt_data_int8_62 = { cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2438" *) { in_wt_data126, in_wt_data62 };
  assign _04822_ = { _07344_, _07344_, _07344_, _07344_, _07344_, _07344_, _07344_, _07344_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24383" *) wt6_sd_data[319:312];
  assign in_wt_data_int8_61 = { cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2439" *) { in_wt_data125, in_wt_data61 };
  assign _04823_ = { _07345_, _07345_, _07345_, _07345_, _07345_, _07345_, _07345_, _07345_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24393" *) wt6_sd_data[327:320];
  assign in_wt_data_int8_60 = { cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2440" *) { in_wt_data124, in_wt_data60 };
  assign _04824_ = { _07346_, _07346_, _07346_, _07346_, _07346_, _07346_, _07346_, _07346_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24403" *) wt6_sd_data[335:328];
  assign in_wt_data_int8_59 = { cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2441" *) { in_wt_data123, in_wt_data59 };
  assign _04825_ = { _07347_, _07347_, _07347_, _07347_, _07347_, _07347_, _07347_, _07347_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24413" *) wt6_sd_data[343:336];
  assign in_wt_data_int8_58 = { cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2442" *) { in_wt_data122, in_wt_data58 };
  assign _04826_ = { _07348_, _07348_, _07348_, _07348_, _07348_, _07348_, _07348_, _07348_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24423" *) wt6_sd_data[351:344];
  assign in_wt_data_int8_57 = { cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2443" *) { in_wt_data121, in_wt_data57 };
  assign _04827_ = { _07349_, _07349_, _07349_, _07349_, _07349_, _07349_, _07349_, _07349_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24433" *) wt6_sd_data[359:352];
  assign in_wt_data_int8_56 = { cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2444" *) { in_wt_data120, in_wt_data56 };
  assign _04828_ = { _07350_, _07350_, _07350_, _07350_, _07350_, _07350_, _07350_, _07350_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24443" *) wt6_sd_data[367:360];
  assign in_wt_data_int8_55 = { cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2445" *) { in_wt_data119, in_wt_data55 };
  assign _04829_ = { _07351_, _07351_, _07351_, _07351_, _07351_, _07351_, _07351_, _07351_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24453" *) wt6_sd_data[375:368];
  assign in_wt_data_int8_54 = { cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2446" *) { in_wt_data118, in_wt_data54 };
  assign _04830_ = { _07352_, _07352_, _07352_, _07352_, _07352_, _07352_, _07352_, _07352_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24463" *) wt6_sd_data[383:376];
  assign in_wt_data_int8_53 = { cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2447" *) { in_wt_data117, in_wt_data53 };
  assign _04831_ = { _07353_, _07353_, _07353_, _07353_, _07353_, _07353_, _07353_, _07353_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24473" *) wt6_sd_data[391:384];
  assign in_wt_data_int8_52 = { cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2448" *) { in_wt_data116, in_wt_data52 };
  assign _04832_ = { _07354_, _07354_, _07354_, _07354_, _07354_, _07354_, _07354_, _07354_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24483" *) wt6_sd_data[399:392];
  assign in_wt_data_int8_51 = { cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2449" *) { in_wt_data115, in_wt_data51 };
  assign _04833_ = { _07355_, _07355_, _07355_, _07355_, _07355_, _07355_, _07355_, _07355_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24493" *) wt6_sd_data[407:400];
  assign in_wt_data_int8_50 = { cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2450" *) { in_wt_data114, in_wt_data50 };
  assign _04834_ = { _07356_, _07356_, _07356_, _07356_, _07356_, _07356_, _07356_, _07356_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24503" *) wt6_sd_data[415:408];
  assign in_wt_data_int8_49 = { cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2451" *) { in_wt_data113, in_wt_data49 };
  assign _04835_ = { _07357_, _07357_, _07357_, _07357_, _07357_, _07357_, _07357_, _07357_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24513" *) wt6_sd_data[423:416];
  assign in_wt_data_int8_48 = { cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2452" *) { in_wt_data112, in_wt_data48 };
  assign _04836_ = { _07358_, _07358_, _07358_, _07358_, _07358_, _07358_, _07358_, _07358_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24523" *) wt6_sd_data[431:424];
  assign in_wt_data_int8_47 = { cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2453" *) { in_wt_data111, in_wt_data47 };
  assign _04837_ = { _07359_, _07359_, _07359_, _07359_, _07359_, _07359_, _07359_, _07359_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24533" *) wt6_sd_data[439:432];
  assign in_wt_data_int8_46 = { cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2454" *) { in_wt_data110, in_wt_data46 };
  assign _04838_ = { _07360_, _07360_, _07360_, _07360_, _07360_, _07360_, _07360_, _07360_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24543" *) wt6_sd_data[447:440];
  assign in_wt_data_int8_45 = { cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2455" *) { in_wt_data109, in_wt_data45 };
  assign _04839_ = { _07361_, _07361_, _07361_, _07361_, _07361_, _07361_, _07361_, _07361_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24553" *) wt6_sd_data[455:448];
  assign in_wt_data_int8_44 = { cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2456" *) { in_wt_data108, in_wt_data44 };
  assign _04840_ = { _07362_, _07362_, _07362_, _07362_, _07362_, _07362_, _07362_, _07362_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24563" *) wt6_sd_data[463:456];
  assign in_wt_data_int8_43 = { cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2457" *) { in_wt_data107, in_wt_data43 };
  assign _04841_ = { _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24573" *) wt6_sd_data[471:464];
  assign in_wt_data_int8_42 = { cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2458" *) { in_wt_data106, in_wt_data42 };
  assign _04842_ = { _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24583" *) wt6_sd_data[479:472];
  assign in_wt_data_int8_41 = { cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2459" *) { in_wt_data105, in_wt_data41 };
  assign _04843_ = { _07365_, _07365_, _07365_, _07365_, _07365_, _07365_, _07365_, _07365_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24593" *) wt6_sd_data[487:480];
  assign in_wt_data_int8_40 = { cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2460" *) { in_wt_data104, in_wt_data40 };
  assign _04844_ = { _07366_, _07366_, _07366_, _07366_, _07366_, _07366_, _07366_, _07366_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24603" *) wt6_sd_data[495:488];
  assign in_wt_data_int8_39 = { cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2461" *) { in_wt_data103, in_wt_data39 };
  assign _04845_ = { _07367_, _07367_, _07367_, _07367_, _07367_, _07367_, _07367_, _07367_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24613" *) wt6_sd_data[503:496];
  assign in_wt_data_int8_38 = { cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2462" *) { in_wt_data102, in_wt_data38 };
  assign _04846_ = { _07368_, _07368_, _07368_, _07368_, _07368_, _07368_, _07368_, _07368_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24623" *) wt6_sd_data[511:504];
  assign in_wt_data_int8_37 = { cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2463" *) { in_wt_data101, in_wt_data37 };
  assign _04847_ = { _07369_, _07369_, _07369_, _07369_, _07369_, _07369_, _07369_, _07369_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24633" *) wt6_sd_data[519:512];
  assign in_wt_data_int8_36 = { cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2464" *) { in_wt_data100, in_wt_data36 };
  assign _04848_ = { _07370_, _07370_, _07370_, _07370_, _07370_, _07370_, _07370_, _07370_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24643" *) wt6_sd_data[527:520];
  assign in_wt_data_int8_35 = { cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2465" *) { in_wt_data99, in_wt_data35 };
  assign _04849_ = { _07371_, _07371_, _07371_, _07371_, _07371_, _07371_, _07371_, _07371_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24653" *) wt6_sd_data[535:528];
  assign in_wt_data_int8_34 = { cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2466" *) { in_wt_data98, in_wt_data34 };
  assign _04850_ = { _07372_, _07372_, _07372_, _07372_, _07372_, _07372_, _07372_, _07372_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24663" *) wt6_sd_data[543:536];
  assign in_wt_data_int8_33 = { cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2467" *) { in_wt_data97, in_wt_data33 };
  assign _04851_ = { _07373_, _07373_, _07373_, _07373_, _07373_, _07373_, _07373_, _07373_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24673" *) wt6_sd_data[551:544];
  assign in_wt_data_int8_32 = { cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2468" *) { in_wt_data96, in_wt_data32 };
  assign _04852_ = { _07374_, _07374_, _07374_, _07374_, _07374_, _07374_, _07374_, _07374_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24683" *) wt6_sd_data[559:552];
  assign in_wt_data_int8_31 = { cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2469" *) { in_wt_data95, in_wt_data31 };
  assign _04853_ = { _07375_, _07375_, _07375_, _07375_, _07375_, _07375_, _07375_, _07375_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24693" *) wt6_sd_data[567:560];
  assign in_wt_data_int8_30 = { cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2470" *) { in_wt_data94, in_wt_data30 };
  assign _04854_ = { _07376_, _07376_, _07376_, _07376_, _07376_, _07376_, _07376_, _07376_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24703" *) wt6_sd_data[575:568];
  assign in_wt_data_int8_29 = { cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2471" *) { in_wt_data93, in_wt_data29 };
  assign _04855_ = { _07377_, _07377_, _07377_, _07377_, _07377_, _07377_, _07377_, _07377_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24713" *) wt6_sd_data[583:576];
  assign in_wt_data_int8_28 = { cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2472" *) { in_wt_data92, in_wt_data28 };
  assign _04856_ = { _07378_, _07378_, _07378_, _07378_, _07378_, _07378_, _07378_, _07378_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24723" *) wt6_sd_data[591:584];
  assign in_wt_data_int8_27 = { cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2473" *) { in_wt_data91, in_wt_data27 };
  assign _04857_ = { _07379_, _07379_, _07379_, _07379_, _07379_, _07379_, _07379_, _07379_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24733" *) wt6_sd_data[599:592];
  assign in_wt_data_int8_26 = { cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2474" *) { in_wt_data90, in_wt_data26 };
  assign _04858_ = { _07380_, _07380_, _07380_, _07380_, _07380_, _07380_, _07380_, _07380_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24743" *) wt6_sd_data[607:600];
  assign in_wt_data_int8_25 = { cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2475" *) { in_wt_data89, in_wt_data25 };
  assign _04859_ = { _07381_, _07381_, _07381_, _07381_, _07381_, _07381_, _07381_, _07381_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24753" *) wt6_sd_data[615:608];
  assign in_wt_data_int8_24 = { cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2476" *) { in_wt_data88, in_wt_data24 };
  assign _04860_ = { _07382_, _07382_, _07382_, _07382_, _07382_, _07382_, _07382_, _07382_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24763" *) wt6_sd_data[623:616];
  assign in_wt_data_int8_23 = { cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2477" *) { in_wt_data87, in_wt_data23 };
  assign _04861_ = { _07383_, _07383_, _07383_, _07383_, _07383_, _07383_, _07383_, _07383_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24773" *) wt6_sd_data[631:624];
  assign in_wt_data_int8_22 = { cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2478" *) { in_wt_data86, in_wt_data22 };
  assign _04862_ = { _07384_, _07384_, _07384_, _07384_, _07384_, _07384_, _07384_, _07384_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24783" *) wt6_sd_data[639:632];
  assign in_wt_data_int8_21 = { cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2479" *) { in_wt_data85, in_wt_data21 };
  assign _04863_ = { _07385_, _07385_, _07385_, _07385_, _07385_, _07385_, _07385_, _07385_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24793" *) wt6_sd_data[647:640];
  assign in_wt_data_int8_20 = { cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2480" *) { in_wt_data84, in_wt_data20 };
  assign _04864_ = { _07386_, _07386_, _07386_, _07386_, _07386_, _07386_, _07386_, _07386_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24803" *) wt6_sd_data[655:648];
  assign in_wt_data_int8_19 = { cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2481" *) { in_wt_data83, in_wt_data19 };
  assign _04865_ = { _07387_, _07387_, _07387_, _07387_, _07387_, _07387_, _07387_, _07387_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24813" *) wt6_sd_data[663:656];
  assign in_wt_data_int8_18 = { cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2482" *) { in_wt_data82, in_wt_data18 };
  assign _04866_ = { _07388_, _07388_, _07388_, _07388_, _07388_, _07388_, _07388_, _07388_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24823" *) wt6_sd_data[671:664];
  assign in_wt_data_int8_17 = { cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2483" *) { in_wt_data81, in_wt_data17 };
  assign _04867_ = { _07389_, _07389_, _07389_, _07389_, _07389_, _07389_, _07389_, _07389_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24833" *) wt6_sd_data[679:672];
  assign in_wt_data_int8_16 = { cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2484" *) { in_wt_data80, in_wt_data16 };
  assign _04868_ = { _07390_, _07390_, _07390_, _07390_, _07390_, _07390_, _07390_, _07390_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24843" *) wt6_sd_data[687:680];
  assign in_wt_data_int8_15 = { cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2485" *) { in_wt_data79, in_wt_data15 };
  assign _04869_ = { _07391_, _07391_, _07391_, _07391_, _07391_, _07391_, _07391_, _07391_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24853" *) wt6_sd_data[695:688];
  assign in_wt_data_int8_14 = { cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2486" *) { in_wt_data78, in_wt_data14 };
  assign _04870_ = { _07392_, _07392_, _07392_, _07392_, _07392_, _07392_, _07392_, _07392_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24863" *) wt6_sd_data[703:696];
  assign in_wt_data_int8_13 = { cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2487" *) { in_wt_data77, in_wt_data13 };
  assign _04871_ = { _07393_, _07393_, _07393_, _07393_, _07393_, _07393_, _07393_, _07393_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24873" *) wt6_sd_data[711:704];
  assign in_wt_data_int8_12 = { cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2488" *) { in_wt_data76, in_wt_data12 };
  assign _04872_ = { _07394_, _07394_, _07394_, _07394_, _07394_, _07394_, _07394_, _07394_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24883" *) wt6_sd_data[719:712];
  assign in_wt_data_int8_11 = { cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2489" *) { in_wt_data75, in_wt_data11 };
  assign _04873_ = { _07395_, _07395_, _07395_, _07395_, _07395_, _07395_, _07395_, _07395_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24893" *) wt6_sd_data[727:720];
  assign in_wt_data_int8_10 = { cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2490" *) { in_wt_data74, in_wt_data10 };
  assign _04874_ = { _07396_, _07396_, _07396_, _07396_, _07396_, _07396_, _07396_, _07396_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24903" *) wt6_sd_data[735:728];
  assign in_wt_data_int8_9 = { cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2491" *) { in_wt_data73, in_wt_data9 };
  assign _04875_ = { _07397_, _07397_, _07397_, _07397_, _07397_, _07397_, _07397_, _07397_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24913" *) wt6_sd_data[743:736];
  assign in_wt_data_int8_8 = { cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2492" *) { in_wt_data72, in_wt_data8 };
  assign _04876_ = { _07398_, _07398_, _07398_, _07398_, _07398_, _07398_, _07398_, _07398_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24923" *) wt6_sd_data[751:744];
  assign in_wt_data_int8_7 = { cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2493" *) { in_wt_data71, in_wt_data7 };
  assign _04877_ = { _07399_, _07399_, _07399_, _07399_, _07399_, _07399_, _07399_, _07399_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24933" *) wt6_sd_data[759:752];
  assign in_wt_data_int8_6 = { cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2494" *) { in_wt_data70, in_wt_data6 };
  assign _04878_ = { _07400_, _07400_, _07400_, _07400_, _07400_, _07400_, _07400_, _07400_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24943" *) wt6_sd_data[767:760];
  assign in_wt_data_int8_5 = { cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2495" *) { in_wt_data69, in_wt_data5 };
  assign _04879_ = { _07401_, _07401_, _07401_, _07401_, _07401_, _07401_, _07401_, _07401_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24953" *) wt6_sd_data[775:768];
  assign in_wt_data_int8_4 = { cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2496" *) { in_wt_data68, in_wt_data4 };
  assign _04880_ = { _07402_, _07402_, _07402_, _07402_, _07402_, _07402_, _07402_, _07402_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24963" *) wt6_sd_data[783:776];
  assign in_wt_data_int8_3 = { cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2497" *) { in_wt_data67, in_wt_data3 };
  assign _04881_ = { _07403_, _07403_, _07403_, _07403_, _07403_, _07403_, _07403_, _07403_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24973" *) wt6_sd_data[791:784];
  assign in_wt_data_int8_2 = { cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2498" *) { in_wt_data66, in_wt_data2 };
  assign _04882_ = { _07404_, _07404_, _07404_, _07404_, _07404_, _07404_, _07404_, _07404_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24983" *) wt6_sd_data[799:792];
  assign in_wt_data_int8_1 = { cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2499" *) { in_wt_data65, in_wt_data1 };
  assign _04883_ = { _07405_, _07405_, _07405_, _07405_, _07405_, _07405_, _07405_, _07405_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24993" *) wt6_sd_data[807:800];
  assign in_wt_data_int8_0 = { cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2500" *) { in_wt_data64, in_wt_data0 };
  assign _04884_ = { _07406_, _07406_, _07406_, _07406_, _07406_, _07406_, _07406_, _07406_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25003" *) wt6_sd_data[815:808];
  assign _04885_ = { _07407_, _07407_, _07407_, _07407_, _07407_, _07407_, _07407_, _07407_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25013" *) wt6_sd_data[823:816];
  assign _04886_ = { _07408_, _07408_, _07408_, _07408_, _07408_, _07408_, _07408_, _07408_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25023" *) wt6_sd_data[831:824];
  assign _04887_ = { _07409_, _07409_, _07409_, _07409_, _07409_, _07409_, _07409_, _07409_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25033" *) wt6_sd_data[839:832];
  assign _04888_ = { _07410_, _07410_, _07410_, _07410_, _07410_, _07410_, _07410_, _07410_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25043" *) wt6_sd_data[847:840];
  assign _04889_ = { _07411_, _07411_, _07411_, _07411_, _07411_, _07411_, _07411_, _07411_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25053" *) wt6_sd_data[855:848];
  assign _04890_ = { _07412_, _07412_, _07412_, _07412_, _07412_, _07412_, _07412_, _07412_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25063" *) wt6_sd_data[863:856];
  assign _04891_ = { _07413_, _07413_, _07413_, _07413_, _07413_, _07413_, _07413_, _07413_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25073" *) wt6_sd_data[871:864];
  assign _04892_ = { _07414_, _07414_, _07414_, _07414_, _07414_, _07414_, _07414_, _07414_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25083" *) wt6_sd_data[879:872];
  assign _04893_ = { _07415_, _07415_, _07415_, _07415_, _07415_, _07415_, _07415_, _07415_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25093" *) wt6_sd_data[887:880];
  assign _04894_ = { _07416_, _07416_, _07416_, _07416_, _07416_, _07416_, _07416_, _07416_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25103" *) wt6_sd_data[895:888];
  assign _04895_ = { _07417_, _07417_, _07417_, _07417_, _07417_, _07417_, _07417_, _07417_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25113" *) wt6_sd_data[903:896];
  assign _04896_ = { _07418_, _07418_, _07418_, _07418_, _07418_, _07418_, _07418_, _07418_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25123" *) wt6_sd_data[911:904];
  assign _04897_ = { _07419_, _07419_, _07419_, _07419_, _07419_, _07419_, _07419_, _07419_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25133" *) wt6_sd_data[919:912];
  assign _04898_ = { _07420_, _07420_, _07420_, _07420_, _07420_, _07420_, _07420_, _07420_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25143" *) wt6_sd_data[927:920];
  assign _04899_ = { _07421_, _07421_, _07421_, _07421_, _07421_, _07421_, _07421_, _07421_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25153" *) wt6_sd_data[935:928];
  assign _04900_ = { _07422_, _07422_, _07422_, _07422_, _07422_, _07422_, _07422_, _07422_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25163" *) wt6_sd_data[943:936];
  assign _04901_ = { _07423_, _07423_, _07423_, _07423_, _07423_, _07423_, _07423_, _07423_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25173" *) wt6_sd_data[951:944];
  assign _04902_ = { _07424_, _07424_, _07424_, _07424_, _07424_, _07424_, _07424_, _07424_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25183" *) wt6_sd_data[959:952];
  assign _04903_ = { _07425_, _07425_, _07425_, _07425_, _07425_, _07425_, _07425_, _07425_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25193" *) wt6_sd_data[967:960];
  assign _04904_ = { _07426_, _07426_, _07426_, _07426_, _07426_, _07426_, _07426_, _07426_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25203" *) wt6_sd_data[975:968];
  assign _04905_ = { _07427_, _07427_, _07427_, _07427_, _07427_, _07427_, _07427_, _07427_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25213" *) wt6_sd_data[983:976];
  assign _04906_ = { _07428_, _07428_, _07428_, _07428_, _07428_, _07428_, _07428_, _07428_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25223" *) wt6_sd_data[991:984];
  assign _04907_ = { _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25233" *) wt6_sd_data[999:992];
  assign _04908_ = { _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25243" *) wt6_sd_data[1007:1000];
  assign _04909_ = { _07431_, _07431_, _07431_, _07431_, _07431_, _07431_, _07431_, _07431_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25253" *) wt6_sd_data[1015:1008];
  assign _04910_ = { _07432_, _07432_, _07432_, _07432_, _07432_, _07432_, _07432_, _07432_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25263" *) wt6_sd_data[1023:1016];
  assign _04911_ = dat_pre_stripe_st[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25296" *) wt7_actv_pvld_w;
  assign _04912_ = _04911_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25306" *) cfg_is_fp16_d1[81];
  assign _04913_ = { _07433_, _07433_, _07433_, _07433_, _07433_, _07433_, _07433_, _07433_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25317" *) wt7_sd_data[7:0];
  assign _04914_ = { _07434_, _07434_, _07434_, _07434_, _07434_, _07434_, _07434_, _07434_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25327" *) wt7_sd_data[15:8];
  assign _04915_ = { _07435_, _07435_, _07435_, _07435_, _07435_, _07435_, _07435_, _07435_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25337" *) wt7_sd_data[23:16];
  assign _04916_ = { _07436_, _07436_, _07436_, _07436_, _07436_, _07436_, _07436_, _07436_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25347" *) wt7_sd_data[31:24];
  assign _04917_ = { _07437_, _07437_, _07437_, _07437_, _07437_, _07437_, _07437_, _07437_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25357" *) wt7_sd_data[39:32];
  assign _04918_ = { _07438_, _07438_, _07438_, _07438_, _07438_, _07438_, _07438_, _07438_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25367" *) wt7_sd_data[47:40];
  assign _04919_ = { _07439_, _07439_, _07439_, _07439_, _07439_, _07439_, _07439_, _07439_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25377" *) wt7_sd_data[55:48];
  assign _04920_ = { _07440_, _07440_, _07440_, _07440_, _07440_, _07440_, _07440_, _07440_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25387" *) wt7_sd_data[63:56];
  assign _04921_ = { _07441_, _07441_, _07441_, _07441_, _07441_, _07441_, _07441_, _07441_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25397" *) wt7_sd_data[71:64];
  assign _04922_ = { _07442_, _07442_, _07442_, _07442_, _07442_, _07442_, _07442_, _07442_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25407" *) wt7_sd_data[79:72];
  assign _04923_ = { _07443_, _07443_, _07443_, _07443_, _07443_, _07443_, _07443_, _07443_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25417" *) wt7_sd_data[87:80];
  assign _04924_ = { _07444_, _07444_, _07444_, _07444_, _07444_, _07444_, _07444_, _07444_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25427" *) wt7_sd_data[95:88];
  assign _04925_ = { _07445_, _07445_, _07445_, _07445_, _07445_, _07445_, _07445_, _07445_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25437" *) wt7_sd_data[103:96];
  assign _04926_ = { _07446_, _07446_, _07446_, _07446_, _07446_, _07446_, _07446_, _07446_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25447" *) wt7_sd_data[111:104];
  assign _04927_ = { _07447_, _07447_, _07447_, _07447_, _07447_, _07447_, _07447_, _07447_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25457" *) wt7_sd_data[119:112];
  assign _04928_ = { _07448_, _07448_, _07448_, _07448_, _07448_, _07448_, _07448_, _07448_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25467" *) wt7_sd_data[127:120];
  assign _04929_ = { _07449_, _07449_, _07449_, _07449_, _07449_, _07449_, _07449_, _07449_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25477" *) wt7_sd_data[135:128];
  assign _04930_ = { _07450_, _07450_, _07450_, _07450_, _07450_, _07450_, _07450_, _07450_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25487" *) wt7_sd_data[143:136];
  assign _04931_ = { _07451_, _07451_, _07451_, _07451_, _07451_, _07451_, _07451_, _07451_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25497" *) wt7_sd_data[151:144];
  assign _04932_ = { _07452_, _07452_, _07452_, _07452_, _07452_, _07452_, _07452_, _07452_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25507" *) wt7_sd_data[159:152];
  assign _04933_ = { _07453_, _07453_, _07453_, _07453_, _07453_, _07453_, _07453_, _07453_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25517" *) wt7_sd_data[167:160];
  assign _04934_ = { _07454_, _07454_, _07454_, _07454_, _07454_, _07454_, _07454_, _07454_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25527" *) wt7_sd_data[175:168];
  assign _04935_ = { _07455_, _07455_, _07455_, _07455_, _07455_, _07455_, _07455_, _07455_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25537" *) wt7_sd_data[183:176];
  assign _04936_ = { _07456_, _07456_, _07456_, _07456_, _07456_, _07456_, _07456_, _07456_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25547" *) wt7_sd_data[191:184];
  assign _04937_ = { _07457_, _07457_, _07457_, _07457_, _07457_, _07457_, _07457_, _07457_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25557" *) wt7_sd_data[199:192];
  assign _04938_ = { _07458_, _07458_, _07458_, _07458_, _07458_, _07458_, _07458_, _07458_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25567" *) wt7_sd_data[207:200];
  assign _04939_ = { _07459_, _07459_, _07459_, _07459_, _07459_, _07459_, _07459_, _07459_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25577" *) wt7_sd_data[215:208];
  assign _04940_ = { _07460_, _07460_, _07460_, _07460_, _07460_, _07460_, _07460_, _07460_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25587" *) wt7_sd_data[223:216];
  assign _04941_ = { _07461_, _07461_, _07461_, _07461_, _07461_, _07461_, _07461_, _07461_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25597" *) wt7_sd_data[231:224];
  assign _04942_ = { _07462_, _07462_, _07462_, _07462_, _07462_, _07462_, _07462_, _07462_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25607" *) wt7_sd_data[239:232];
  assign _04943_ = { _07463_, _07463_, _07463_, _07463_, _07463_, _07463_, _07463_, _07463_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25617" *) wt7_sd_data[247:240];
  assign _04944_ = { _07464_, _07464_, _07464_, _07464_, _07464_, _07464_, _07464_, _07464_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25627" *) wt7_sd_data[255:248];
  assign _04945_ = { _07465_, _07465_, _07465_, _07465_, _07465_, _07465_, _07465_, _07465_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25637" *) wt7_sd_data[263:256];
  assign _04946_ = { _07466_, _07466_, _07466_, _07466_, _07466_, _07466_, _07466_, _07466_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25647" *) wt7_sd_data[271:264];
  assign _04947_ = { _07467_, _07467_, _07467_, _07467_, _07467_, _07467_, _07467_, _07467_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25657" *) wt7_sd_data[279:272];
  assign _04948_ = { _07468_, _07468_, _07468_, _07468_, _07468_, _07468_, _07468_, _07468_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25667" *) wt7_sd_data[287:280];
  assign _04949_ = { _07469_, _07469_, _07469_, _07469_, _07469_, _07469_, _07469_, _07469_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25677" *) wt7_sd_data[295:288];
  assign _04950_ = { _07470_, _07470_, _07470_, _07470_, _07470_, _07470_, _07470_, _07470_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25687" *) wt7_sd_data[303:296];
  assign _04951_ = { _07471_, _07471_, _07471_, _07471_, _07471_, _07471_, _07471_, _07471_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25697" *) wt7_sd_data[311:304];
  assign _04952_ = { _07472_, _07472_, _07472_, _07472_, _07472_, _07472_, _07472_, _07472_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25707" *) wt7_sd_data[319:312];
  assign _04953_ = { _07473_, _07473_, _07473_, _07473_, _07473_, _07473_, _07473_, _07473_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25717" *) wt7_sd_data[327:320];
  assign _04954_ = { _07474_, _07474_, _07474_, _07474_, _07474_, _07474_, _07474_, _07474_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25727" *) wt7_sd_data[335:328];
  assign _04955_ = { _07475_, _07475_, _07475_, _07475_, _07475_, _07475_, _07475_, _07475_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25737" *) wt7_sd_data[343:336];
  assign _04956_ = { _07476_, _07476_, _07476_, _07476_, _07476_, _07476_, _07476_, _07476_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25747" *) wt7_sd_data[351:344];
  assign _04957_ = { _07477_, _07477_, _07477_, _07477_, _07477_, _07477_, _07477_, _07477_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25757" *) wt7_sd_data[359:352];
  assign _04958_ = { _07478_, _07478_, _07478_, _07478_, _07478_, _07478_, _07478_, _07478_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25767" *) wt7_sd_data[367:360];
  assign _04959_ = { _07479_, _07479_, _07479_, _07479_, _07479_, _07479_, _07479_, _07479_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25777" *) wt7_sd_data[375:368];
  assign _04960_ = { _07480_, _07480_, _07480_, _07480_, _07480_, _07480_, _07480_, _07480_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25787" *) wt7_sd_data[383:376];
  assign _04961_ = { _07481_, _07481_, _07481_, _07481_, _07481_, _07481_, _07481_, _07481_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25797" *) wt7_sd_data[391:384];
  assign _04962_ = { _07482_, _07482_, _07482_, _07482_, _07482_, _07482_, _07482_, _07482_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25807" *) wt7_sd_data[399:392];
  assign _04963_ = { _07483_, _07483_, _07483_, _07483_, _07483_, _07483_, _07483_, _07483_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25817" *) wt7_sd_data[407:400];
  assign _04964_ = { _07484_, _07484_, _07484_, _07484_, _07484_, _07484_, _07484_, _07484_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25827" *) wt7_sd_data[415:408];
  assign _04965_ = { _07485_, _07485_, _07485_, _07485_, _07485_, _07485_, _07485_, _07485_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25837" *) wt7_sd_data[423:416];
  assign _04966_ = { _07486_, _07486_, _07486_, _07486_, _07486_, _07486_, _07486_, _07486_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25847" *) wt7_sd_data[431:424];
  assign _04967_ = { _07487_, _07487_, _07487_, _07487_, _07487_, _07487_, _07487_, _07487_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25857" *) wt7_sd_data[439:432];
  assign _04968_ = { _07488_, _07488_, _07488_, _07488_, _07488_, _07488_, _07488_, _07488_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25867" *) wt7_sd_data[447:440];
  assign _04969_ = { _07489_, _07489_, _07489_, _07489_, _07489_, _07489_, _07489_, _07489_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25877" *) wt7_sd_data[455:448];
  assign _04970_ = cfg_is_fp16_d1[63] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *) _07947_;
  assign _04971_ = _04970_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *) _08075_;
  assign in_wt_nan[63] = _04971_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *) in_wt_mask[126];
  assign _04972_ = { _07490_, _07490_, _07490_, _07490_, _07490_, _07490_, _07490_, _07490_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25887" *) wt7_sd_data[463:456];
  assign _04973_ = cfg_is_fp16_d1[62] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *) _07948_;
  assign _04974_ = _04973_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *) _08076_;
  assign in_wt_nan[62] = _04974_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *) in_wt_mask[124];
  assign _04975_ = { _07491_, _07491_, _07491_, _07491_, _07491_, _07491_, _07491_, _07491_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25897" *) wt7_sd_data[471:464];
  assign _04976_ = cfg_is_fp16_d1[61] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *) _07949_;
  assign _04977_ = _04976_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *) _08077_;
  assign in_wt_nan[61] = _04977_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *) in_wt_mask[122];
  assign _04978_ = { _07492_, _07492_, _07492_, _07492_, _07492_, _07492_, _07492_, _07492_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25907" *) wt7_sd_data[479:472];
  assign _04979_ = cfg_is_fp16_d1[60] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *) _07950_;
  assign _04980_ = _04979_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *) _08078_;
  assign in_wt_nan[60] = _04980_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *) in_wt_mask[120];
  assign _04981_ = { _07493_, _07493_, _07493_, _07493_, _07493_, _07493_, _07493_, _07493_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25917" *) wt7_sd_data[487:480];
  assign _04982_ = cfg_is_fp16_d1[59] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *) _07951_;
  assign _04983_ = _04982_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *) _08079_;
  assign in_wt_nan[59] = _04983_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *) in_wt_mask[118];
  assign _04984_ = { _07494_, _07494_, _07494_, _07494_, _07494_, _07494_, _07494_, _07494_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25927" *) wt7_sd_data[495:488];
  assign _04985_ = cfg_is_fp16_d1[58] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *) _07952_;
  assign _04986_ = _04985_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *) _08080_;
  assign in_wt_nan[58] = _04986_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *) in_wt_mask[116];
  assign _04987_ = { _07495_, _07495_, _07495_, _07495_, _07495_, _07495_, _07495_, _07495_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25937" *) wt7_sd_data[503:496];
  assign _04988_ = cfg_is_fp16_d1[57] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *) _07953_;
  assign _04989_ = _04988_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *) _08081_;
  assign in_wt_nan[57] = _04989_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *) in_wt_mask[114];
  assign _04990_ = { _07496_, _07496_, _07496_, _07496_, _07496_, _07496_, _07496_, _07496_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25947" *) wt7_sd_data[511:504];
  assign _04991_ = cfg_is_fp16_d1[56] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *) _07954_;
  assign _04992_ = _04991_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *) _08082_;
  assign in_wt_nan[56] = _04992_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *) in_wt_mask[112];
  assign _04993_ = { _07497_, _07497_, _07497_, _07497_, _07497_, _07497_, _07497_, _07497_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25957" *) wt7_sd_data[519:512];
  assign _04994_ = cfg_is_fp16_d1[55] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *) _07955_;
  assign _04995_ = _04994_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *) _08083_;
  assign in_wt_nan[55] = _04995_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *) in_wt_mask[110];
  assign _04996_ = { _07498_, _07498_, _07498_, _07498_, _07498_, _07498_, _07498_, _07498_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25967" *) wt7_sd_data[527:520];
  assign _04997_ = cfg_is_fp16_d1[54] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *) _07956_;
  assign _04998_ = _04997_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *) _08084_;
  assign in_wt_nan[54] = _04998_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *) in_wt_mask[108];
  assign _04999_ = { _07499_, _07499_, _07499_, _07499_, _07499_, _07499_, _07499_, _07499_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25977" *) wt7_sd_data[535:528];
  assign _05000_ = cfg_is_fp16_d1[53] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *) _07957_;
  assign _05001_ = _05000_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *) _08085_;
  assign in_wt_nan[53] = _05001_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *) in_wt_mask[106];
  assign _05002_ = { _07500_, _07500_, _07500_, _07500_, _07500_, _07500_, _07500_, _07500_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25987" *) wt7_sd_data[543:536];
  assign _05003_ = cfg_is_fp16_d1[52] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *) _07958_;
  assign _05004_ = _05003_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *) _08086_;
  assign in_wt_nan[52] = _05004_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *) in_wt_mask[104];
  assign _05005_ = { _07501_, _07501_, _07501_, _07501_, _07501_, _07501_, _07501_, _07501_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25997" *) wt7_sd_data[551:544];
  assign _05006_ = cfg_is_fp16_d1[51] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *) _07959_;
  assign _05007_ = _05006_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *) _08087_;
  assign in_wt_nan[51] = _05007_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *) in_wt_mask[102];
  assign _05008_ = { _07502_, _07502_, _07502_, _07502_, _07502_, _07502_, _07502_, _07502_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26007" *) wt7_sd_data[559:552];
  assign _05009_ = cfg_is_fp16_d1[50] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *) _07960_;
  assign _05010_ = _05009_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *) _08088_;
  assign in_wt_nan[50] = _05010_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *) in_wt_mask[100];
  assign _05011_ = { _07503_, _07503_, _07503_, _07503_, _07503_, _07503_, _07503_, _07503_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26017" *) wt7_sd_data[567:560];
  assign _05012_ = cfg_is_fp16_d1[49] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *) _07961_;
  assign _05013_ = _05012_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *) _08089_;
  assign in_wt_nan[49] = _05013_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *) in_wt_mask[98];
  assign _05014_ = { _07504_, _07504_, _07504_, _07504_, _07504_, _07504_, _07504_, _07504_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26027" *) wt7_sd_data[575:568];
  assign _05015_ = cfg_is_fp16_d1[48] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *) _07962_;
  assign _05016_ = _05015_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *) _08090_;
  assign in_wt_nan[48] = _05016_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *) in_wt_mask[96];
  assign _05017_ = { _07505_, _07505_, _07505_, _07505_, _07505_, _07505_, _07505_, _07505_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26037" *) wt7_sd_data[583:576];
  assign _05018_ = cfg_is_fp16_d1[47] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *) _07963_;
  assign _05019_ = _05018_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *) _08091_;
  assign in_wt_nan[47] = _05019_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *) in_wt_mask[94];
  assign _05020_ = { _07506_, _07506_, _07506_, _07506_, _07506_, _07506_, _07506_, _07506_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26047" *) wt7_sd_data[591:584];
  assign _05021_ = cfg_is_fp16_d1[46] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *) _07964_;
  assign _05022_ = _05021_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *) _08092_;
  assign in_wt_nan[46] = _05022_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *) in_wt_mask[92];
  assign _05023_ = { _07507_, _07507_, _07507_, _07507_, _07507_, _07507_, _07507_, _07507_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26057" *) wt7_sd_data[599:592];
  assign _05024_ = cfg_is_fp16_d1[45] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *) _07965_;
  assign _05025_ = _05024_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *) _08093_;
  assign in_wt_nan[45] = _05025_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *) in_wt_mask[90];
  assign _05026_ = { _07508_, _07508_, _07508_, _07508_, _07508_, _07508_, _07508_, _07508_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26067" *) wt7_sd_data[607:600];
  assign _05027_ = cfg_is_fp16_d1[44] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *) _07966_;
  assign _05028_ = _05027_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *) _08094_;
  assign in_wt_nan[44] = _05028_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *) in_wt_mask[88];
  assign _05029_ = { _07509_, _07509_, _07509_, _07509_, _07509_, _07509_, _07509_, _07509_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26077" *) wt7_sd_data[615:608];
  assign _05030_ = cfg_is_fp16_d1[43] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *) _07967_;
  assign _05031_ = _05030_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *) _08095_;
  assign in_wt_nan[43] = _05031_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *) in_wt_mask[86];
  assign _05032_ = { _07510_, _07510_, _07510_, _07510_, _07510_, _07510_, _07510_, _07510_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26087" *) wt7_sd_data[623:616];
  assign _05033_ = cfg_is_fp16_d1[42] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *) _07968_;
  assign _05034_ = _05033_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *) _08096_;
  assign in_wt_nan[42] = _05034_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *) in_wt_mask[84];
  assign _05035_ = { _07511_, _07511_, _07511_, _07511_, _07511_, _07511_, _07511_, _07511_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26097" *) wt7_sd_data[631:624];
  assign _05036_ = cfg_is_fp16_d1[41] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *) _07969_;
  assign _05037_ = _05036_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *) _08097_;
  assign in_wt_nan[41] = _05037_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *) in_wt_mask[82];
  assign _05038_ = { _07512_, _07512_, _07512_, _07512_, _07512_, _07512_, _07512_, _07512_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26107" *) wt7_sd_data[639:632];
  assign _05039_ = cfg_is_fp16_d1[40] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *) _07970_;
  assign _05040_ = _05039_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *) _08098_;
  assign in_wt_nan[40] = _05040_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *) in_wt_mask[80];
  assign _05041_ = { _07513_, _07513_, _07513_, _07513_, _07513_, _07513_, _07513_, _07513_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26117" *) wt7_sd_data[647:640];
  assign _05042_ = cfg_is_fp16_d1[39] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *) _07971_;
  assign _05043_ = _05042_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *) _08099_;
  assign in_wt_nan[39] = _05043_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *) in_wt_mask[78];
  assign _05044_ = { _07514_, _07514_, _07514_, _07514_, _07514_, _07514_, _07514_, _07514_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26127" *) wt7_sd_data[655:648];
  assign _05045_ = cfg_is_fp16_d1[38] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *) _07972_;
  assign _05046_ = _05045_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *) _08100_;
  assign in_wt_nan[38] = _05046_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *) in_wt_mask[76];
  assign _05047_ = { _07515_, _07515_, _07515_, _07515_, _07515_, _07515_, _07515_, _07515_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26137" *) wt7_sd_data[663:656];
  assign _05048_ = cfg_is_fp16_d1[37] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *) _07973_;
  assign _05049_ = _05048_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *) _08101_;
  assign in_wt_nan[37] = _05049_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *) in_wt_mask[74];
  assign _05050_ = { _07516_, _07516_, _07516_, _07516_, _07516_, _07516_, _07516_, _07516_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26147" *) wt7_sd_data[671:664];
  assign _05051_ = cfg_is_fp16_d1[36] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *) _07974_;
  assign _05052_ = _05051_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *) _08102_;
  assign in_wt_nan[36] = _05052_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *) in_wt_mask[72];
  assign _05053_ = { _07517_, _07517_, _07517_, _07517_, _07517_, _07517_, _07517_, _07517_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26157" *) wt7_sd_data[679:672];
  assign _05054_ = cfg_is_fp16_d1[35] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *) _07975_;
  assign _05055_ = _05054_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *) _08103_;
  assign in_wt_nan[35] = _05055_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *) in_wt_mask[70];
  assign _05056_ = { _07518_, _07518_, _07518_, _07518_, _07518_, _07518_, _07518_, _07518_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26167" *) wt7_sd_data[687:680];
  assign _05057_ = cfg_is_fp16_d1[34] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *) _07976_;
  assign _05058_ = _05057_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *) _08104_;
  assign in_wt_nan[34] = _05058_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *) in_wt_mask[68];
  assign _05059_ = { _07519_, _07519_, _07519_, _07519_, _07519_, _07519_, _07519_, _07519_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26177" *) wt7_sd_data[695:688];
  assign _05060_ = cfg_is_fp16_d1[33] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *) _07977_;
  assign _05061_ = _05060_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *) _08105_;
  assign in_wt_nan[33] = _05061_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *) in_wt_mask[66];
  assign _05062_ = { _07520_, _07520_, _07520_, _07520_, _07520_, _07520_, _07520_, _07520_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26187" *) wt7_sd_data[703:696];
  assign _05063_ = cfg_is_fp16_d1[32] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *) _07978_;
  assign _05064_ = _05063_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *) _08106_;
  assign in_wt_nan[32] = _05064_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *) in_wt_mask[64];
  assign _05065_ = { _07521_, _07521_, _07521_, _07521_, _07521_, _07521_, _07521_, _07521_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26197" *) wt7_sd_data[711:704];
  assign _05066_ = cfg_is_fp16_d1[31] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *) _07979_;
  assign _05067_ = _05066_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *) _08107_;
  assign in_wt_nan[31] = _05067_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *) in_wt_mask[62];
  assign _05068_ = { _07522_, _07522_, _07522_, _07522_, _07522_, _07522_, _07522_, _07522_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26207" *) wt7_sd_data[719:712];
  assign _05069_ = cfg_is_fp16_d1[30] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *) _07980_;
  assign _05070_ = _05069_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *) _08108_;
  assign in_wt_nan[30] = _05070_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *) in_wt_mask[60];
  assign _05071_ = { _07523_, _07523_, _07523_, _07523_, _07523_, _07523_, _07523_, _07523_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26217" *) wt7_sd_data[727:720];
  assign _05072_ = cfg_is_fp16_d1[29] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *) _07981_;
  assign _05073_ = _05072_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *) _08109_;
  assign in_wt_nan[29] = _05073_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *) in_wt_mask[58];
  assign _05074_ = { _07524_, _07524_, _07524_, _07524_, _07524_, _07524_, _07524_, _07524_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26227" *) wt7_sd_data[735:728];
  assign _05075_ = cfg_is_fp16_d1[28] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *) _07982_;
  assign _05076_ = _05075_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *) _08110_;
  assign in_wt_nan[28] = _05076_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *) in_wt_mask[56];
  assign _05077_ = { _07525_, _07525_, _07525_, _07525_, _07525_, _07525_, _07525_, _07525_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26237" *) wt7_sd_data[743:736];
  assign _05078_ = cfg_is_fp16_d1[27] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *) _07983_;
  assign _05079_ = _05078_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *) _08111_;
  assign in_wt_nan[27] = _05079_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *) in_wt_mask[54];
  assign _05080_ = { _07526_, _07526_, _07526_, _07526_, _07526_, _07526_, _07526_, _07526_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26247" *) wt7_sd_data[751:744];
  assign _05081_ = cfg_is_fp16_d1[26] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *) _07984_;
  assign _05082_ = _05081_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *) _08112_;
  assign in_wt_nan[26] = _05082_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *) in_wt_mask[52];
  assign _05083_ = { _07527_, _07527_, _07527_, _07527_, _07527_, _07527_, _07527_, _07527_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26257" *) wt7_sd_data[759:752];
  assign _05084_ = cfg_is_fp16_d1[25] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *) _07985_;
  assign _05085_ = _05084_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *) _08113_;
  assign in_wt_nan[25] = _05085_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *) in_wt_mask[50];
  assign _05086_ = { _07528_, _07528_, _07528_, _07528_, _07528_, _07528_, _07528_, _07528_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26267" *) wt7_sd_data[767:760];
  assign _05087_ = cfg_is_fp16_d1[24] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *) _07986_;
  assign _05088_ = _05087_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *) _08114_;
  assign in_wt_nan[24] = _05088_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *) in_wt_mask[48];
  assign _05089_ = { _07529_, _07529_, _07529_, _07529_, _07529_, _07529_, _07529_, _07529_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26277" *) wt7_sd_data[775:768];
  assign _05090_ = cfg_is_fp16_d1[23] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *) _07987_;
  assign _05091_ = _05090_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *) _08115_;
  assign in_wt_nan[23] = _05091_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *) in_wt_mask[46];
  assign _05092_ = { _07530_, _07530_, _07530_, _07530_, _07530_, _07530_, _07530_, _07530_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26287" *) wt7_sd_data[783:776];
  assign _05093_ = cfg_is_fp16_d1[22] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *) _07988_;
  assign _05094_ = _05093_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *) _08116_;
  assign in_wt_nan[22] = _05094_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *) in_wt_mask[44];
  assign _05095_ = { _07531_, _07531_, _07531_, _07531_, _07531_, _07531_, _07531_, _07531_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26297" *) wt7_sd_data[791:784];
  assign _05096_ = cfg_is_fp16_d1[21] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *) _07989_;
  assign _05097_ = _05096_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *) _08117_;
  assign in_wt_nan[21] = _05097_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *) in_wt_mask[42];
  assign _05098_ = { _07532_, _07532_, _07532_, _07532_, _07532_, _07532_, _07532_, _07532_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26307" *) wt7_sd_data[799:792];
  assign _05099_ = cfg_is_fp16_d1[20] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *) _07990_;
  assign _05100_ = _05099_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *) _08118_;
  assign in_wt_nan[20] = _05100_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *) in_wt_mask[40];
  assign _05101_ = { _07533_, _07533_, _07533_, _07533_, _07533_, _07533_, _07533_, _07533_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26317" *) wt7_sd_data[807:800];
  assign _05102_ = cfg_is_fp16_d1[19] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *) _07991_;
  assign _05103_ = _05102_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *) _08119_;
  assign in_wt_nan[19] = _05103_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *) in_wt_mask[38];
  assign _05104_ = { _07534_, _07534_, _07534_, _07534_, _07534_, _07534_, _07534_, _07534_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26327" *) wt7_sd_data[815:808];
  assign _05105_ = cfg_is_fp16_d1[18] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *) _07992_;
  assign _05106_ = _05105_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *) _08120_;
  assign in_wt_nan[18] = _05106_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *) in_wt_mask[36];
  assign _05107_ = { _07535_, _07535_, _07535_, _07535_, _07535_, _07535_, _07535_, _07535_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26337" *) wt7_sd_data[823:816];
  assign _05108_ = cfg_is_fp16_d1[17] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *) _07993_;
  assign _05109_ = _05108_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *) _08121_;
  assign in_wt_nan[17] = _05109_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *) in_wt_mask[34];
  assign _05110_ = { _07536_, _07536_, _07536_, _07536_, _07536_, _07536_, _07536_, _07536_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26347" *) wt7_sd_data[831:824];
  assign _05111_ = cfg_is_fp16_d1[16] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *) _07994_;
  assign _05112_ = _05111_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *) _08122_;
  assign in_wt_nan[16] = _05112_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *) in_wt_mask[32];
  assign _05113_ = { _07537_, _07537_, _07537_, _07537_, _07537_, _07537_, _07537_, _07537_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26357" *) wt7_sd_data[839:832];
  assign _05114_ = cfg_is_fp16_d1[15] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *) _07995_;
  assign _05115_ = _05114_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *) _08123_;
  assign in_wt_nan[15] = _05115_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *) in_wt_mask[30];
  assign _05116_ = { _07538_, _07538_, _07538_, _07538_, _07538_, _07538_, _07538_, _07538_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26367" *) wt7_sd_data[847:840];
  assign _05117_ = cfg_is_fp16_d1[14] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *) _07996_;
  assign _05118_ = _05117_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *) _08124_;
  assign in_wt_nan[14] = _05118_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *) in_wt_mask[28];
  assign _05119_ = { _07539_, _07539_, _07539_, _07539_, _07539_, _07539_, _07539_, _07539_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26377" *) wt7_sd_data[855:848];
  assign _05120_ = cfg_is_fp16_d1[13] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *) _07997_;
  assign _05121_ = _05120_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *) _08125_;
  assign in_wt_nan[13] = _05121_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *) in_wt_mask[26];
  assign _05122_ = { _07540_, _07540_, _07540_, _07540_, _07540_, _07540_, _07540_, _07540_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26387" *) wt7_sd_data[863:856];
  assign _05123_ = cfg_is_fp16_d1[12] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *) _07998_;
  assign _05124_ = _05123_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *) _08126_;
  assign in_wt_nan[12] = _05124_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *) in_wt_mask[24];
  assign _05125_ = { _07541_, _07541_, _07541_, _07541_, _07541_, _07541_, _07541_, _07541_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26397" *) wt7_sd_data[871:864];
  assign _05126_ = cfg_is_fp16_d1[11] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *) _07999_;
  assign _05127_ = _05126_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *) _08127_;
  assign in_wt_nan[11] = _05127_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *) in_wt_mask[22];
  assign _05128_ = { _07542_, _07542_, _07542_, _07542_, _07542_, _07542_, _07542_, _07542_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26407" *) wt7_sd_data[879:872];
  assign _05129_ = cfg_is_fp16_d1[10] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *) _08000_;
  assign _05130_ = _05129_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *) _08128_;
  assign in_wt_nan[10] = _05130_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *) in_wt_mask[20];
  assign _05131_ = { _07543_, _07543_, _07543_, _07543_, _07543_, _07543_, _07543_, _07543_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26417" *) wt7_sd_data[887:880];
  assign _05132_ = cfg_is_fp16_d1[9] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *) _08001_;
  assign _05133_ = _05132_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *) _08129_;
  assign in_wt_nan[9] = _05133_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *) in_wt_mask[18];
  assign _05134_ = { _07544_, _07544_, _07544_, _07544_, _07544_, _07544_, _07544_, _07544_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26427" *) wt7_sd_data[895:888];
  assign _05135_ = cfg_is_fp16_d1[8] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *) _08002_;
  assign _05136_ = _05135_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *) _08130_;
  assign in_wt_nan[8] = _05136_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *) in_wt_mask[16];
  assign _05137_ = { _07545_, _07545_, _07545_, _07545_, _07545_, _07545_, _07545_, _07545_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26437" *) wt7_sd_data[903:896];
  assign _05138_ = cfg_is_fp16_d1[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *) _08003_;
  assign _05139_ = _05138_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *) _08131_;
  assign in_wt_nan[7] = _05139_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *) in_wt_mask[14];
  assign _05140_ = { _07546_, _07546_, _07546_, _07546_, _07546_, _07546_, _07546_, _07546_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26447" *) wt7_sd_data[911:904];
  assign _05141_ = cfg_is_fp16_d1[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *) _08004_;
  assign _05142_ = _05141_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *) _08132_;
  assign in_wt_nan[6] = _05142_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *) in_wt_mask[12];
  assign _05143_ = { _07547_, _07547_, _07547_, _07547_, _07547_, _07547_, _07547_, _07547_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26457" *) wt7_sd_data[919:912];
  assign _05144_ = cfg_is_fp16_d1[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *) _08005_;
  assign _05145_ = _05144_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *) _08133_;
  assign in_wt_nan[5] = _05145_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *) in_wt_mask[10];
  assign _05146_ = { _07548_, _07548_, _07548_, _07548_, _07548_, _07548_, _07548_, _07548_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26467" *) wt7_sd_data[927:920];
  assign _05147_ = cfg_is_fp16_d1[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *) _08006_;
  assign _05148_ = _05147_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *) _08134_;
  assign in_wt_nan[4] = _05148_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *) in_wt_mask[8];
  assign _05149_ = { _07549_, _07549_, _07549_, _07549_, _07549_, _07549_, _07549_, _07549_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26477" *) wt7_sd_data[935:928];
  assign _05150_ = cfg_is_fp16_d1[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *) _08007_;
  assign _05151_ = _05150_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *) _08135_;
  assign in_wt_nan[3] = _05151_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *) in_wt_mask[6];
  assign _05152_ = { _07550_, _07550_, _07550_, _07550_, _07550_, _07550_, _07550_, _07550_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26487" *) wt7_sd_data[943:936];
  assign _05153_ = cfg_is_fp16_d1[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *) _08008_;
  assign _05154_ = _05153_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *) _08136_;
  assign in_wt_nan[2] = _05154_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *) in_wt_mask[4];
  assign _05155_ = { _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26497" *) wt7_sd_data[951:944];
  assign _05156_ = cfg_is_fp16_d1[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *) _08009_;
  assign _05157_ = _05156_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *) _08137_;
  assign in_wt_nan[1] = _05157_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *) in_wt_mask[2];
  assign _05158_ = { _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26507" *) wt7_sd_data[959:952];
  assign _05159_ = cfg_is_fp16_d1[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *) _08010_;
  assign _05160_ = _05159_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *) _08138_;
  assign in_wt_nan[0] = _05160_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *) in_wt_mask[0];
  assign _05161_ = { _07553_, _07553_, _07553_, _07553_, _07553_, _07553_, _07553_, _07553_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26517" *) wt7_sd_data[967:960];
  assign _05162_ = { _07554_, _07554_, _07554_, _07554_, _07554_, _07554_, _07554_, _07554_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26527" *) wt7_sd_data[975:968];
  assign _05163_ = { _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26537" *) wt7_sd_data[983:976];
  assign _05164_ = { _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26547" *) wt7_sd_data[991:984];
  assign _05165_ = { _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26557" *) wt7_sd_data[999:992];
  assign _05166_ = { _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26567" *) wt7_sd_data[1007:1000];
  assign _05167_ = { _07559_, _07559_, _07559_, _07559_, _07559_, _07559_, _07559_, _07559_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26577" *) wt7_sd_data[1015:1008];
  assign _05168_ = cfg_is_fp16_d1[63] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2658" *) in_wt_mask[127];
  assign wt_pre_exp_w[191:189] = { _05168_, _05168_, _05168_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2658" *) in_wt_data127[6:4];
  assign _05169_ = { _07560_, _07560_, _07560_, _07560_, _07560_, _07560_, _07560_, _07560_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26587" *) wt7_sd_data[1023:1016];
  assign _05170_ = cfg_is_fp16_d1[62] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2659" *) in_wt_mask[125];
  assign wt_pre_exp_w[188:186] = { _05170_, _05170_, _05170_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2659" *) in_wt_data125[6:4];
  assign _05171_ = cfg_is_fp16_d1[61] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2660" *) in_wt_mask[123];
  assign wt_pre_exp_w[185:183] = { _05171_, _05171_, _05171_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2660" *) in_wt_data123[6:4];
  assign _05172_ = cfg_is_fp16_d1[60] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2661" *) in_wt_mask[121];
  assign wt_pre_exp_w[182:180] = { _05172_, _05172_, _05172_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2661" *) in_wt_data121[6:4];
  assign _05173_ = cfg_is_fp16_d1[59] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2662" *) in_wt_mask[119];
  assign wt_pre_exp_w[179:177] = { _05173_, _05173_, _05173_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2662" *) in_wt_data119[6:4];
  assign _05174_ = cfg_is_fp16_d1[58] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2663" *) in_wt_mask[117];
  assign wt_pre_exp_w[176:174] = { _05174_, _05174_, _05174_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2663" *) in_wt_data117[6:4];
  assign _05175_ = cfg_is_fp16_d1[57] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2664" *) in_wt_mask[115];
  assign wt_pre_exp_w[173:171] = { _05175_, _05175_, _05175_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2664" *) in_wt_data115[6:4];
  assign _05176_ = cfg_is_fp16_d1[56] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2665" *) in_wt_mask[113];
  assign wt_pre_exp_w[170:168] = { _05176_, _05176_, _05176_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2665" *) in_wt_data113[6:4];
  assign _05177_ = cfg_is_fp16_d1[55] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2666" *) in_wt_mask[111];
  assign wt_pre_exp_w[167:165] = { _05177_, _05177_, _05177_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2666" *) in_wt_data111[6:4];
  assign _05178_ = cfg_is_fp16_d1[54] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2667" *) in_wt_mask[109];
  assign wt_pre_exp_w[164:162] = { _05178_, _05178_, _05178_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2667" *) in_wt_data109[6:4];
  assign _05179_ = cfg_is_fp16_d1[53] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2668" *) in_wt_mask[107];
  assign wt_pre_exp_w[161:159] = { _05179_, _05179_, _05179_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2668" *) in_wt_data107[6:4];
  assign _05180_ = cfg_is_fp16_d1[52] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2669" *) in_wt_mask[105];
  assign wt_pre_exp_w[158:156] = { _05180_, _05180_, _05180_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2669" *) in_wt_data105[6:4];
  assign _05181_ = cfg_is_fp16_d1[51] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2670" *) in_wt_mask[103];
  assign wt_pre_exp_w[155:153] = { _05181_, _05181_, _05181_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2670" *) in_wt_data103[6:4];
  assign _05182_ = cfg_is_fp16_d1[50] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2671" *) in_wt_mask[101];
  assign wt_pre_exp_w[152:150] = { _05182_, _05182_, _05182_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2671" *) in_wt_data101[6:4];
  assign _05183_ = cfg_is_fp16_d1[49] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2672" *) in_wt_mask[99];
  assign wt_pre_exp_w[149:147] = { _05183_, _05183_, _05183_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2672" *) in_wt_data99[6:4];
  assign _05184_ = cfg_is_fp16_d1[48] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2673" *) in_wt_mask[97];
  assign wt_pre_exp_w[146:144] = { _05184_, _05184_, _05184_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2673" *) in_wt_data97[6:4];
  assign _05185_ = cfg_is_fp16_d1[47] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2674" *) in_wt_mask[95];
  assign wt_pre_exp_w[143:141] = { _05185_, _05185_, _05185_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2674" *) in_wt_data95[6:4];
  assign _05186_ = cfg_is_fp16_d1[46] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2675" *) in_wt_mask[93];
  assign wt_pre_exp_w[140:138] = { _05186_, _05186_, _05186_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2675" *) in_wt_data93[6:4];
  assign _05187_ = cfg_is_fp16_d1[45] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2676" *) in_wt_mask[91];
  assign wt_pre_exp_w[137:135] = { _05187_, _05187_, _05187_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2676" *) in_wt_data91[6:4];
  assign _05188_ = cfg_is_fp16_d1[44] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2677" *) in_wt_mask[89];
  assign wt_pre_exp_w[134:132] = { _05188_, _05188_, _05188_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2677" *) in_wt_data89[6:4];
  assign _05189_ = cfg_is_fp16_d1[43] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2678" *) in_wt_mask[87];
  assign wt_pre_exp_w[131:129] = { _05189_, _05189_, _05189_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2678" *) in_wt_data87[6:4];
  assign _05190_ = cfg_is_fp16_d1[42] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2679" *) in_wt_mask[85];
  assign wt_pre_exp_w[128:126] = { _05190_, _05190_, _05190_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2679" *) in_wt_data85[6:4];
  assign _05191_ = cfg_is_fp16_d1[41] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2680" *) in_wt_mask[83];
  assign wt_pre_exp_w[125:123] = { _05191_, _05191_, _05191_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2680" *) in_wt_data83[6:4];
  assign _05192_ = cfg_is_fp16_d1[40] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2681" *) in_wt_mask[81];
  assign wt_pre_exp_w[122:120] = { _05192_, _05192_, _05192_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2681" *) in_wt_data81[6:4];
  assign _05193_ = cfg_is_fp16_d1[39] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2682" *) in_wt_mask[79];
  assign wt_pre_exp_w[119:117] = { _05193_, _05193_, _05193_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2682" *) in_wt_data79[6:4];
  assign _05194_ = cfg_is_fp16_d1[38] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2683" *) in_wt_mask[77];
  assign wt_pre_exp_w[116:114] = { _05194_, _05194_, _05194_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2683" *) in_wt_data77[6:4];
  assign _05195_ = cfg_is_fp16_d1[37] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2684" *) in_wt_mask[75];
  assign wt_pre_exp_w[113:111] = { _05195_, _05195_, _05195_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2684" *) in_wt_data75[6:4];
  assign _05196_ = cfg_is_fp16_d1[36] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2685" *) in_wt_mask[73];
  assign wt_pre_exp_w[110:108] = { _05196_, _05196_, _05196_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2685" *) in_wt_data73[6:4];
  assign _05197_ = cfg_is_fp16_d1[35] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2686" *) in_wt_mask[71];
  assign wt_pre_exp_w[107:105] = { _05197_, _05197_, _05197_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2686" *) in_wt_data71[6:4];
  assign _05198_ = cfg_is_fp16_d1[34] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2687" *) in_wt_mask[69];
  assign wt_pre_exp_w[104:102] = { _05198_, _05198_, _05198_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2687" *) in_wt_data69[6:4];
  assign _05199_ = cfg_is_fp16_d1[33] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2688" *) in_wt_mask[67];
  assign wt_pre_exp_w[101:99] = { _05199_, _05199_, _05199_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2688" *) in_wt_data67[6:4];
  assign _05200_ = cfg_is_fp16_d1[32] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2689" *) in_wt_mask[65];
  assign wt_pre_exp_w[98:96] = { _05200_, _05200_, _05200_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2689" *) in_wt_data65[6:4];
  assign _05201_ = cfg_is_fp16_d1[31] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2690" *) in_wt_mask[63];
  assign wt_pre_exp_w[95:93] = { _05201_, _05201_, _05201_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2690" *) in_wt_data63[6:4];
  assign _05202_ = cfg_is_fp16_d1[30] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2691" *) in_wt_mask[61];
  assign wt_pre_exp_w[92:90] = { _05202_, _05202_, _05202_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2691" *) in_wt_data61[6:4];
  assign _05203_ = cfg_is_fp16_d1[29] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2692" *) in_wt_mask[59];
  assign wt_pre_exp_w[89:87] = { _05203_, _05203_, _05203_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2692" *) in_wt_data59[6:4];
  assign _05204_ = cfg_is_fp16_d1[28] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2693" *) in_wt_mask[57];
  assign wt_pre_exp_w[86:84] = { _05204_, _05204_, _05204_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2693" *) in_wt_data57[6:4];
  assign _05205_ = cfg_is_fp16_d1[27] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2694" *) in_wt_mask[55];
  assign wt_pre_exp_w[83:81] = { _05205_, _05205_, _05205_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2694" *) in_wt_data55[6:4];
  assign _05206_ = cfg_is_fp16_d1[26] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2695" *) in_wt_mask[53];
  assign wt_pre_exp_w[80:78] = { _05206_, _05206_, _05206_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2695" *) in_wt_data53[6:4];
  assign _05207_ = cfg_is_fp16_d1[25] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2696" *) in_wt_mask[51];
  assign wt_pre_exp_w[77:75] = { _05207_, _05207_, _05207_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2696" *) in_wt_data51[6:4];
  assign _05208_ = cfg_is_fp16_d1[24] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2697" *) in_wt_mask[49];
  assign wt_pre_exp_w[74:72] = { _05208_, _05208_, _05208_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2697" *) in_wt_data49[6:4];
  assign _05209_ = cfg_is_fp16_d1[23] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2698" *) in_wt_mask[47];
  assign wt_pre_exp_w[71:69] = { _05209_, _05209_, _05209_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2698" *) in_wt_data47[6:4];
  assign _05210_ = cfg_is_fp16_d1[22] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2699" *) in_wt_mask[45];
  assign wt_pre_exp_w[68:66] = { _05210_, _05210_, _05210_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2699" *) in_wt_data45[6:4];
  assign _05211_ = cfg_is_fp16_d1[21] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2700" *) in_wt_mask[43];
  assign wt_pre_exp_w[65:63] = { _05211_, _05211_, _05211_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2700" *) in_wt_data43[6:4];
  assign _05212_ = cfg_is_fp16_d1[20] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2701" *) in_wt_mask[41];
  assign wt_pre_exp_w[62:60] = { _05212_, _05212_, _05212_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2701" *) in_wt_data41[6:4];
  assign _05213_ = cfg_is_fp16_d1[19] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2702" *) in_wt_mask[39];
  assign wt_pre_exp_w[59:57] = { _05213_, _05213_, _05213_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2702" *) in_wt_data39[6:4];
  assign _05214_ = cfg_is_fp16_d1[18] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2703" *) in_wt_mask[37];
  assign wt_pre_exp_w[56:54] = { _05214_, _05214_, _05214_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2703" *) in_wt_data37[6:4];
  assign _05215_ = cfg_is_fp16_d1[17] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2704" *) in_wt_mask[35];
  assign wt_pre_exp_w[53:51] = { _05215_, _05215_, _05215_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2704" *) in_wt_data35[6:4];
  assign _05216_ = cfg_is_fp16_d1[16] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2705" *) in_wt_mask[33];
  assign wt_pre_exp_w[50:48] = { _05216_, _05216_, _05216_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2705" *) in_wt_data33[6:4];
  assign _05217_ = cfg_is_fp16_d1[15] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2706" *) in_wt_mask[31];
  assign wt_pre_exp_w[47:45] = { _05217_, _05217_, _05217_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2706" *) in_wt_data31[6:4];
  assign _05218_ = cfg_is_fp16_d1[14] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2707" *) in_wt_mask[29];
  assign wt_pre_exp_w[44:42] = { _05218_, _05218_, _05218_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2707" *) in_wt_data29[6:4];
  assign _05219_ = cfg_is_fp16_d1[13] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2708" *) in_wt_mask[27];
  assign wt_pre_exp_w[41:39] = { _05219_, _05219_, _05219_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2708" *) in_wt_data27[6:4];
  assign _05220_ = cfg_is_fp16_d1[12] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2709" *) in_wt_mask[25];
  assign wt_pre_exp_w[38:36] = { _05220_, _05220_, _05220_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2709" *) in_wt_data25[6:4];
  assign _05221_ = cfg_is_fp16_d1[11] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2710" *) in_wt_mask[23];
  assign wt_pre_exp_w[35:33] = { _05221_, _05221_, _05221_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2710" *) in_wt_data23[6:4];
  assign _05222_ = cfg_is_fp16_d1[10] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2711" *) in_wt_mask[21];
  assign wt_pre_exp_w[32:30] = { _05222_, _05222_, _05222_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2711" *) in_wt_data21[6:4];
  assign _05223_ = cfg_is_fp16_d1[9] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2712" *) in_wt_mask[19];
  assign wt_pre_exp_w[29:27] = { _05223_, _05223_, _05223_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2712" *) in_wt_data19[6:4];
  assign _05224_ = cfg_is_fp16_d1[8] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2713" *) in_wt_mask[17];
  assign wt_pre_exp_w[26:24] = { _05224_, _05224_, _05224_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2713" *) in_wt_data17[6:4];
  assign _05225_ = cfg_is_fp16_d1[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2714" *) in_wt_mask[15];
  assign wt_pre_exp_w[23:21] = { _05225_, _05225_, _05225_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2714" *) in_wt_data15[6:4];
  assign _05226_ = cfg_is_fp16_d1[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2715" *) in_wt_mask[13];
  assign wt_pre_exp_w[20:18] = { _05226_, _05226_, _05226_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2715" *) in_wt_data13[6:4];
  assign _05227_ = cfg_is_fp16_d1[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2716" *) in_wt_mask[11];
  assign wt_pre_exp_w[17:15] = { _05227_, _05227_, _05227_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2716" *) in_wt_data11[6:4];
  assign _05228_ = cfg_is_fp16_d1[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2717" *) in_wt_mask[9];
  assign wt_pre_exp_w[14:12] = { _05228_, _05228_, _05228_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2717" *) in_wt_data9[6:4];
  assign _05229_ = cfg_is_fp16_d1[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2718" *) in_wt_mask[7];
  assign wt_pre_exp_w[11:9] = { _05229_, _05229_, _05229_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2718" *) in_wt_data7[6:4];
  assign _05230_ = cfg_is_fp16_d1[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2719" *) in_wt_mask[5];
  assign wt_pre_exp_w[8:6] = { _05230_, _05230_, _05230_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2719" *) in_wt_data5[6:4];
  assign _05231_ = cfg_is_fp16_d1[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2720" *) in_wt_mask[3];
  assign wt_pre_exp_w[5:3] = { _05231_, _05231_, _05231_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2720" *) in_wt_data3[6:4];
  assign _05232_ = cfg_is_fp16_d1[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2721" *) in_wt_mask[1];
  assign wt_pre_exp_w[2:0] = { _05232_, _05232_, _05232_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2721" *) in_wt_data1[6:4];
  assign in_dat_data_int16_63 = { cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63], cfg_is_int16_d1[63] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27245" *) { in_dat_data127, in_dat_data126 };
  assign in_dat_data_int16_62 = { cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62], cfg_is_int16_d1[62] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27246" *) { in_dat_data125, in_dat_data124 };
  assign in_dat_data_int16_61 = { cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61], cfg_is_int16_d1[61] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27247" *) { in_dat_data123, in_dat_data122 };
  assign in_dat_data_int16_60 = { cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60], cfg_is_int16_d1[60] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27248" *) { in_dat_data121, in_dat_data120 };
  assign in_dat_data_int16_59 = { cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59], cfg_is_int16_d1[59] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27249" *) { in_dat_data119, in_dat_data118 };
  assign in_dat_data_int16_58 = { cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58], cfg_is_int16_d1[58] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27250" *) { in_dat_data117, in_dat_data116 };
  assign in_dat_data_int16_57 = { cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57], cfg_is_int16_d1[57] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27251" *) { in_dat_data115, in_dat_data114 };
  assign in_dat_data_int16_56 = { cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56], cfg_is_int16_d1[56] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27252" *) { in_dat_data113, in_dat_data112 };
  assign in_dat_data_int16_55 = { cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55], cfg_is_int16_d1[55] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27253" *) { in_dat_data111, in_dat_data110 };
  assign in_dat_data_int16_54 = { cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54], cfg_is_int16_d1[54] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27254" *) { in_dat_data109, in_dat_data108 };
  assign in_dat_data_int16_53 = { cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53], cfg_is_int16_d1[53] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27255" *) { in_dat_data107, in_dat_data106 };
  assign in_dat_data_int16_52 = { cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52], cfg_is_int16_d1[52] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27256" *) { in_dat_data105, in_dat_data104 };
  assign in_dat_data_int16_51 = { cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51], cfg_is_int16_d1[51] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27257" *) { in_dat_data103, in_dat_data102 };
  assign in_dat_data_int16_50 = { cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50], cfg_is_int16_d1[50] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27258" *) { in_dat_data101, in_dat_data100 };
  assign in_dat_data_int16_49 = { cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49], cfg_is_int16_d1[49] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27259" *) { in_dat_data99, in_dat_data98 };
  assign in_dat_data_int16_48 = { cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48], cfg_is_int16_d1[48] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27260" *) { in_dat_data97, in_dat_data96 };
  assign in_dat_data_int16_47 = { cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47], cfg_is_int16_d1[47] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27261" *) { in_dat_data95, in_dat_data94 };
  assign in_dat_data_int16_46 = { cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46], cfg_is_int16_d1[46] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27262" *) { in_dat_data93, in_dat_data92 };
  assign in_dat_data_int16_45 = { cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45], cfg_is_int16_d1[45] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27263" *) { in_dat_data91, in_dat_data90 };
  assign in_dat_data_int16_44 = { cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44], cfg_is_int16_d1[44] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27264" *) { in_dat_data89, in_dat_data88 };
  assign in_dat_data_int16_43 = { cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43], cfg_is_int16_d1[43] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27265" *) { in_dat_data87, in_dat_data86 };
  assign in_dat_data_int16_42 = { cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42], cfg_is_int16_d1[42] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27266" *) { in_dat_data85, in_dat_data84 };
  assign in_dat_data_int16_41 = { cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41], cfg_is_int16_d1[41] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27267" *) { in_dat_data83, in_dat_data82 };
  assign in_dat_data_int16_40 = { cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40], cfg_is_int16_d1[40] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27268" *) { in_dat_data81, in_dat_data80 };
  assign in_dat_data_int16_39 = { cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39], cfg_is_int16_d1[39] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27269" *) { in_dat_data79, in_dat_data78 };
  assign in_wt_norm[63] = cfg_is_fp16_d1[63] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2727" *) _08139_;
  assign in_dat_data_int16_38 = { cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38], cfg_is_int16_d1[38] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27270" *) { in_dat_data77, in_dat_data76 };
  assign in_dat_data_int16_37 = { cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37], cfg_is_int16_d1[37] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27271" *) { in_dat_data75, in_dat_data74 };
  assign in_dat_data_int16_36 = { cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36], cfg_is_int16_d1[36] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27272" *) { in_dat_data73, in_dat_data72 };
  assign in_dat_data_int16_35 = { cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35], cfg_is_int16_d1[35] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27273" *) { in_dat_data71, in_dat_data70 };
  assign in_dat_data_int16_34 = { cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34], cfg_is_int16_d1[34] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27274" *) { in_dat_data69, in_dat_data68 };
  assign in_dat_data_int16_33 = { cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33], cfg_is_int16_d1[33] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27275" *) { in_dat_data67, in_dat_data66 };
  assign in_dat_data_int16_32 = { cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32], cfg_is_int16_d1[32] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27276" *) { in_dat_data65, in_dat_data64 };
  assign in_dat_data_int16_31 = { cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31], cfg_is_int16_d1[31] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27277" *) { in_dat_data63, in_dat_data62 };
  assign in_dat_data_int16_30 = { cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30], cfg_is_int16_d1[30] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27278" *) { in_dat_data61, in_dat_data60 };
  assign in_dat_data_int16_29 = { cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29], cfg_is_int16_d1[29] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27279" *) { in_dat_data59, in_dat_data58 };
  assign in_wt_norm[62] = cfg_is_fp16_d1[62] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2728" *) _08140_;
  assign in_dat_data_int16_28 = { cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28], cfg_is_int16_d1[28] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27280" *) { in_dat_data57, in_dat_data56 };
  assign in_dat_data_int16_27 = { cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27], cfg_is_int16_d1[27] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27281" *) { in_dat_data55, in_dat_data54 };
  assign in_dat_data_int16_26 = { cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26], cfg_is_int16_d1[26] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27282" *) { in_dat_data53, in_dat_data52 };
  assign in_dat_data_int16_25 = { cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25], cfg_is_int16_d1[25] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27283" *) { in_dat_data51, in_dat_data50 };
  assign in_dat_data_int16_24 = { cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24], cfg_is_int16_d1[24] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27284" *) { in_dat_data49, in_dat_data48 };
  assign in_dat_data_int16_23 = { cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23], cfg_is_int16_d1[23] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27285" *) { in_dat_data47, in_dat_data46 };
  assign in_dat_data_int16_22 = { cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22], cfg_is_int16_d1[22] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27286" *) { in_dat_data45, in_dat_data44 };
  assign in_dat_data_int16_21 = { cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21], cfg_is_int16_d1[21] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27287" *) { in_dat_data43, in_dat_data42 };
  assign in_dat_data_int16_20 = { cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20], cfg_is_int16_d1[20] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27288" *) { in_dat_data41, in_dat_data40 };
  assign in_dat_data_int16_19 = { cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19], cfg_is_int16_d1[19] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27289" *) { in_dat_data39, in_dat_data38 };
  assign in_wt_norm[61] = cfg_is_fp16_d1[61] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2729" *) _08141_;
  assign in_dat_data_int16_18 = { cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18], cfg_is_int16_d1[18] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27290" *) { in_dat_data37, in_dat_data36 };
  assign in_dat_data_int16_17 = { cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17], cfg_is_int16_d1[17] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27291" *) { in_dat_data35, in_dat_data34 };
  assign in_dat_data_int16_16 = { cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16], cfg_is_int16_d1[16] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27292" *) { in_dat_data33, in_dat_data32 };
  assign in_dat_data_int16_15 = { cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15], cfg_is_int16_d1[15] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27293" *) { in_dat_data31, in_dat_data30 };
  assign in_dat_data_int16_14 = { cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14], cfg_is_int16_d1[14] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27294" *) { in_dat_data29, in_dat_data28 };
  assign in_dat_data_int16_13 = { cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13], cfg_is_int16_d1[13] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27295" *) { in_dat_data27, in_dat_data26 };
  assign in_dat_data_int16_12 = { cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12], cfg_is_int16_d1[12] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27296" *) { in_dat_data25, in_dat_data24 };
  assign in_dat_data_int16_11 = { cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11], cfg_is_int16_d1[11] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27297" *) { in_dat_data23, in_dat_data22 };
  assign in_dat_data_int16_10 = { cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10], cfg_is_int16_d1[10] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27298" *) { in_dat_data21, in_dat_data20 };
  assign in_dat_data_int16_9 = { cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9], cfg_is_int16_d1[9] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27299" *) { in_dat_data19, in_dat_data18 };
  assign in_wt_norm[60] = cfg_is_fp16_d1[60] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2730" *) _08142_;
  assign in_dat_data_int16_8 = { cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8], cfg_is_int16_d1[8] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27300" *) { in_dat_data17, in_dat_data16 };
  assign in_dat_data_int16_7 = { cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7], cfg_is_int16_d1[7] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27301" *) { in_dat_data15, in_dat_data14 };
  assign in_dat_data_int16_6 = { cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6], cfg_is_int16_d1[6] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27302" *) { in_dat_data13, in_dat_data12 };
  assign in_dat_data_int16_5 = { cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5], cfg_is_int16_d1[5] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27303" *) { in_dat_data11, in_dat_data10 };
  assign in_dat_data_int16_4 = { cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4], cfg_is_int16_d1[4] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27304" *) { in_dat_data9, in_dat_data8 };
  assign in_dat_data_int16_3 = { cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3], cfg_is_int16_d1[3] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27305" *) { in_dat_data7, in_dat_data6 };
  assign in_dat_data_int16_2 = { cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2], cfg_is_int16_d1[2] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27306" *) { in_dat_data5, in_dat_data4 };
  assign in_dat_data_int16_1 = { cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1], cfg_is_int16_d1[1] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27307" *) { in_dat_data3, in_dat_data2 };
  assign in_dat_data_int16_0 = { cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0], cfg_is_int16_d1[0] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27308" *) { in_dat_data1, in_dat_data0 };
  assign in_wt_norm[59] = cfg_is_fp16_d1[59] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2731" *) _08143_;
  assign in_wt_norm[58] = cfg_is_fp16_d1[58] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2732" *) _08144_;
  assign in_wt_norm[57] = cfg_is_fp16_d1[57] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2733" *) _08145_;
  assign in_wt_norm[56] = cfg_is_fp16_d1[56] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2734" *) _08146_;
  assign in_wt_norm[55] = cfg_is_fp16_d1[55] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2735" *) _08147_;
  assign in_wt_norm[54] = cfg_is_fp16_d1[54] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2736" *) _08148_;
  assign in_wt_norm[53] = cfg_is_fp16_d1[53] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2737" *) _08149_;
  assign in_wt_norm[52] = cfg_is_fp16_d1[52] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2738" *) _08150_;
  assign in_wt_norm[51] = cfg_is_fp16_d1[51] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2739" *) _08151_;
  assign in_wt_norm[50] = cfg_is_fp16_d1[50] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2740" *) _08152_;
  assign in_wt_norm[49] = cfg_is_fp16_d1[49] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2741" *) _08153_;
  assign in_wt_norm[48] = cfg_is_fp16_d1[48] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2742" *) _08154_;
  assign in_wt_norm[47] = cfg_is_fp16_d1[47] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2743" *) _08155_;
  assign in_wt_norm[46] = cfg_is_fp16_d1[46] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2744" *) _08156_;
  assign in_wt_norm[45] = cfg_is_fp16_d1[45] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2745" *) _08157_;
  assign in_wt_norm[44] = cfg_is_fp16_d1[44] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2746" *) _08158_;
  assign in_wt_norm[43] = cfg_is_fp16_d1[43] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2747" *) _08159_;
  assign in_wt_norm[42] = cfg_is_fp16_d1[42] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2748" *) _08160_;
  assign in_wt_norm[41] = cfg_is_fp16_d1[41] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2749" *) _08161_;
  assign in_wt_norm[40] = cfg_is_fp16_d1[40] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2750" *) _08162_;
  assign in_wt_norm[39] = cfg_is_fp16_d1[39] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2751" *) _08163_;
  assign in_dat_data_int8_63 = { cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63], cfg_is_int8_d1[63] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27510" *) { in_dat_data127, in_dat_data63 };
  assign in_dat_data_int8_62 = { cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62], cfg_is_int8_d1[62] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27511" *) { in_dat_data126, in_dat_data62 };
  assign in_dat_data_int8_61 = { cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61], cfg_is_int8_d1[61] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27512" *) { in_dat_data125, in_dat_data61 };
  assign in_dat_data_int8_60 = { cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60], cfg_is_int8_d1[60] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27513" *) { in_dat_data124, in_dat_data60 };
  assign in_dat_data_int8_59 = { cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59], cfg_is_int8_d1[59] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27514" *) { in_dat_data123, in_dat_data59 };
  assign in_dat_data_int8_58 = { cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58], cfg_is_int8_d1[58] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27515" *) { in_dat_data122, in_dat_data58 };
  assign in_dat_data_int8_57 = { cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57], cfg_is_int8_d1[57] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27516" *) { in_dat_data121, in_dat_data57 };
  assign in_dat_data_int8_56 = { cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56], cfg_is_int8_d1[56] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27517" *) { in_dat_data120, in_dat_data56 };
  assign in_dat_data_int8_55 = { cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55], cfg_is_int8_d1[55] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27518" *) { in_dat_data119, in_dat_data55 };
  assign in_dat_data_int8_54 = { cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54], cfg_is_int8_d1[54] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27519" *) { in_dat_data118, in_dat_data54 };
  assign in_wt_norm[38] = cfg_is_fp16_d1[38] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2752" *) _08164_;
  assign in_dat_data_int8_53 = { cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53], cfg_is_int8_d1[53] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27520" *) { in_dat_data117, in_dat_data53 };
  assign in_dat_data_int8_52 = { cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52], cfg_is_int8_d1[52] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27521" *) { in_dat_data116, in_dat_data52 };
  assign in_dat_data_int8_51 = { cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51], cfg_is_int8_d1[51] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27522" *) { in_dat_data115, in_dat_data51 };
  assign in_dat_data_int8_50 = { cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50], cfg_is_int8_d1[50] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27523" *) { in_dat_data114, in_dat_data50 };
  assign in_dat_data_int8_49 = { cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49], cfg_is_int8_d1[49] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27524" *) { in_dat_data113, in_dat_data49 };
  assign in_dat_data_int8_48 = { cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48], cfg_is_int8_d1[48] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27525" *) { in_dat_data112, in_dat_data48 };
  assign in_dat_data_int8_47 = { cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47], cfg_is_int8_d1[47] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27526" *) { in_dat_data111, in_dat_data47 };
  assign in_dat_data_int8_46 = { cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46], cfg_is_int8_d1[46] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27527" *) { in_dat_data110, in_dat_data46 };
  assign in_dat_data_int8_45 = { cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45], cfg_is_int8_d1[45] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27528" *) { in_dat_data109, in_dat_data45 };
  assign in_dat_data_int8_44 = { cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44], cfg_is_int8_d1[44] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27529" *) { in_dat_data108, in_dat_data44 };
  assign in_wt_norm[37] = cfg_is_fp16_d1[37] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2753" *) _08165_;
  assign in_dat_data_int8_43 = { cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43], cfg_is_int8_d1[43] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27530" *) { in_dat_data107, in_dat_data43 };
  assign in_dat_data_int8_42 = { cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42], cfg_is_int8_d1[42] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27531" *) { in_dat_data106, in_dat_data42 };
  assign in_dat_data_int8_41 = { cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41], cfg_is_int8_d1[41] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27532" *) { in_dat_data105, in_dat_data41 };
  assign in_dat_data_int8_40 = { cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40], cfg_is_int8_d1[40] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27533" *) { in_dat_data104, in_dat_data40 };
  assign in_dat_data_int8_39 = { cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39], cfg_is_int8_d1[39] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27534" *) { in_dat_data103, in_dat_data39 };
  assign in_dat_data_int8_38 = { cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38], cfg_is_int8_d1[38] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27535" *) { in_dat_data102, in_dat_data38 };
  assign in_dat_data_int8_37 = { cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37], cfg_is_int8_d1[37] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27536" *) { in_dat_data101, in_dat_data37 };
  assign in_dat_data_int8_36 = { cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36], cfg_is_int8_d1[36] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27537" *) { in_dat_data100, in_dat_data36 };
  assign in_dat_data_int8_35 = { cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35], cfg_is_int8_d1[35] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27538" *) { in_dat_data99, in_dat_data35 };
  assign in_dat_data_int8_34 = { cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34], cfg_is_int8_d1[34] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27539" *) { in_dat_data98, in_dat_data34 };
  assign in_wt_norm[36] = cfg_is_fp16_d1[36] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2754" *) _08166_;
  assign in_dat_data_int8_33 = { cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33], cfg_is_int8_d1[33] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27540" *) { in_dat_data97, in_dat_data33 };
  assign in_dat_data_int8_32 = { cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32], cfg_is_int8_d1[32] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27541" *) { in_dat_data96, in_dat_data32 };
  assign in_dat_data_int8_31 = { cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31], cfg_is_int8_d1[31] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27542" *) { in_dat_data95, in_dat_data31 };
  assign in_dat_data_int8_30 = { cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30], cfg_is_int8_d1[30] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27543" *) { in_dat_data94, in_dat_data30 };
  assign in_dat_data_int8_29 = { cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29], cfg_is_int8_d1[29] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27544" *) { in_dat_data93, in_dat_data29 };
  assign in_dat_data_int8_28 = { cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28], cfg_is_int8_d1[28] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27545" *) { in_dat_data92, in_dat_data28 };
  assign in_dat_data_int8_27 = { cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27], cfg_is_int8_d1[27] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27546" *) { in_dat_data91, in_dat_data27 };
  assign in_dat_data_int8_26 = { cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26], cfg_is_int8_d1[26] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27547" *) { in_dat_data90, in_dat_data26 };
  assign in_dat_data_int8_25 = { cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25], cfg_is_int8_d1[25] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27548" *) { in_dat_data89, in_dat_data25 };
  assign in_dat_data_int8_24 = { cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24], cfg_is_int8_d1[24] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27549" *) { in_dat_data88, in_dat_data24 };
  assign in_wt_norm[35] = cfg_is_fp16_d1[35] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2755" *) _08167_;
  assign in_dat_data_int8_23 = { cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23], cfg_is_int8_d1[23] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27550" *) { in_dat_data87, in_dat_data23 };
  assign in_dat_data_int8_22 = { cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22], cfg_is_int8_d1[22] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27551" *) { in_dat_data86, in_dat_data22 };
  assign in_dat_data_int8_21 = { cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21], cfg_is_int8_d1[21] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27552" *) { in_dat_data85, in_dat_data21 };
  assign in_dat_data_int8_20 = { cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20], cfg_is_int8_d1[20] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27553" *) { in_dat_data84, in_dat_data20 };
  assign in_dat_data_int8_19 = { cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19], cfg_is_int8_d1[19] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27554" *) { in_dat_data83, in_dat_data19 };
  assign in_dat_data_int8_18 = { cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18], cfg_is_int8_d1[18] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27555" *) { in_dat_data82, in_dat_data18 };
  assign in_dat_data_int8_17 = { cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17], cfg_is_int8_d1[17] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27556" *) { in_dat_data81, in_dat_data17 };
  assign in_dat_data_int8_16 = { cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16], cfg_is_int8_d1[16] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27557" *) { in_dat_data80, in_dat_data16 };
  assign in_dat_data_int8_15 = { cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15], cfg_is_int8_d1[15] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27558" *) { in_dat_data79, in_dat_data15 };
  assign in_dat_data_int8_14 = { cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14], cfg_is_int8_d1[14] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27559" *) { in_dat_data78, in_dat_data14 };
  assign in_wt_norm[34] = cfg_is_fp16_d1[34] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2756" *) _08168_;
  assign in_dat_data_int8_13 = { cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13], cfg_is_int8_d1[13] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27560" *) { in_dat_data77, in_dat_data13 };
  assign in_dat_data_int8_12 = { cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12], cfg_is_int8_d1[12] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27561" *) { in_dat_data76, in_dat_data12 };
  assign in_dat_data_int8_11 = { cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11], cfg_is_int8_d1[11] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27562" *) { in_dat_data75, in_dat_data11 };
  assign in_dat_data_int8_10 = { cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10], cfg_is_int8_d1[10] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27563" *) { in_dat_data74, in_dat_data10 };
  assign in_dat_data_int8_9 = { cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9], cfg_is_int8_d1[9] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27564" *) { in_dat_data73, in_dat_data9 };
  assign in_dat_data_int8_8 = { cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8], cfg_is_int8_d1[8] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27565" *) { in_dat_data72, in_dat_data8 };
  assign in_dat_data_int8_7 = { cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7], cfg_is_int8_d1[7] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27566" *) { in_dat_data71, in_dat_data7 };
  assign in_dat_data_int8_6 = { cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6], cfg_is_int8_d1[6] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27567" *) { in_dat_data70, in_dat_data6 };
  assign in_dat_data_int8_5 = { cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5], cfg_is_int8_d1[5] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27568" *) { in_dat_data69, in_dat_data5 };
  assign in_dat_data_int8_4 = { cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4], cfg_is_int8_d1[4] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27569" *) { in_dat_data68, in_dat_data4 };
  assign in_wt_norm[33] = cfg_is_fp16_d1[33] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2757" *) _08169_;
  assign in_dat_data_int8_3 = { cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3], cfg_is_int8_d1[3] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27570" *) { in_dat_data67, in_dat_data3 };
  assign in_dat_data_int8_2 = { cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2], cfg_is_int8_d1[2] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27571" *) { in_dat_data66, in_dat_data2 };
  assign in_dat_data_int8_1 = { cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1], cfg_is_int8_d1[1] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27572" *) { in_dat_data65, in_dat_data1 };
  assign in_dat_data_int8_0 = { cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0], cfg_is_int8_d1[0] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27573" *) { in_dat_data64, in_dat_data0 };
  assign in_wt_norm[32] = cfg_is_fp16_d1[32] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2758" *) _08170_;
  assign in_wt_norm[31] = cfg_is_fp16_d1[31] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2759" *) _08171_;
  assign in_wt_norm[30] = cfg_is_fp16_d1[30] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2760" *) _08172_;
  assign in_wt_norm[29] = cfg_is_fp16_d1[29] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2761" *) _08173_;
  assign in_wt_norm[28] = cfg_is_fp16_d1[28] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2762" *) _08174_;
  assign in_wt_norm[27] = cfg_is_fp16_d1[27] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2763" *) _08175_;
  assign in_wt_norm[26] = cfg_is_fp16_d1[26] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2764" *) _08176_;
  assign in_wt_norm[25] = cfg_is_fp16_d1[25] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2765" *) _08177_;
  assign in_wt_norm[24] = cfg_is_fp16_d1[24] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2766" *) _08178_;
  assign _05233_ = cfg_is_fp16_d1[63] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *) _08011_;
  assign _05234_ = _05233_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *) _08179_;
  assign in_dat_nan[63] = _05234_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *) in_dat_mask[126];
  assign _05235_ = cfg_is_fp16_d1[62] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *) _08012_;
  assign _05236_ = _05235_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *) _08180_;
  assign in_dat_nan[62] = _05236_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *) in_dat_mask[124];
  assign _05237_ = cfg_is_fp16_d1[61] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *) _08013_;
  assign _05238_ = _05237_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *) _08181_;
  assign in_dat_nan[61] = _05238_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *) in_dat_mask[122];
  assign _05239_ = cfg_is_fp16_d1[60] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *) _08014_;
  assign _05240_ = _05239_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *) _08182_;
  assign in_dat_nan[60] = _05240_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *) in_dat_mask[120];
  assign _05241_ = cfg_is_fp16_d1[59] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *) _08015_;
  assign _05242_ = _05241_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *) _08183_;
  assign in_dat_nan[59] = _05242_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *) in_dat_mask[118];
  assign _05243_ = cfg_is_fp16_d1[58] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *) _08016_;
  assign _05244_ = _05243_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *) _08184_;
  assign in_dat_nan[58] = _05244_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *) in_dat_mask[116];
  assign _05245_ = cfg_is_fp16_d1[57] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *) _08017_;
  assign _05246_ = _05245_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *) _08185_;
  assign in_dat_nan[57] = _05246_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *) in_dat_mask[114];
  assign _05247_ = cfg_is_fp16_d1[56] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *) _08018_;
  assign _05248_ = _05247_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *) _08186_;
  assign in_dat_nan[56] = _05248_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *) in_dat_mask[112];
  assign _05249_ = cfg_is_fp16_d1[55] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *) _08019_;
  assign _05250_ = _05249_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *) _08187_;
  assign in_dat_nan[55] = _05250_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *) in_dat_mask[110];
  assign in_wt_norm[23] = cfg_is_fp16_d1[23] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2767" *) _08188_;
  assign _05251_ = cfg_is_fp16_d1[54] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *) _08020_;
  assign _05252_ = _05251_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *) _08189_;
  assign in_dat_nan[54] = _05252_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *) in_dat_mask[108];
  assign _05253_ = cfg_is_fp16_d1[53] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *) _08021_;
  assign _05254_ = _05253_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *) _08190_;
  assign in_dat_nan[53] = _05254_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *) in_dat_mask[106];
  assign _05255_ = cfg_is_fp16_d1[52] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *) _08022_;
  assign _05256_ = _05255_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *) _08191_;
  assign in_dat_nan[52] = _05256_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *) in_dat_mask[104];
  assign _05257_ = cfg_is_fp16_d1[51] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *) _08023_;
  assign _05258_ = _05257_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *) _08192_;
  assign in_dat_nan[51] = _05258_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *) in_dat_mask[102];
  assign _05259_ = cfg_is_fp16_d1[50] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *) _08024_;
  assign _05260_ = _05259_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *) _08193_;
  assign in_dat_nan[50] = _05260_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *) in_dat_mask[100];
  assign _05261_ = cfg_is_fp16_d1[49] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *) _08025_;
  assign _05262_ = _05261_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *) _08194_;
  assign in_dat_nan[49] = _05262_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *) in_dat_mask[98];
  assign _05263_ = cfg_is_fp16_d1[48] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *) _08026_;
  assign _05264_ = _05263_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *) _08195_;
  assign in_dat_nan[48] = _05264_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *) in_dat_mask[96];
  assign _05265_ = cfg_is_fp16_d1[47] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *) _08027_;
  assign _05266_ = _05265_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *) _08196_;
  assign in_dat_nan[47] = _05266_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *) in_dat_mask[94];
  assign _05267_ = cfg_is_fp16_d1[46] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *) _08028_;
  assign _05268_ = _05267_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *) _08197_;
  assign in_dat_nan[46] = _05268_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *) in_dat_mask[92];
  assign _05269_ = cfg_is_fp16_d1[45] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *) _08029_;
  assign _05270_ = _05269_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *) _08198_;
  assign in_dat_nan[45] = _05270_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *) in_dat_mask[90];
  assign in_wt_norm[22] = cfg_is_fp16_d1[22] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2768" *) _08199_;
  assign _05271_ = cfg_is_fp16_d1[44] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *) _08030_;
  assign _05272_ = _05271_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *) _08200_;
  assign in_dat_nan[44] = _05272_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *) in_dat_mask[88];
  assign _05273_ = cfg_is_fp16_d1[43] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *) _08031_;
  assign _05274_ = _05273_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *) _08201_;
  assign in_dat_nan[43] = _05274_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *) in_dat_mask[86];
  assign _05275_ = cfg_is_fp16_d1[42] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *) _08032_;
  assign _05276_ = _05275_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *) _08202_;
  assign in_dat_nan[42] = _05276_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *) in_dat_mask[84];
  assign _05277_ = cfg_is_fp16_d1[41] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *) _08033_;
  assign _05278_ = _05277_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *) _08203_;
  assign in_dat_nan[41] = _05278_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *) in_dat_mask[82];
  assign _05279_ = cfg_is_fp16_d1[40] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *) _08034_;
  assign _05280_ = _05279_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *) _08204_;
  assign in_dat_nan[40] = _05280_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *) in_dat_mask[80];
  assign _05281_ = cfg_is_fp16_d1[39] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *) _08035_;
  assign _05282_ = _05281_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *) _08205_;
  assign in_dat_nan[39] = _05282_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *) in_dat_mask[78];
  assign _05283_ = cfg_is_fp16_d1[38] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *) _08036_;
  assign _05284_ = _05283_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *) _08206_;
  assign in_dat_nan[38] = _05284_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *) in_dat_mask[76];
  assign _05285_ = cfg_is_fp16_d1[37] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *) _08037_;
  assign _05286_ = _05285_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *) _08207_;
  assign in_dat_nan[37] = _05286_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *) in_dat_mask[74];
  assign _05287_ = cfg_is_fp16_d1[36] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *) _08038_;
  assign _05288_ = _05287_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *) _08208_;
  assign in_dat_nan[36] = _05288_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *) in_dat_mask[72];
  assign _05289_ = cfg_is_fp16_d1[35] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *) _08039_;
  assign _05290_ = _05289_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *) _08209_;
  assign in_dat_nan[35] = _05290_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *) in_dat_mask[70];
  assign in_wt_norm[21] = cfg_is_fp16_d1[21] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2769" *) _08210_;
  assign _05291_ = cfg_is_fp16_d1[34] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *) _08040_;
  assign _05292_ = _05291_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *) _08211_;
  assign in_dat_nan[34] = _05292_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *) in_dat_mask[68];
  assign _05293_ = cfg_is_fp16_d1[33] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *) _08041_;
  assign _05294_ = _05293_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *) _08212_;
  assign in_dat_nan[33] = _05294_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *) in_dat_mask[66];
  assign _05295_ = cfg_is_fp16_d1[32] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *) _08042_;
  assign _05296_ = _05295_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *) _08213_;
  assign in_dat_nan[32] = _05296_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *) in_dat_mask[64];
  assign _05297_ = cfg_is_fp16_d1[31] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *) _08043_;
  assign _05298_ = _05297_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *) _08214_;
  assign in_dat_nan[31] = _05298_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *) in_dat_mask[62];
  assign _05299_ = cfg_is_fp16_d1[30] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *) _08044_;
  assign _05300_ = _05299_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *) _08215_;
  assign in_dat_nan[30] = _05300_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *) in_dat_mask[60];
  assign _05301_ = cfg_is_fp16_d1[29] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *) _08045_;
  assign _05302_ = _05301_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *) _08216_;
  assign in_dat_nan[29] = _05302_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *) in_dat_mask[58];
  assign _05303_ = cfg_is_fp16_d1[28] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *) _08046_;
  assign _05304_ = _05303_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *) _08217_;
  assign in_dat_nan[28] = _05304_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *) in_dat_mask[56];
  assign _05305_ = cfg_is_fp16_d1[27] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *) _08047_;
  assign _05306_ = _05305_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *) _08218_;
  assign in_dat_nan[27] = _05306_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *) in_dat_mask[54];
  assign _05307_ = cfg_is_fp16_d1[26] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *) _08048_;
  assign _05308_ = _05307_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *) _08219_;
  assign in_dat_nan[26] = _05308_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *) in_dat_mask[52];
  assign _05309_ = cfg_is_fp16_d1[25] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *) _08049_;
  assign _05310_ = _05309_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *) _08220_;
  assign in_dat_nan[25] = _05310_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *) in_dat_mask[50];
  assign in_wt_norm[20] = cfg_is_fp16_d1[20] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2770" *) _08221_;
  assign _05311_ = cfg_is_fp16_d1[24] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *) _08050_;
  assign _05312_ = _05311_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *) _08222_;
  assign in_dat_nan[24] = _05312_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *) in_dat_mask[48];
  assign _05313_ = cfg_is_fp16_d1[23] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *) _08051_;
  assign _05314_ = _05313_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *) _08223_;
  assign in_dat_nan[23] = _05314_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *) in_dat_mask[46];
  assign _05315_ = cfg_is_fp16_d1[22] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *) _08052_;
  assign _05316_ = _05315_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *) _08224_;
  assign in_dat_nan[22] = _05316_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *) in_dat_mask[44];
  assign _05317_ = cfg_is_fp16_d1[21] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *) _08053_;
  assign _05318_ = _05317_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *) _08225_;
  assign in_dat_nan[21] = _05318_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *) in_dat_mask[42];
  assign _05319_ = cfg_is_fp16_d1[20] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *) _08054_;
  assign _05320_ = _05319_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *) _08226_;
  assign in_dat_nan[20] = _05320_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *) in_dat_mask[40];
  assign _05321_ = cfg_is_fp16_d1[19] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *) _08055_;
  assign _05322_ = _05321_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *) _08227_;
  assign in_dat_nan[19] = _05322_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *) in_dat_mask[38];
  assign _05323_ = cfg_is_fp16_d1[18] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *) _08056_;
  assign _05324_ = _05323_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *) _08228_;
  assign in_dat_nan[18] = _05324_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *) in_dat_mask[36];
  assign _05325_ = cfg_is_fp16_d1[17] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *) _08057_;
  assign _05326_ = _05325_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *) _08229_;
  assign in_dat_nan[17] = _05326_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *) in_dat_mask[34];
  assign _05327_ = cfg_is_fp16_d1[16] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *) _08058_;
  assign _05328_ = _05327_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *) _08230_;
  assign in_dat_nan[16] = _05328_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *) in_dat_mask[32];
  assign _05329_ = cfg_is_fp16_d1[15] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *) _08059_;
  assign _05330_ = _05329_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *) _08231_;
  assign in_dat_nan[15] = _05330_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *) in_dat_mask[30];
  assign in_wt_norm[19] = cfg_is_fp16_d1[19] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2771" *) _08232_;
  assign _05331_ = cfg_is_fp16_d1[14] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *) _08060_;
  assign _05332_ = _05331_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *) _08233_;
  assign in_dat_nan[14] = _05332_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *) in_dat_mask[28];
  assign _05333_ = cfg_is_fp16_d1[13] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *) _08061_;
  assign _05334_ = _05333_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *) _08234_;
  assign in_dat_nan[13] = _05334_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *) in_dat_mask[26];
  assign _05335_ = cfg_is_fp16_d1[12] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *) _08062_;
  assign _05336_ = _05335_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *) _08235_;
  assign in_dat_nan[12] = _05336_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *) in_dat_mask[24];
  assign _05337_ = cfg_is_fp16_d1[11] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *) _08063_;
  assign _05338_ = _05337_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *) _08236_;
  assign in_dat_nan[11] = _05338_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *) in_dat_mask[22];
  assign _05339_ = cfg_is_fp16_d1[10] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *) _08064_;
  assign _05340_ = _05339_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *) _08237_;
  assign in_dat_nan[10] = _05340_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *) in_dat_mask[20];
  assign _05341_ = cfg_is_fp16_d1[9] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *) _08065_;
  assign _05342_ = _05341_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *) _08238_;
  assign in_dat_nan[9] = _05342_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *) in_dat_mask[18];
  assign _05343_ = cfg_is_fp16_d1[8] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *) _08066_;
  assign _05344_ = _05343_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *) _08239_;
  assign in_dat_nan[8] = _05344_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *) in_dat_mask[16];
  assign _05345_ = cfg_is_fp16_d1[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *) _08067_;
  assign _05346_ = _05345_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *) _08240_;
  assign in_dat_nan[7] = _05346_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *) in_dat_mask[14];
  assign _05347_ = cfg_is_fp16_d1[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *) _08068_;
  assign _05348_ = _05347_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *) _08241_;
  assign in_dat_nan[6] = _05348_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *) in_dat_mask[12];
  assign _05349_ = cfg_is_fp16_d1[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *) _08069_;
  assign _05350_ = _05349_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *) _08242_;
  assign in_dat_nan[5] = _05350_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *) in_dat_mask[10];
  assign in_wt_norm[18] = cfg_is_fp16_d1[18] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2772" *) _08243_;
  assign _05351_ = cfg_is_fp16_d1[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *) _08070_;
  assign _05352_ = _05351_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *) _08244_;
  assign in_dat_nan[4] = _05352_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *) in_dat_mask[8];
  assign _05353_ = cfg_is_fp16_d1[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *) _08071_;
  assign _05354_ = _05353_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *) _08245_;
  assign in_dat_nan[3] = _05354_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *) in_dat_mask[6];
  assign _05355_ = cfg_is_fp16_d1[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *) _08072_;
  assign _05356_ = _05355_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *) _08246_;
  assign in_dat_nan[2] = _05356_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *) in_dat_mask[4];
  assign _05357_ = cfg_is_fp16_d1[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *) _08073_;
  assign _05358_ = _05357_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *) _08247_;
  assign in_dat_nan[1] = _05358_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *) in_dat_mask[2];
  assign _05359_ = cfg_is_fp16_d1[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *) _08074_;
  assign _05360_ = _05359_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *) _08248_;
  assign in_dat_nan[0] = _05360_ & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *) in_dat_mask[0];
  assign in_wt_norm[17] = cfg_is_fp16_d1[17] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2773" *) _08249_;
  assign _05361_ = cfg_is_fp16_d1[63] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27731" *) in_dat_mask[127];
  assign dat_pre_exp_w[191:189] = { _05361_, _05361_, _05361_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27731" *) in_dat_data127[6:4];
  assign _05362_ = cfg_is_fp16_d1[62] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27732" *) in_dat_mask[125];
  assign dat_pre_exp_w[188:186] = { _05362_, _05362_, _05362_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27732" *) in_dat_data125[6:4];
  assign _05363_ = cfg_is_fp16_d1[61] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27733" *) in_dat_mask[123];
  assign dat_pre_exp_w[185:183] = { _05363_, _05363_, _05363_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27733" *) in_dat_data123[6:4];
  assign _05364_ = cfg_is_fp16_d1[60] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27734" *) in_dat_mask[121];
  assign dat_pre_exp_w[182:180] = { _05364_, _05364_, _05364_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27734" *) in_dat_data121[6:4];
  assign _05365_ = cfg_is_fp16_d1[59] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27735" *) in_dat_mask[119];
  assign dat_pre_exp_w[179:177] = { _05365_, _05365_, _05365_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27735" *) in_dat_data119[6:4];
  assign _05366_ = cfg_is_fp16_d1[58] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27736" *) in_dat_mask[117];
  assign dat_pre_exp_w[176:174] = { _05366_, _05366_, _05366_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27736" *) in_dat_data117[6:4];
  assign _05367_ = cfg_is_fp16_d1[57] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27737" *) in_dat_mask[115];
  assign dat_pre_exp_w[173:171] = { _05367_, _05367_, _05367_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27737" *) in_dat_data115[6:4];
  assign _05368_ = cfg_is_fp16_d1[56] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27738" *) in_dat_mask[113];
  assign dat_pre_exp_w[170:168] = { _05368_, _05368_, _05368_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27738" *) in_dat_data113[6:4];
  assign _05369_ = cfg_is_fp16_d1[55] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27739" *) in_dat_mask[111];
  assign dat_pre_exp_w[167:165] = { _05369_, _05369_, _05369_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27739" *) in_dat_data111[6:4];
  assign in_wt_norm[16] = cfg_is_fp16_d1[16] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2774" *) _08250_;
  assign _05370_ = cfg_is_fp16_d1[54] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27740" *) in_dat_mask[109];
  assign dat_pre_exp_w[164:162] = { _05370_, _05370_, _05370_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27740" *) in_dat_data109[6:4];
  assign _05371_ = cfg_is_fp16_d1[53] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27741" *) in_dat_mask[107];
  assign dat_pre_exp_w[161:159] = { _05371_, _05371_, _05371_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27741" *) in_dat_data107[6:4];
  assign _05372_ = cfg_is_fp16_d1[52] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27742" *) in_dat_mask[105];
  assign dat_pre_exp_w[158:156] = { _05372_, _05372_, _05372_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27742" *) in_dat_data105[6:4];
  assign _05373_ = cfg_is_fp16_d1[51] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27743" *) in_dat_mask[103];
  assign dat_pre_exp_w[155:153] = { _05373_, _05373_, _05373_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27743" *) in_dat_data103[6:4];
  assign _05374_ = cfg_is_fp16_d1[50] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27744" *) in_dat_mask[101];
  assign dat_pre_exp_w[152:150] = { _05374_, _05374_, _05374_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27744" *) in_dat_data101[6:4];
  assign _05375_ = cfg_is_fp16_d1[49] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27745" *) in_dat_mask[99];
  assign dat_pre_exp_w[149:147] = { _05375_, _05375_, _05375_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27745" *) in_dat_data99[6:4];
  assign _05376_ = cfg_is_fp16_d1[48] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27746" *) in_dat_mask[97];
  assign dat_pre_exp_w[146:144] = { _05376_, _05376_, _05376_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27746" *) in_dat_data97[6:4];
  assign _05377_ = cfg_is_fp16_d1[47] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27747" *) in_dat_mask[95];
  assign dat_pre_exp_w[143:141] = { _05377_, _05377_, _05377_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27747" *) in_dat_data95[6:4];
  assign _05378_ = cfg_is_fp16_d1[46] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27748" *) in_dat_mask[93];
  assign dat_pre_exp_w[140:138] = { _05378_, _05378_, _05378_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27748" *) in_dat_data93[6:4];
  assign _05379_ = cfg_is_fp16_d1[45] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27749" *) in_dat_mask[91];
  assign dat_pre_exp_w[137:135] = { _05379_, _05379_, _05379_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27749" *) in_dat_data91[6:4];
  assign in_wt_norm[15] = cfg_is_fp16_d1[15] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2775" *) _08251_;
  assign _05380_ = cfg_is_fp16_d1[44] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27750" *) in_dat_mask[89];
  assign dat_pre_exp_w[134:132] = { _05380_, _05380_, _05380_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27750" *) in_dat_data89[6:4];
  assign _05381_ = cfg_is_fp16_d1[43] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27751" *) in_dat_mask[87];
  assign dat_pre_exp_w[131:129] = { _05381_, _05381_, _05381_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27751" *) in_dat_data87[6:4];
  assign _05382_ = cfg_is_fp16_d1[42] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27752" *) in_dat_mask[85];
  assign dat_pre_exp_w[128:126] = { _05382_, _05382_, _05382_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27752" *) in_dat_data85[6:4];
  assign _05383_ = cfg_is_fp16_d1[41] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27753" *) in_dat_mask[83];
  assign dat_pre_exp_w[125:123] = { _05383_, _05383_, _05383_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27753" *) in_dat_data83[6:4];
  assign _05384_ = cfg_is_fp16_d1[40] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27754" *) in_dat_mask[81];
  assign dat_pre_exp_w[122:120] = { _05384_, _05384_, _05384_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27754" *) in_dat_data81[6:4];
  assign _05385_ = cfg_is_fp16_d1[39] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27755" *) in_dat_mask[79];
  assign dat_pre_exp_w[119:117] = { _05385_, _05385_, _05385_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27755" *) in_dat_data79[6:4];
  assign _05386_ = cfg_is_fp16_d1[38] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27756" *) in_dat_mask[77];
  assign dat_pre_exp_w[116:114] = { _05386_, _05386_, _05386_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27756" *) in_dat_data77[6:4];
  assign _05387_ = cfg_is_fp16_d1[37] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27757" *) in_dat_mask[75];
  assign dat_pre_exp_w[113:111] = { _05387_, _05387_, _05387_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27757" *) in_dat_data75[6:4];
  assign _05388_ = cfg_is_fp16_d1[36] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27758" *) in_dat_mask[73];
  assign dat_pre_exp_w[110:108] = { _05388_, _05388_, _05388_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27758" *) in_dat_data73[6:4];
  assign _05389_ = cfg_is_fp16_d1[35] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27759" *) in_dat_mask[71];
  assign dat_pre_exp_w[107:105] = { _05389_, _05389_, _05389_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27759" *) in_dat_data71[6:4];
  assign in_wt_norm[14] = cfg_is_fp16_d1[14] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2776" *) _08252_;
  assign _05390_ = cfg_is_fp16_d1[34] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27760" *) in_dat_mask[69];
  assign dat_pre_exp_w[104:102] = { _05390_, _05390_, _05390_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27760" *) in_dat_data69[6:4];
  assign _05391_ = cfg_is_fp16_d1[33] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27761" *) in_dat_mask[67];
  assign dat_pre_exp_w[101:99] = { _05391_, _05391_, _05391_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27761" *) in_dat_data67[6:4];
  assign _05392_ = cfg_is_fp16_d1[32] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27762" *) in_dat_mask[65];
  assign dat_pre_exp_w[98:96] = { _05392_, _05392_, _05392_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27762" *) in_dat_data65[6:4];
  assign _05393_ = cfg_is_fp16_d1[31] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27763" *) in_dat_mask[63];
  assign dat_pre_exp_w[95:93] = { _05393_, _05393_, _05393_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27763" *) in_dat_data63[6:4];
  assign _05394_ = cfg_is_fp16_d1[30] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27764" *) in_dat_mask[61];
  assign dat_pre_exp_w[92:90] = { _05394_, _05394_, _05394_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27764" *) in_dat_data61[6:4];
  assign _05395_ = cfg_is_fp16_d1[29] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27765" *) in_dat_mask[59];
  assign dat_pre_exp_w[89:87] = { _05395_, _05395_, _05395_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27765" *) in_dat_data59[6:4];
  assign _05396_ = cfg_is_fp16_d1[28] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27766" *) in_dat_mask[57];
  assign dat_pre_exp_w[86:84] = { _05396_, _05396_, _05396_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27766" *) in_dat_data57[6:4];
  assign _05397_ = cfg_is_fp16_d1[27] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27767" *) in_dat_mask[55];
  assign dat_pre_exp_w[83:81] = { _05397_, _05397_, _05397_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27767" *) in_dat_data55[6:4];
  assign _05398_ = cfg_is_fp16_d1[26] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27768" *) in_dat_mask[53];
  assign dat_pre_exp_w[80:78] = { _05398_, _05398_, _05398_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27768" *) in_dat_data53[6:4];
  assign _05399_ = cfg_is_fp16_d1[25] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27769" *) in_dat_mask[51];
  assign dat_pre_exp_w[77:75] = { _05399_, _05399_, _05399_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27769" *) in_dat_data51[6:4];
  assign in_wt_norm[13] = cfg_is_fp16_d1[13] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2777" *) _08253_;
  assign _05400_ = cfg_is_fp16_d1[24] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27770" *) in_dat_mask[49];
  assign dat_pre_exp_w[74:72] = { _05400_, _05400_, _05400_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27770" *) in_dat_data49[6:4];
  assign _05401_ = cfg_is_fp16_d1[23] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27771" *) in_dat_mask[47];
  assign dat_pre_exp_w[71:69] = { _05401_, _05401_, _05401_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27771" *) in_dat_data47[6:4];
  assign _05402_ = cfg_is_fp16_d1[22] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27772" *) in_dat_mask[45];
  assign dat_pre_exp_w[68:66] = { _05402_, _05402_, _05402_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27772" *) in_dat_data45[6:4];
  assign _05403_ = cfg_is_fp16_d1[21] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27773" *) in_dat_mask[43];
  assign dat_pre_exp_w[65:63] = { _05403_, _05403_, _05403_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27773" *) in_dat_data43[6:4];
  assign _05404_ = cfg_is_fp16_d1[20] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27774" *) in_dat_mask[41];
  assign dat_pre_exp_w[62:60] = { _05404_, _05404_, _05404_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27774" *) in_dat_data41[6:4];
  assign _05405_ = cfg_is_fp16_d1[19] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27775" *) in_dat_mask[39];
  assign dat_pre_exp_w[59:57] = { _05405_, _05405_, _05405_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27775" *) in_dat_data39[6:4];
  assign _05406_ = cfg_is_fp16_d1[18] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27776" *) in_dat_mask[37];
  assign dat_pre_exp_w[56:54] = { _05406_, _05406_, _05406_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27776" *) in_dat_data37[6:4];
  assign _05407_ = cfg_is_fp16_d1[17] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27777" *) in_dat_mask[35];
  assign dat_pre_exp_w[53:51] = { _05407_, _05407_, _05407_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27777" *) in_dat_data35[6:4];
  assign _05408_ = cfg_is_fp16_d1[16] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27778" *) in_dat_mask[33];
  assign dat_pre_exp_w[50:48] = { _05408_, _05408_, _05408_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27778" *) in_dat_data33[6:4];
  assign _05409_ = cfg_is_fp16_d1[15] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27779" *) in_dat_mask[31];
  assign dat_pre_exp_w[47:45] = { _05409_, _05409_, _05409_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27779" *) in_dat_data31[6:4];
  assign in_wt_norm[12] = cfg_is_fp16_d1[12] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2778" *) _08254_;
  assign _05410_ = cfg_is_fp16_d1[14] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27780" *) in_dat_mask[29];
  assign dat_pre_exp_w[44:42] = { _05410_, _05410_, _05410_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27780" *) in_dat_data29[6:4];
  assign _05411_ = cfg_is_fp16_d1[13] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27781" *) in_dat_mask[27];
  assign dat_pre_exp_w[41:39] = { _05411_, _05411_, _05411_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27781" *) in_dat_data27[6:4];
  assign _05412_ = cfg_is_fp16_d1[12] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27782" *) in_dat_mask[25];
  assign dat_pre_exp_w[38:36] = { _05412_, _05412_, _05412_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27782" *) in_dat_data25[6:4];
  assign _05413_ = cfg_is_fp16_d1[11] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27783" *) in_dat_mask[23];
  assign dat_pre_exp_w[35:33] = { _05413_, _05413_, _05413_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27783" *) in_dat_data23[6:4];
  assign _05414_ = cfg_is_fp16_d1[10] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27784" *) in_dat_mask[21];
  assign dat_pre_exp_w[32:30] = { _05414_, _05414_, _05414_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27784" *) in_dat_data21[6:4];
  assign _05415_ = cfg_is_fp16_d1[9] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27785" *) in_dat_mask[19];
  assign dat_pre_exp_w[29:27] = { _05415_, _05415_, _05415_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27785" *) in_dat_data19[6:4];
  assign _05416_ = cfg_is_fp16_d1[8] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27786" *) in_dat_mask[17];
  assign dat_pre_exp_w[26:24] = { _05416_, _05416_, _05416_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27786" *) in_dat_data17[6:4];
  assign _05417_ = cfg_is_fp16_d1[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27787" *) in_dat_mask[15];
  assign dat_pre_exp_w[23:21] = { _05417_, _05417_, _05417_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27787" *) in_dat_data15[6:4];
  assign _05418_ = cfg_is_fp16_d1[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27788" *) in_dat_mask[13];
  assign dat_pre_exp_w[20:18] = { _05418_, _05418_, _05418_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27788" *) in_dat_data13[6:4];
  assign _05419_ = cfg_is_fp16_d1[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27789" *) in_dat_mask[11];
  assign dat_pre_exp_w[17:15] = { _05419_, _05419_, _05419_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27789" *) in_dat_data11[6:4];
  assign in_wt_norm[11] = cfg_is_fp16_d1[11] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2779" *) _08255_;
  assign _05420_ = cfg_is_fp16_d1[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27790" *) in_dat_mask[9];
  assign dat_pre_exp_w[14:12] = { _05420_, _05420_, _05420_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27790" *) in_dat_data9[6:4];
  assign _05421_ = cfg_is_fp16_d1[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27791" *) in_dat_mask[7];
  assign dat_pre_exp_w[11:9] = { _05421_, _05421_, _05421_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27791" *) in_dat_data7[6:4];
  assign _05422_ = cfg_is_fp16_d1[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27792" *) in_dat_mask[5];
  assign dat_pre_exp_w[8:6] = { _05422_, _05422_, _05422_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27792" *) in_dat_data5[6:4];
  assign _05423_ = cfg_is_fp16_d1[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27793" *) in_dat_mask[3];
  assign dat_pre_exp_w[5:3] = { _05423_, _05423_, _05423_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27793" *) in_dat_data3[6:4];
  assign _05424_ = cfg_is_fp16_d1[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27794" *) in_dat_mask[1];
  assign dat_pre_exp_w[2:0] = { _05424_, _05424_, _05424_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27794" *) in_dat_data1[6:4];
  assign in_wt_norm[10] = cfg_is_fp16_d1[10] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2780" *) _08256_;
  assign in_dat_norm[63] = cfg_is_fp16_d1[63] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27800" *) _08257_;
  assign in_dat_norm[62] = cfg_is_fp16_d1[62] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27801" *) _08258_;
  assign in_dat_norm[61] = cfg_is_fp16_d1[61] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27802" *) _08259_;
  assign in_dat_norm[60] = cfg_is_fp16_d1[60] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27803" *) _08260_;
  assign in_dat_norm[59] = cfg_is_fp16_d1[59] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27804" *) _08261_;
  assign in_dat_norm[58] = cfg_is_fp16_d1[58] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27805" *) _08262_;
  assign in_dat_norm[57] = cfg_is_fp16_d1[57] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27806" *) _08263_;
  assign in_dat_norm[56] = cfg_is_fp16_d1[56] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27807" *) _08264_;
  assign in_dat_norm[55] = cfg_is_fp16_d1[55] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27808" *) _08265_;
  assign in_dat_norm[54] = cfg_is_fp16_d1[54] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27809" *) _08266_;
  assign in_wt_norm[9] = cfg_is_fp16_d1[9] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2781" *) _08267_;
  assign in_dat_norm[53] = cfg_is_fp16_d1[53] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27810" *) _08268_;
  assign in_dat_norm[52] = cfg_is_fp16_d1[52] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27811" *) _08269_;
  assign in_dat_norm[51] = cfg_is_fp16_d1[51] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27812" *) _08270_;
  assign in_dat_norm[50] = cfg_is_fp16_d1[50] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27813" *) _08271_;
  assign in_dat_norm[49] = cfg_is_fp16_d1[49] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27814" *) _08272_;
  assign in_dat_norm[48] = cfg_is_fp16_d1[48] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27815" *) _08273_;
  assign in_dat_norm[47] = cfg_is_fp16_d1[47] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27816" *) _08274_;
  assign in_dat_norm[46] = cfg_is_fp16_d1[46] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27817" *) _08275_;
  assign in_dat_norm[45] = cfg_is_fp16_d1[45] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27818" *) _08276_;
  assign in_dat_norm[44] = cfg_is_fp16_d1[44] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27819" *) _08277_;
  assign in_wt_norm[8] = cfg_is_fp16_d1[8] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2782" *) _08278_;
  assign in_dat_norm[43] = cfg_is_fp16_d1[43] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27820" *) _08279_;
  assign in_dat_norm[42] = cfg_is_fp16_d1[42] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27821" *) _08280_;
  assign in_dat_norm[41] = cfg_is_fp16_d1[41] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27822" *) _08281_;
  assign in_dat_norm[40] = cfg_is_fp16_d1[40] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27823" *) _08282_;
  assign in_dat_norm[39] = cfg_is_fp16_d1[39] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27824" *) _08283_;
  assign in_dat_norm[38] = cfg_is_fp16_d1[38] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27825" *) _08284_;
  assign in_dat_norm[37] = cfg_is_fp16_d1[37] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27826" *) _08285_;
  assign in_dat_norm[36] = cfg_is_fp16_d1[36] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27827" *) _08286_;
  assign in_dat_norm[35] = cfg_is_fp16_d1[35] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27828" *) _08287_;
  assign in_dat_norm[34] = cfg_is_fp16_d1[34] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27829" *) _08288_;
  assign in_wt_norm[7] = cfg_is_fp16_d1[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2783" *) _08289_;
  assign in_dat_norm[33] = cfg_is_fp16_d1[33] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27830" *) _08290_;
  assign in_dat_norm[32] = cfg_is_fp16_d1[32] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27831" *) _08291_;
  assign in_dat_norm[31] = cfg_is_fp16_d1[31] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27832" *) _08292_;
  assign in_dat_norm[30] = cfg_is_fp16_d1[30] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27833" *) _08293_;
  assign in_dat_norm[29] = cfg_is_fp16_d1[29] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27834" *) _08294_;
  assign in_dat_norm[28] = cfg_is_fp16_d1[28] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27835" *) _08295_;
  assign in_dat_norm[27] = cfg_is_fp16_d1[27] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27836" *) _08296_;
  assign in_dat_norm[26] = cfg_is_fp16_d1[26] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27837" *) _08297_;
  assign in_dat_norm[25] = cfg_is_fp16_d1[25] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27838" *) _08298_;
  assign in_dat_norm[24] = cfg_is_fp16_d1[24] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27839" *) _08299_;
  assign in_wt_norm[6] = cfg_is_fp16_d1[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2784" *) _08300_;
  assign in_dat_norm[23] = cfg_is_fp16_d1[23] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27840" *) _08301_;
  assign in_dat_norm[22] = cfg_is_fp16_d1[22] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27841" *) _08302_;
  assign in_dat_norm[21] = cfg_is_fp16_d1[21] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27842" *) _08303_;
  assign in_dat_norm[20] = cfg_is_fp16_d1[20] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27843" *) _08304_;
  assign in_dat_norm[19] = cfg_is_fp16_d1[19] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27844" *) _08305_;
  assign in_dat_norm[18] = cfg_is_fp16_d1[18] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27845" *) _08306_;
  assign in_dat_norm[17] = cfg_is_fp16_d1[17] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27846" *) _08307_;
  assign in_dat_norm[16] = cfg_is_fp16_d1[16] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27847" *) _08308_;
  assign in_dat_norm[15] = cfg_is_fp16_d1[15] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27848" *) _08309_;
  assign in_dat_norm[14] = cfg_is_fp16_d1[14] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27849" *) _08310_;
  assign in_wt_norm[5] = cfg_is_fp16_d1[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2785" *) _08311_;
  assign in_dat_norm[13] = cfg_is_fp16_d1[13] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27850" *) _08312_;
  assign in_dat_norm[12] = cfg_is_fp16_d1[12] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27851" *) _08313_;
  assign in_dat_norm[11] = cfg_is_fp16_d1[11] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27852" *) _08314_;
  assign in_dat_norm[10] = cfg_is_fp16_d1[10] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27853" *) _08315_;
  assign in_dat_norm[9] = cfg_is_fp16_d1[9] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27854" *) _08316_;
  assign in_dat_norm[8] = cfg_is_fp16_d1[8] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27855" *) _08317_;
  assign in_dat_norm[7] = cfg_is_fp16_d1[7] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27856" *) _08318_;
  assign in_dat_norm[6] = cfg_is_fp16_d1[6] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27857" *) _08319_;
  assign in_dat_norm[5] = cfg_is_fp16_d1[5] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27858" *) _08320_;
  assign in_dat_norm[4] = cfg_is_fp16_d1[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27859" *) _08321_;
  assign in_wt_norm[4] = cfg_is_fp16_d1[4] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2786" *) _08322_;
  assign in_dat_norm[3] = cfg_is_fp16_d1[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27860" *) _08323_;
  assign in_dat_norm[2] = cfg_is_fp16_d1[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27861" *) _08324_;
  assign in_dat_norm[1] = cfg_is_fp16_d1[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27862" *) _08325_;
  assign in_dat_norm[0] = cfg_is_fp16_d1[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27863" *) _08326_;
  assign in_wt_norm[3] = cfg_is_fp16_d1[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2787" *) _08327_;
  assign in_wt_norm[2] = cfg_is_fp16_d1[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2788" *) _08328_;
  assign in_wt_norm[1] = cfg_is_fp16_d1[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2789" *) _08329_;
  assign in_wt_norm[0] = cfg_is_fp16_d1[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2790" *) _08330_;
  assign in_dat_data_fp16_63 = { cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28447" *) { in_dat_data127[7], in_dat_data_fp16_mts_sft63 };
  assign in_dat_data_fp16_62 = { cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28455" *) { in_dat_data125[7], in_dat_data_fp16_mts_sft62 };
  assign in_dat_data_fp16_61 = { cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28463" *) { in_dat_data123[7], in_dat_data_fp16_mts_sft61 };
  assign in_dat_data_fp16_60 = { cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28471" *) { in_dat_data121[7], in_dat_data_fp16_mts_sft60 };
  assign in_dat_data_fp16_59 = { cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28479" *) { in_dat_data119[7], in_dat_data_fp16_mts_sft59 };
  assign in_dat_data_fp16_58 = { cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28487" *) { in_dat_data117[7], in_dat_data_fp16_mts_sft58 };
  assign in_dat_data_fp16_57 = { cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28495" *) { in_dat_data115[7], in_dat_data_fp16_mts_sft57 };
  assign in_dat_data_fp16_56 = { cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28503" *) { in_dat_data113[7], in_dat_data_fp16_mts_sft56 };
  assign in_dat_data_fp16_55 = { cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28511" *) { in_dat_data111[7], in_dat_data_fp16_mts_sft55 };
  assign in_dat_data_fp16_54 = { cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28519" *) { in_dat_data109[7], in_dat_data_fp16_mts_sft54 };
  assign in_dat_data_fp16_53 = { cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28527" *) { in_dat_data107[7], in_dat_data_fp16_mts_sft53 };
  assign in_dat_data_fp16_52 = { cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28535" *) { in_dat_data105[7], in_dat_data_fp16_mts_sft52 };
  assign in_dat_data_fp16_51 = { cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28543" *) { in_dat_data103[7], in_dat_data_fp16_mts_sft51 };
  assign in_dat_data_fp16_50 = { cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28551" *) { in_dat_data101[7], in_dat_data_fp16_mts_sft50 };
  assign in_dat_data_fp16_49 = { cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28559" *) { in_dat_data99[7], in_dat_data_fp16_mts_sft49 };
  assign in_dat_data_fp16_48 = { cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28567" *) { in_dat_data97[7], in_dat_data_fp16_mts_sft48 };
  assign in_dat_data_fp16_47 = { cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28575" *) { in_dat_data95[7], in_dat_data_fp16_mts_sft47 };
  assign in_dat_data_fp16_46 = { cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28583" *) { in_dat_data93[7], in_dat_data_fp16_mts_sft46 };
  assign in_dat_data_fp16_45 = { cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28591" *) { in_dat_data91[7], in_dat_data_fp16_mts_sft45 };
  assign in_dat_data_fp16_44 = { cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28599" *) { in_dat_data89[7], in_dat_data_fp16_mts_sft44 };
  assign in_dat_data_fp16_43 = { cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28607" *) { in_dat_data87[7], in_dat_data_fp16_mts_sft43 };
  assign in_dat_data_fp16_42 = { cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28615" *) { in_dat_data85[7], in_dat_data_fp16_mts_sft42 };
  assign in_dat_data_fp16_41 = { cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28623" *) { in_dat_data83[7], in_dat_data_fp16_mts_sft41 };
  assign in_dat_data_fp16_40 = { cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28631" *) { in_dat_data81[7], in_dat_data_fp16_mts_sft40 };
  assign in_dat_data_fp16_39 = { cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28639" *) { in_dat_data79[7], in_dat_data_fp16_mts_sft39 };
  assign in_dat_data_fp16_38 = { cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28647" *) { in_dat_data77[7], in_dat_data_fp16_mts_sft38 };
  assign in_dat_data_fp16_37 = { cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28655" *) { in_dat_data75[7], in_dat_data_fp16_mts_sft37 };
  assign in_dat_data_fp16_36 = { cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28663" *) { in_dat_data73[7], in_dat_data_fp16_mts_sft36 };
  assign in_dat_data_fp16_35 = { cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28671" *) { in_dat_data71[7], in_dat_data_fp16_mts_sft35 };
  assign in_dat_data_fp16_34 = { cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28679" *) { in_dat_data69[7], in_dat_data_fp16_mts_sft34 };
  assign in_dat_data_fp16_33 = { cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28687" *) { in_dat_data67[7], in_dat_data_fp16_mts_sft33 };
  assign in_dat_data_fp16_32 = { cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28695" *) { in_dat_data65[7], in_dat_data_fp16_mts_sft32 };
  assign in_dat_data_fp16_31 = { cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28703" *) { in_dat_data63[7], in_dat_data_fp16_mts_sft31 };
  assign in_dat_data_fp16_30 = { cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28711" *) { in_dat_data61[7], in_dat_data_fp16_mts_sft30 };
  assign in_dat_data_fp16_29 = { cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28719" *) { in_dat_data59[7], in_dat_data_fp16_mts_sft29 };
  assign in_dat_data_fp16_28 = { cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28727" *) { in_dat_data57[7], in_dat_data_fp16_mts_sft28 };
  assign in_dat_data_fp16_27 = { cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28735" *) { in_dat_data55[7], in_dat_data_fp16_mts_sft27 };
  assign in_dat_data_fp16_26 = { cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28743" *) { in_dat_data53[7], in_dat_data_fp16_mts_sft26 };
  assign in_dat_data_fp16_25 = { cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28751" *) { in_dat_data51[7], in_dat_data_fp16_mts_sft25 };
  assign in_dat_data_fp16_24 = { cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28759" *) { in_dat_data49[7], in_dat_data_fp16_mts_sft24 };
  assign in_dat_data_fp16_23 = { cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28767" *) { in_dat_data47[7], in_dat_data_fp16_mts_sft23 };
  assign in_dat_data_fp16_22 = { cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28775" *) { in_dat_data45[7], in_dat_data_fp16_mts_sft22 };
  assign in_dat_data_fp16_21 = { cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28783" *) { in_dat_data43[7], in_dat_data_fp16_mts_sft21 };
  assign in_dat_data_fp16_20 = { cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28791" *) { in_dat_data41[7], in_dat_data_fp16_mts_sft20 };
  assign in_dat_data_fp16_19 = { cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28799" *) { in_dat_data39[7], in_dat_data_fp16_mts_sft19 };
  assign in_dat_data_fp16_18 = { cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28807" *) { in_dat_data37[7], in_dat_data_fp16_mts_sft18 };
  assign in_dat_data_fp16_17 = { cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28815" *) { in_dat_data35[7], in_dat_data_fp16_mts_sft17 };
  assign in_dat_data_fp16_16 = { cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28823" *) { in_dat_data33[7], in_dat_data_fp16_mts_sft16 };
  assign in_dat_data_fp16_15 = { cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28831" *) { in_dat_data31[7], in_dat_data_fp16_mts_sft15 };
  assign in_dat_data_fp16_14 = { cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28839" *) { in_dat_data29[7], in_dat_data_fp16_mts_sft14 };
  assign in_dat_data_fp16_13 = { cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28847" *) { in_dat_data27[7], in_dat_data_fp16_mts_sft13 };
  assign in_dat_data_fp16_12 = { cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28855" *) { in_dat_data25[7], in_dat_data_fp16_mts_sft12 };
  assign in_dat_data_fp16_11 = { cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28863" *) { in_dat_data23[7], in_dat_data_fp16_mts_sft11 };
  assign in_dat_data_fp16_10 = { cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28871" *) { in_dat_data21[7], in_dat_data_fp16_mts_sft10 };
  assign in_dat_data_fp16_9 = { cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28879" *) { in_dat_data19[7], in_dat_data_fp16_mts_sft9 };
  assign in_dat_data_fp16_8 = { cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28887" *) { in_dat_data17[7], in_dat_data_fp16_mts_sft8 };
  assign in_dat_data_fp16_7 = { cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28895" *) { in_dat_data15[7], in_dat_data_fp16_mts_sft7 };
  assign in_dat_data_fp16_6 = { cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28903" *) { in_dat_data13[7], in_dat_data_fp16_mts_sft6 };
  assign in_dat_data_fp16_5 = { cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28911" *) { in_dat_data11[7], in_dat_data_fp16_mts_sft5 };
  assign in_dat_data_fp16_4 = { cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28919" *) { in_dat_data9[7], in_dat_data_fp16_mts_sft4 };
  assign in_dat_data_fp16_3 = { cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28927" *) { in_dat_data7[7], in_dat_data_fp16_mts_sft3 };
  assign in_dat_data_fp16_2 = { cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28935" *) { in_dat_data5[7], in_dat_data_fp16_mts_sft2 };
  assign in_dat_data_fp16_1 = { cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28943" *) { in_dat_data3[7], in_dat_data_fp16_mts_sft1 };
  assign in_dat_data_fp16_0 = { cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28951" *) { in_dat_data1[7], in_dat_data_fp16_mts_sft0 };
  assign _05425_ = { _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_, _06407_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29041" *) in_dat_mask;
  assign _05426_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29076" *) cfg_is_fp16_d1[65];
  assign _05427_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29086" *) _07562_;
  assign _05428_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29096" *) _07563_;
  assign _05429_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29106" *) _07564_;
  assign _05430_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29116" *) _07565_;
  assign _05431_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29126" *) _07566_;
  assign _05432_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29136" *) _07567_;
  assign _05433_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29146" *) _07568_;
  assign _05434_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29156" *) _07569_;
  assign _05435_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29166" *) _07570_;
  assign _05436_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29176" *) _07571_;
  assign _05437_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29186" *) _07572_;
  assign _05438_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29196" *) _07573_;
  assign _05439_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29206" *) _07574_;
  assign _05440_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29216" *) _07575_;
  assign _05441_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29226" *) _07576_;
  assign _05442_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29236" *) _07577_;
  assign _05443_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29246" *) _07578_;
  assign _05444_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29256" *) _07579_;
  assign _05445_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29266" *) _07580_;
  assign _05446_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29276" *) _07581_;
  assign _05447_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29286" *) _07582_;
  assign _05448_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29296" *) _07583_;
  assign _05449_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29306" *) _07584_;
  assign _05450_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29316" *) _07585_;
  assign _05451_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29326" *) _07586_;
  assign _05452_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29336" *) _07587_;
  assign _05453_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29346" *) _07588_;
  assign _05454_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29356" *) _07589_;
  assign _05455_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29366" *) _07590_;
  assign _05456_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29376" *) _07591_;
  assign _05457_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29386" *) _07592_;
  assign _05458_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29396" *) _07593_;
  assign _05459_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29406" *) _07594_;
  assign _05460_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29416" *) _07595_;
  assign _05461_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29426" *) _07596_;
  assign _05462_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29436" *) _07597_;
  assign _05463_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29446" *) _07598_;
  assign _05464_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29456" *) _07599_;
  assign _05465_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29466" *) _07600_;
  assign _05466_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29476" *) _07601_;
  assign _05467_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29486" *) _07602_;
  assign _05468_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29496" *) _07603_;
  assign _05469_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29506" *) _07604_;
  assign _05470_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29516" *) _07605_;
  assign _05471_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29526" *) _07606_;
  assign _05472_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29536" *) _07607_;
  assign _05473_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29546" *) _07608_;
  assign _05474_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29556" *) _07609_;
  assign _05475_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29566" *) _07610_;
  assign _05476_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29576" *) _07611_;
  assign _05477_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29586" *) _07612_;
  assign _05478_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29596" *) _07613_;
  assign _05479_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29606" *) _07614_;
  assign _05480_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29616" *) _07615_;
  assign _05481_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29626" *) _07616_;
  assign _05482_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29636" *) _07617_;
  assign _05483_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29646" *) _07618_;
  assign _05484_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29656" *) _07619_;
  assign _05485_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29666" *) _07620_;
  assign _05486_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29676" *) _07621_;
  assign _05487_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29686" *) _07622_;
  assign _05488_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29696" *) _07623_;
  assign _05489_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29706" *) _07624_;
  assign _05490_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29716" *) _07625_;
  assign _05491_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29726" *) _07626_;
  assign _05492_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29736" *) _07627_;
  assign _05493_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29746" *) _07628_;
  assign _05494_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29756" *) _07629_;
  assign _05495_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29766" *) _07630_;
  assign _05496_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29776" *) _07631_;
  assign _05497_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29786" *) _07632_;
  assign _05498_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29796" *) _07633_;
  assign _05499_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29806" *) _07634_;
  assign _05500_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29816" *) _07635_;
  assign _05501_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29826" *) _07636_;
  assign _05502_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29836" *) _07637_;
  assign _05503_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29846" *) _07638_;
  assign _05504_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29856" *) _07639_;
  assign _05505_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29866" *) _07640_;
  assign _05506_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29876" *) _07641_;
  assign _05507_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29886" *) _07642_;
  assign _05508_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29896" *) _07643_;
  assign _05509_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29906" *) _07644_;
  assign _05510_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29916" *) _07645_;
  assign _05511_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29926" *) _07646_;
  assign _05512_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29936" *) _07647_;
  assign _05513_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29946" *) _07648_;
  assign _05514_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29956" *) _07649_;
  assign _05515_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29966" *) _07650_;
  assign _05516_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29976" *) _07651_;
  assign _05517_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29986" *) _07652_;
  assign _05518_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29996" *) _07653_;
  assign _05519_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30006" *) _07654_;
  assign _05520_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30016" *) _07655_;
  assign _05521_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30026" *) _07656_;
  assign _05522_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30036" *) _07657_;
  assign _05523_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30046" *) _07658_;
  assign _05524_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30056" *) _07659_;
  assign _05525_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30066" *) _07660_;
  assign _05526_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30076" *) _07661_;
  assign _05527_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30086" *) _07662_;
  assign _05528_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30096" *) _07663_;
  assign _05529_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30106" *) _07664_;
  assign _05530_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30116" *) _07665_;
  assign _05531_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30126" *) _07666_;
  assign _05532_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30136" *) _07667_;
  assign _05533_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30146" *) _07668_;
  assign _05534_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30156" *) _07669_;
  assign _05535_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30166" *) _07670_;
  assign _05536_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30176" *) _07671_;
  assign _05537_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30186" *) _07672_;
  assign _05538_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30196" *) _07673_;
  assign _05539_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30206" *) _07674_;
  assign _05540_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30216" *) _07675_;
  assign _05541_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30226" *) _07676_;
  assign _05542_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30236" *) _07677_;
  assign _05543_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30246" *) _07678_;
  assign _05544_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30256" *) _07679_;
  assign _05545_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30266" *) _07680_;
  assign _05546_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30276" *) _07681_;
  assign _05547_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30286" *) _07682_;
  assign _05548_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30296" *) _07683_;
  assign _05549_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30306" *) _07684_;
  assign _05550_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30316" *) _07685_;
  assign _05551_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30326" *) _07686_;
  assign _05552_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30336" *) _07687_;
  assign _05553_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30346" *) _07688_;
  assign _05554_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30356" *) _07689_;
  assign _01190_[15] = in_dat_stripe_st & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30369" *) in_dat_pvld;
  assign _01189_[8] = in_dat_stripe_end & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30376" *) in_dat_pvld;
  assign _05555_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30380" *) cfg_is_fp16_d1[82];
  assign _05556_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30400" *) cfg_is_fp16_d1[83];
  assign _05557_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30420" *) cfg_is_fp16_d1[84];
  assign _05558_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30440" *) cfg_is_fp16_d1[85];
  assign _05559_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30460" *) cfg_is_fp16_d1[86];
  assign _05560_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30480" *) cfg_is_fp16_d1[87];
  assign _05561_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30500" *) cfg_is_fp16_d1[88];
  assign _05562_ = in_dat_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30520" *) cfg_is_fp16_d1[89];
  assign _05563_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30664" *) cfg_is_fp16_d1[90];
  assign _05564_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30674" *) _07690_;
  assign _05565_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30684" *) _07691_;
  assign _05566_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30694" *) _07692_;
  assign _05567_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30704" *) _07693_;
  assign _05568_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30714" *) _07694_;
  assign _05569_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30724" *) _07695_;
  assign _05570_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30734" *) _07696_;
  assign _05571_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30744" *) _07697_;
  assign _05572_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30754" *) _07698_;
  assign _05573_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30764" *) _07699_;
  assign _05574_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30774" *) _07700_;
  assign _05575_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30784" *) _07701_;
  assign _05576_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30794" *) _07702_;
  assign _05577_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30804" *) _07703_;
  assign _05578_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30814" *) _07704_;
  assign _05579_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30824" *) _07705_;
  assign _05580_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30834" *) _07706_;
  assign _05581_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30844" *) _07707_;
  assign _05582_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30854" *) _07708_;
  assign _05583_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30864" *) _07709_;
  assign _05584_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30874" *) _07710_;
  assign _05585_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30884" *) _07711_;
  assign _05586_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30894" *) _07712_;
  assign _05587_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30904" *) _07713_;
  assign _05588_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30914" *) _07714_;
  assign _05589_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30924" *) _07715_;
  assign _05590_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30934" *) _07716_;
  assign _05591_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30944" *) _07717_;
  assign _05592_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30954" *) _07718_;
  assign _05593_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30964" *) _07719_;
  assign _05594_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30974" *) _07720_;
  assign _05595_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30984" *) _07721_;
  assign _05596_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30994" *) _07722_;
  assign _05597_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31004" *) _07723_;
  assign _05598_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31014" *) _07724_;
  assign _05599_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31024" *) _07725_;
  assign _05600_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31034" *) _07726_;
  assign _05601_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31044" *) _07727_;
  assign _05602_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31054" *) _07728_;
  assign _05603_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31064" *) _07729_;
  assign _05604_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31074" *) _07730_;
  assign _05605_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31084" *) _07731_;
  assign _05606_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31094" *) _07732_;
  assign _05607_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31104" *) _07733_;
  assign _05608_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31114" *) _07734_;
  assign _05609_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31124" *) _07735_;
  assign _05610_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31134" *) _07736_;
  assign _05611_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31144" *) _07737_;
  assign _05612_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31154" *) _07738_;
  assign _05613_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31164" *) _07739_;
  assign _05614_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31174" *) _07740_;
  assign _05615_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31184" *) _07741_;
  assign _05616_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31194" *) _07742_;
  assign _05617_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31204" *) _07743_;
  assign _05618_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31214" *) _07744_;
  assign _05619_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31224" *) _07745_;
  assign _05620_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31234" *) _07746_;
  assign _05621_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31244" *) _07747_;
  assign _05622_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31254" *) _07748_;
  assign _05623_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31264" *) _07749_;
  assign _05624_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31274" *) _07750_;
  assign _05625_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31284" *) _07751_;
  assign _05626_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31294" *) _07752_;
  assign _05627_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31304" *) _07753_;
  assign _05628_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31314" *) _07754_;
  assign _05629_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31324" *) _07755_;
  assign _05630_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31334" *) _07756_;
  assign _05631_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31344" *) _07757_;
  assign _05632_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31354" *) _07758_;
  assign _05633_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31364" *) _07759_;
  assign _05634_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31374" *) _07760_;
  assign _05635_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31384" *) _07761_;
  assign _05636_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31394" *) _07762_;
  assign _05637_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31404" *) _07763_;
  assign _05638_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31414" *) _07764_;
  assign _05639_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31424" *) _07765_;
  assign _05640_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31434" *) _07766_;
  assign _05641_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31444" *) _07767_;
  assign _05642_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31454" *) _07768_;
  assign _05643_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31464" *) _07769_;
  assign _05644_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31474" *) _07770_;
  assign _05645_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31484" *) _07771_;
  assign _05646_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31494" *) _07772_;
  assign _05647_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31504" *) _07773_;
  assign _05648_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31514" *) _07774_;
  assign _05649_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31524" *) _07775_;
  assign _05650_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31534" *) _07776_;
  assign _05651_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31544" *) _07777_;
  assign _05652_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31554" *) _07778_;
  assign _05653_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31564" *) _07779_;
  assign _05654_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31574" *) _07780_;
  assign _05655_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31584" *) _07781_;
  assign _05656_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31594" *) _07782_;
  assign _05657_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31604" *) _07783_;
  assign _05658_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31614" *) _07784_;
  assign _05659_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31624" *) _07785_;
  assign _05660_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31634" *) _07786_;
  assign _05661_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31644" *) _07787_;
  assign _05662_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31654" *) _07788_;
  assign _05663_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31664" *) _07789_;
  assign _05664_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31674" *) _07790_;
  assign _05665_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31684" *) _07791_;
  assign _05666_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31694" *) _07792_;
  assign _05667_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31704" *) _07793_;
  assign _05668_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31714" *) _07794_;
  assign _05669_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31724" *) _07795_;
  assign _05670_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31734" *) _07796_;
  assign _05671_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31744" *) _07797_;
  assign _05672_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31754" *) _07798_;
  assign _05673_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31764" *) _07799_;
  assign _05674_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31774" *) _07800_;
  assign _05675_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31784" *) _07801_;
  assign _05676_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31794" *) _07802_;
  assign _05677_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31804" *) _07803_;
  assign _05678_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31814" *) _07804_;
  assign _05679_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31824" *) _07805_;
  assign _05680_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31834" *) _07806_;
  assign _05681_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31844" *) _07807_;
  assign _05682_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31854" *) _07808_;
  assign _05683_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31864" *) _07809_;
  assign _05684_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31874" *) _07810_;
  assign _05685_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31884" *) _07811_;
  assign _05686_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31894" *) _07812_;
  assign _05687_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31904" *) _07813_;
  assign _05688_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31914" *) _07814_;
  assign _05689_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31924" *) _07815_;
  assign _05690_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31934" *) _07816_;
  assign _05691_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31944" *) _07817_;
  assign _05692_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31971" *) cfg_is_fp16_d1[91];
  assign _05693_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33278" *) cfg_is_fp16_d1[92];
  assign in_wt_data_fp16_63 = { cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63], cfg_is_fp16_d1[63] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3374" *) { in_wt_data127[7], in_wt_data_fp16_mts_sft63 };
  assign in_wt_data_fp16_62 = { cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62], cfg_is_fp16_d1[62] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3382" *) { in_wt_data125[7], in_wt_data_fp16_mts_sft62 };
  assign in_wt_data_fp16_61 = { cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61], cfg_is_fp16_d1[61] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3390" *) { in_wt_data123[7], in_wt_data_fp16_mts_sft61 };
  assign in_wt_data_fp16_60 = { cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60], cfg_is_fp16_d1[60] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3398" *) { in_wt_data121[7], in_wt_data_fp16_mts_sft60 };
  assign in_wt_data_fp16_59 = { cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59], cfg_is_fp16_d1[59] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3406" *) { in_wt_data119[7], in_wt_data_fp16_mts_sft59 };
  assign in_wt_data_fp16_58 = { cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58], cfg_is_fp16_d1[58] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3414" *) { in_wt_data117[7], in_wt_data_fp16_mts_sft58 };
  assign in_wt_data_fp16_57 = { cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57], cfg_is_fp16_d1[57] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3422" *) { in_wt_data115[7], in_wt_data_fp16_mts_sft57 };
  assign in_wt_data_fp16_56 = { cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56], cfg_is_fp16_d1[56] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3430" *) { in_wt_data113[7], in_wt_data_fp16_mts_sft56 };
  assign in_wt_data_fp16_55 = { cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55], cfg_is_fp16_d1[55] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3438" *) { in_wt_data111[7], in_wt_data_fp16_mts_sft55 };
  assign in_wt_data_fp16_54 = { cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54], cfg_is_fp16_d1[54] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3446" *) { in_wt_data109[7], in_wt_data_fp16_mts_sft54 };
  assign in_wt_data_fp16_53 = { cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53], cfg_is_fp16_d1[53] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3454" *) { in_wt_data107[7], in_wt_data_fp16_mts_sft53 };
  assign _05694_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34585" *) cfg_is_fp16_d1[93];
  assign in_wt_data_fp16_52 = { cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52], cfg_is_fp16_d1[52] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3462" *) { in_wt_data105[7], in_wt_data_fp16_mts_sft52 };
  assign in_wt_data_fp16_51 = { cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51], cfg_is_fp16_d1[51] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3470" *) { in_wt_data103[7], in_wt_data_fp16_mts_sft51 };
  assign in_wt_data_fp16_50 = { cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50], cfg_is_fp16_d1[50] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3478" *) { in_wt_data101[7], in_wt_data_fp16_mts_sft50 };
  assign in_wt_data_fp16_49 = { cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49], cfg_is_fp16_d1[49] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3486" *) { in_wt_data99[7], in_wt_data_fp16_mts_sft49 };
  assign in_wt_data_fp16_48 = { cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48], cfg_is_fp16_d1[48] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3494" *) { in_wt_data97[7], in_wt_data_fp16_mts_sft48 };
  assign in_wt_data_fp16_47 = { cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47], cfg_is_fp16_d1[47] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3502" *) { in_wt_data95[7], in_wt_data_fp16_mts_sft47 };
  assign in_wt_data_fp16_46 = { cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46], cfg_is_fp16_d1[46] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3510" *) { in_wt_data93[7], in_wt_data_fp16_mts_sft46 };
  assign in_wt_data_fp16_45 = { cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45], cfg_is_fp16_d1[45] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3518" *) { in_wt_data91[7], in_wt_data_fp16_mts_sft45 };
  assign in_wt_data_fp16_44 = { cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44], cfg_is_fp16_d1[44] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3526" *) { in_wt_data89[7], in_wt_data_fp16_mts_sft44 };
  assign in_wt_data_fp16_43 = { cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43], cfg_is_fp16_d1[43] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3534" *) { in_wt_data87[7], in_wt_data_fp16_mts_sft43 };
  assign in_wt_data_fp16_42 = { cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42], cfg_is_fp16_d1[42] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3542" *) { in_wt_data85[7], in_wt_data_fp16_mts_sft42 };
  assign in_wt_data_fp16_41 = { cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41], cfg_is_fp16_d1[41] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3550" *) { in_wt_data83[7], in_wt_data_fp16_mts_sft41 };
  assign in_wt_data_fp16_40 = { cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40], cfg_is_fp16_d1[40] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3558" *) { in_wt_data81[7], in_wt_data_fp16_mts_sft40 };
  assign in_wt_data_fp16_39 = { cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39], cfg_is_fp16_d1[39] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3566" *) { in_wt_data79[7], in_wt_data_fp16_mts_sft39 };
  assign in_wt_data_fp16_38 = { cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38], cfg_is_fp16_d1[38] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3574" *) { in_wt_data77[7], in_wt_data_fp16_mts_sft38 };
  assign in_wt_data_fp16_37 = { cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37], cfg_is_fp16_d1[37] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3582" *) { in_wt_data75[7], in_wt_data_fp16_mts_sft37 };
  assign _05695_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35892" *) cfg_is_fp16_d1[94];
  assign in_wt_data_fp16_36 = { cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36], cfg_is_fp16_d1[36] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3590" *) { in_wt_data73[7], in_wt_data_fp16_mts_sft36 };
  assign in_wt_data_fp16_35 = { cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35], cfg_is_fp16_d1[35] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3598" *) { in_wt_data71[7], in_wt_data_fp16_mts_sft35 };
  assign in_wt_data_fp16_34 = { cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34], cfg_is_fp16_d1[34] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3606" *) { in_wt_data69[7], in_wt_data_fp16_mts_sft34 };
  assign in_wt_data_fp16_33 = { cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33], cfg_is_fp16_d1[33] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3614" *) { in_wt_data67[7], in_wt_data_fp16_mts_sft33 };
  assign in_wt_data_fp16_32 = { cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32], cfg_is_fp16_d1[32] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3622" *) { in_wt_data65[7], in_wt_data_fp16_mts_sft32 };
  assign in_wt_data_fp16_31 = { cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31], cfg_is_fp16_d1[31] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3630" *) { in_wt_data63[7], in_wt_data_fp16_mts_sft31 };
  assign in_wt_data_fp16_30 = { cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30], cfg_is_fp16_d1[30] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3638" *) { in_wt_data61[7], in_wt_data_fp16_mts_sft30 };
  assign in_wt_data_fp16_29 = { cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29], cfg_is_fp16_d1[29] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3646" *) { in_wt_data59[7], in_wt_data_fp16_mts_sft29 };
  assign in_wt_data_fp16_28 = { cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28], cfg_is_fp16_d1[28] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3654" *) { in_wt_data57[7], in_wt_data_fp16_mts_sft28 };
  assign in_wt_data_fp16_27 = { cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27], cfg_is_fp16_d1[27] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3662" *) { in_wt_data55[7], in_wt_data_fp16_mts_sft27 };
  assign in_wt_data_fp16_26 = { cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26], cfg_is_fp16_d1[26] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3670" *) { in_wt_data53[7], in_wt_data_fp16_mts_sft26 };
  assign in_wt_data_fp16_25 = { cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25], cfg_is_fp16_d1[25] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3678" *) { in_wt_data51[7], in_wt_data_fp16_mts_sft25 };
  assign in_wt_data_fp16_24 = { cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24], cfg_is_fp16_d1[24] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3686" *) { in_wt_data49[7], in_wt_data_fp16_mts_sft24 };
  assign in_wt_data_fp16_23 = { cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23], cfg_is_fp16_d1[23] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3694" *) { in_wt_data47[7], in_wt_data_fp16_mts_sft23 };
  assign in_wt_data_fp16_22 = { cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22], cfg_is_fp16_d1[22] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3702" *) { in_wt_data45[7], in_wt_data_fp16_mts_sft22 };
  assign in_wt_data_fp16_21 = { cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21], cfg_is_fp16_d1[21] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3710" *) { in_wt_data43[7], in_wt_data_fp16_mts_sft21 };
  assign in_wt_data_fp16_20 = { cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20], cfg_is_fp16_d1[20] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3718" *) { in_wt_data41[7], in_wt_data_fp16_mts_sft20 };
  assign _05696_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37199" *) cfg_is_fp16_d1[95];
  assign in_wt_data_fp16_19 = { cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19], cfg_is_fp16_d1[19] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3726" *) { in_wt_data39[7], in_wt_data_fp16_mts_sft19 };
  assign in_wt_data_fp16_18 = { cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18], cfg_is_fp16_d1[18] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3734" *) { in_wt_data37[7], in_wt_data_fp16_mts_sft18 };
  assign in_wt_data_fp16_17 = { cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17], cfg_is_fp16_d1[17] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3742" *) { in_wt_data35[7], in_wt_data_fp16_mts_sft17 };
  assign in_wt_data_fp16_16 = { cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16], cfg_is_fp16_d1[16] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3750" *) { in_wt_data33[7], in_wt_data_fp16_mts_sft16 };
  assign in_wt_data_fp16_15 = { cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15], cfg_is_fp16_d1[15] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3758" *) { in_wt_data31[7], in_wt_data_fp16_mts_sft15 };
  assign in_wt_data_fp16_14 = { cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14], cfg_is_fp16_d1[14] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3766" *) { in_wt_data29[7], in_wt_data_fp16_mts_sft14 };
  assign in_wt_data_fp16_13 = { cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13], cfg_is_fp16_d1[13] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3774" *) { in_wt_data27[7], in_wt_data_fp16_mts_sft13 };
  assign in_wt_data_fp16_12 = { cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12], cfg_is_fp16_d1[12] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3782" *) { in_wt_data25[7], in_wt_data_fp16_mts_sft12 };
  assign in_wt_data_fp16_11 = { cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11], cfg_is_fp16_d1[11] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3790" *) { in_wt_data23[7], in_wt_data_fp16_mts_sft11 };
  assign in_wt_data_fp16_10 = { cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10], cfg_is_fp16_d1[10] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3798" *) { in_wt_data21[7], in_wt_data_fp16_mts_sft10 };
  assign in_wt_data_fp16_9 = { cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9], cfg_is_fp16_d1[9] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3806" *) { in_wt_data19[7], in_wt_data_fp16_mts_sft9 };
  assign in_wt_data_fp16_8 = { cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8], cfg_is_fp16_d1[8] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3814" *) { in_wt_data17[7], in_wt_data_fp16_mts_sft8 };
  assign in_wt_data_fp16_7 = { cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7], cfg_is_fp16_d1[7] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3822" *) { in_wt_data15[7], in_wt_data_fp16_mts_sft7 };
  assign in_wt_data_fp16_6 = { cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6], cfg_is_fp16_d1[6] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3830" *) { in_wt_data13[7], in_wt_data_fp16_mts_sft6 };
  assign in_wt_data_fp16_5 = { cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5], cfg_is_fp16_d1[5] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3838" *) { in_wt_data11[7], in_wt_data_fp16_mts_sft5 };
  assign in_wt_data_fp16_4 = { cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4], cfg_is_fp16_d1[4] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3846" *) { in_wt_data9[7], in_wt_data_fp16_mts_sft4 };
  assign _05697_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38506" *) cfg_is_fp16_d1[96];
  assign in_wt_data_fp16_3 = { cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3], cfg_is_fp16_d1[3] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3854" *) { in_wt_data7[7], in_wt_data_fp16_mts_sft3 };
  assign in_wt_data_fp16_2 = { cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2], cfg_is_fp16_d1[2] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3862" *) { in_wt_data5[7], in_wt_data_fp16_mts_sft2 };
  assign in_wt_data_fp16_1 = { cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1], cfg_is_fp16_d1[1] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3870" *) { in_wt_data3[7], in_wt_data_fp16_mts_sft1 };
  assign in_wt_data_fp16_0 = { cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0], cfg_is_fp16_d1[0] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3878" *) { in_wt_data1[7], in_wt_data_fp16_mts_sft0 };
  assign _05698_ = { _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_, _06408_ } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3968" *) in_wt_mask;
  assign _05699_ = dat_pre_pvld[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39813" *) cfg_is_fp16_d1[97];
  assign _05700_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4003" *) cfg_is_fp16_d1[65];
  assign _05701_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4033" *) _07819_;
  assign _05702_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4043" *) _07820_;
  assign _05703_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4053" *) _07821_;
  assign _05704_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4063" *) _07822_;
  assign _05705_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4073" *) _07823_;
  assign _05706_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4083" *) _07824_;
  assign _05707_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4093" *) _07825_;
  assign _05708_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4103" *) _07826_;
  assign _05709_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4113" *) _07827_;
  assign _05710_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4123" *) _07828_;
  assign _05711_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4133" *) _07829_;
  assign _05712_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4143" *) _07830_;
  assign _05713_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4153" *) _07831_;
  assign _05714_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4163" *) _07832_;
  assign _05715_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4173" *) _07833_;
  assign _05716_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4183" *) _07834_;
  assign _05717_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4193" *) _07835_;
  assign _05718_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4203" *) _07836_;
  assign _05719_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4213" *) _07837_;
  assign _05720_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4223" *) _07838_;
  assign _05721_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4233" *) _07839_;
  assign _05722_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4243" *) _07840_;
  assign _05723_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4253" *) _07841_;
  assign _05724_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4263" *) _07842_;
  assign _05725_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4273" *) _07843_;
  assign _05726_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4283" *) _07844_;
  assign _05727_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4293" *) _07845_;
  assign _05728_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4303" *) _07846_;
  assign _05729_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4313" *) _07847_;
  assign _05730_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4323" *) _07848_;
  assign _05731_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4333" *) _07849_;
  assign _05732_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4343" *) _07850_;
  assign _05733_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4353" *) _07851_;
  assign _05734_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4363" *) _07852_;
  assign _05735_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4373" *) _07853_;
  assign _05736_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4383" *) _07854_;
  assign _05737_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4393" *) _07855_;
  assign _05738_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4403" *) _07856_;
  assign _05739_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4413" *) _07857_;
  assign _05740_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4423" *) _07858_;
  assign _05741_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4433" *) _07859_;
  assign _05742_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4443" *) _07860_;
  assign _05743_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4453" *) _07861_;
  assign _05744_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4463" *) _07862_;
  assign _05745_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4473" *) _07863_;
  assign _05746_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4483" *) _07864_;
  assign _05747_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4493" *) _07865_;
  assign _05748_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4503" *) _07866_;
  assign _05749_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4513" *) _07867_;
  assign _05750_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4523" *) _07868_;
  assign _05751_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4533" *) _07869_;
  assign _05752_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4543" *) _07870_;
  assign _05753_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4553" *) _07871_;
  assign _05754_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4563" *) _07872_;
  assign _05755_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4573" *) _07873_;
  assign _05756_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4583" *) _07874_;
  assign _05757_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4593" *) _07875_;
  assign _05758_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4603" *) _07876_;
  assign _05759_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4613" *) _07877_;
  assign _05760_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4623" *) _07878_;
  assign _05761_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4633" *) _07879_;
  assign _05762_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4643" *) _07880_;
  assign _05763_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4653" *) _07881_;
  assign _05764_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4663" *) _07882_;
  assign _05765_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4673" *) _07883_;
  assign _05766_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4683" *) _07884_;
  assign _05767_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4693" *) _07885_;
  assign _05768_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4703" *) _07886_;
  assign _05769_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4713" *) _07887_;
  assign _05770_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4723" *) _07888_;
  assign _05771_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4733" *) _07889_;
  assign _05772_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4743" *) _07890_;
  assign _05773_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4753" *) _07891_;
  assign _05774_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4763" *) _07892_;
  assign _05775_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4773" *) _07893_;
  assign _05776_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4783" *) _07894_;
  assign _05777_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4793" *) _07895_;
  assign _05778_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4803" *) _07896_;
  assign _05779_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4813" *) _07897_;
  assign _05780_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4823" *) _07898_;
  assign _05781_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4833" *) _07899_;
  assign _05782_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4843" *) _07900_;
  assign _05783_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4853" *) _07901_;
  assign _05784_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4863" *) _07902_;
  assign _05785_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4873" *) _07903_;
  assign _05786_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4883" *) _07904_;
  assign _05787_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4893" *) _07905_;
  assign _05788_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4903" *) _07906_;
  assign _05789_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4913" *) _07907_;
  assign _05790_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4923" *) _07908_;
  assign _05791_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4933" *) _07909_;
  assign _05792_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4943" *) _07910_;
  assign _05793_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4953" *) _07911_;
  assign _05794_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4963" *) _07912_;
  assign _05795_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4973" *) _07913_;
  assign _05796_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4983" *) _07914_;
  assign _05797_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4993" *) _07915_;
  assign _05798_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5003" *) _07916_;
  assign _05799_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5013" *) _07917_;
  assign _05800_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5023" *) _07918_;
  assign _05801_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5033" *) _07919_;
  assign _05802_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5043" *) _07920_;
  assign _05803_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5053" *) _07921_;
  assign _05804_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5063" *) _07922_;
  assign _05805_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5073" *) _07923_;
  assign _05806_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5083" *) _07924_;
  assign _05807_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5093" *) _07925_;
  assign _05808_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5103" *) _07926_;
  assign _05809_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5113" *) _07927_;
  assign _05810_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5123" *) _07928_;
  assign _05811_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5133" *) _07929_;
  assign _05812_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5143" *) _07930_;
  assign _05813_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5153" *) _07931_;
  assign _05814_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5163" *) _07932_;
  assign _05815_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5173" *) _07933_;
  assign _05816_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5183" *) _07934_;
  assign _05817_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5193" *) _07935_;
  assign _05818_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5203" *) _07936_;
  assign _05819_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5213" *) _07937_;
  assign _05820_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5223" *) _07938_;
  assign _05821_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5233" *) _07939_;
  assign _05822_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5243" *) _07940_;
  assign _05823_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5253" *) _07941_;
  assign _05824_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5263" *) _07942_;
  assign _05825_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5273" *) _07943_;
  assign _05826_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5283" *) _07944_;
  assign _05827_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5293" *) _07945_;
  assign _05828_ = in_wt_pvld & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5303" *) _07946_;
  assign _05829_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5342" *) cfg_is_fp16_d1[66];
  assign _05830_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5372" *) _06475_;
  assign _05831_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5382" *) _06476_;
  assign _05832_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5392" *) _06477_;
  assign _05833_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5402" *) _06478_;
  assign _05834_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5412" *) _06479_;
  assign _05835_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5422" *) _06480_;
  assign _05836_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5432" *) _06481_;
  assign _05837_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5442" *) _06482_;
  assign _05838_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5452" *) _06483_;
  assign _05839_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5462" *) _06484_;
  assign _05840_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5472" *) _06485_;
  assign _05841_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5482" *) _06486_;
  assign _05842_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5492" *) _06487_;
  assign _05843_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5502" *) _06488_;
  assign _05844_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5512" *) _06489_;
  assign _05845_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5522" *) _06490_;
  assign _05846_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5532" *) _06491_;
  assign _05847_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5542" *) _06492_;
  assign _05848_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5552" *) _06493_;
  assign _05849_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5562" *) _06494_;
  assign _05850_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5572" *) _06495_;
  assign _05851_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5582" *) _06496_;
  assign _05852_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5592" *) _06497_;
  assign _05853_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5602" *) _06498_;
  assign _05854_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5612" *) _06499_;
  assign _05855_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5622" *) _06500_;
  assign _05856_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5632" *) _06501_;
  assign _05857_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5642" *) _06502_;
  assign _05858_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5652" *) _06503_;
  assign _05859_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5662" *) _06504_;
  assign _05860_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5672" *) _06505_;
  assign _05861_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5682" *) _06506_;
  assign _05862_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5692" *) _06507_;
  assign _05863_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5702" *) _06508_;
  assign _05864_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5712" *) _06509_;
  assign _05865_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5722" *) _06510_;
  assign _05866_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5732" *) _06511_;
  assign _05867_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5742" *) _06512_;
  assign _05868_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5752" *) _06513_;
  assign _05869_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5762" *) _06514_;
  assign _05870_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5772" *) _06515_;
  assign _05871_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5782" *) _06516_;
  assign _05872_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5792" *) _06517_;
  assign _05873_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5802" *) _06518_;
  assign _05874_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5812" *) _06519_;
  assign _05875_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5822" *) _06520_;
  assign _05876_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5832" *) _06521_;
  assign _05877_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5842" *) _06522_;
  assign _05878_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5852" *) _06523_;
  assign _05879_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5862" *) _06524_;
  assign _05880_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5872" *) _06525_;
  assign _05881_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5882" *) _06526_;
  assign _05882_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5892" *) _06527_;
  assign _05883_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5902" *) _06528_;
  assign _05884_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5912" *) _06529_;
  assign _05885_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5922" *) _06530_;
  assign _05886_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5932" *) _06531_;
  assign _05887_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5942" *) _06532_;
  assign _05888_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5952" *) _06533_;
  assign _05889_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5962" *) _06534_;
  assign _05890_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5972" *) _06535_;
  assign _05891_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5982" *) _06536_;
  assign _05892_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5992" *) _06409_;
  assign _05893_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6002" *) _06410_;
  assign _05894_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6012" *) _06411_;
  assign _05895_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6022" *) _06412_;
  assign _05896_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6032" *) _06413_;
  assign _05897_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6042" *) _06414_;
  assign _05898_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6052" *) _06415_;
  assign _05899_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6062" *) _06416_;
  assign _05900_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6072" *) _06417_;
  assign _05901_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6082" *) _06418_;
  assign _05902_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6092" *) _06419_;
  assign _05903_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6102" *) _06420_;
  assign _05904_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6112" *) _06421_;
  assign _05905_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6122" *) _06422_;
  assign _05906_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6132" *) _06423_;
  assign _05907_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6142" *) _06424_;
  assign _05908_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6152" *) _06425_;
  assign _05909_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6162" *) _06426_;
  assign _05910_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6172" *) _06427_;
  assign _05911_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6182" *) _06428_;
  assign _05912_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6192" *) _06429_;
  assign _05913_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6202" *) _06430_;
  assign _05914_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6212" *) _06431_;
  assign _05915_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6222" *) _06432_;
  assign _05916_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6232" *) _06433_;
  assign _05917_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6242" *) _06434_;
  assign _05918_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6252" *) _06435_;
  assign _05919_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6262" *) _06436_;
  assign _05920_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6272" *) _06437_;
  assign _05921_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6282" *) _06438_;
  assign _05922_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6292" *) _06439_;
  assign _05923_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6302" *) _06440_;
  assign _05924_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6312" *) _06441_;
  assign _05925_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6322" *) _06442_;
  assign _05926_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6332" *) _06443_;
  assign _05927_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6342" *) _06444_;
  assign _05928_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6352" *) _06445_;
  assign _05929_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6362" *) _06446_;
  assign _05930_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6372" *) _06447_;
  assign _05931_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6382" *) _06448_;
  assign _05932_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6392" *) _06449_;
  assign _05933_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6402" *) _06450_;
  assign _05934_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6412" *) _06451_;
  assign _05935_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6422" *) _06452_;
  assign _05936_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6432" *) _06453_;
  assign _05937_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6442" *) _06454_;
  assign _05938_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6452" *) _06455_;
  assign _05939_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6462" *) _06456_;
  assign _05940_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6472" *) _06457_;
  assign _05941_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6482" *) _06458_;
  assign _05942_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6492" *) _06459_;
  assign _05943_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6502" *) _06460_;
  assign _05944_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6512" *) _06461_;
  assign _05945_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6522" *) _06462_;
  assign _05946_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6532" *) _06463_;
  assign _05947_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6542" *) _06464_;
  assign _05948_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6552" *) _06465_;
  assign _05949_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6562" *) _06466_;
  assign _05950_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6572" *) _06467_;
  assign _05951_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6582" *) _06468_;
  assign _05952_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6592" *) _06469_;
  assign _05953_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6602" *) _06470_;
  assign _05954_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6612" *) _06471_;
  assign _05955_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6622" *) _06472_;
  assign _05956_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6632" *) _06473_;
  assign _05957_ = wt_pre_sel[0] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6642" *) _06474_;
  assign _05958_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6678" *) cfg_is_fp16_d1[67];
  assign _05959_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6708" *) _06475_;
  assign _05960_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6718" *) _06476_;
  assign _05961_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6728" *) _06477_;
  assign _05962_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6738" *) _06478_;
  assign _05963_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6748" *) _06479_;
  assign _05964_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6758" *) _06480_;
  assign _05965_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6768" *) _06481_;
  assign _05966_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6778" *) _06482_;
  assign _05967_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6788" *) _06483_;
  assign _05968_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6798" *) _06484_;
  assign _05969_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6808" *) _06485_;
  assign _05970_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6818" *) _06486_;
  assign _05971_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6828" *) _06487_;
  assign _05972_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6838" *) _06488_;
  assign _05973_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6848" *) _06489_;
  assign _05974_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6858" *) _06490_;
  assign _05975_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6868" *) _06491_;
  assign _05976_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6878" *) _06492_;
  assign _05977_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6888" *) _06493_;
  assign _05978_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6898" *) _06494_;
  assign _05979_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6908" *) _06495_;
  assign _05980_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6918" *) _06496_;
  assign _05981_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6928" *) _06497_;
  assign _05982_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6938" *) _06498_;
  assign _05983_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6948" *) _06499_;
  assign _05984_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6958" *) _06500_;
  assign _05985_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6968" *) _06501_;
  assign _05986_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6978" *) _06502_;
  assign _05987_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6988" *) _06503_;
  assign _05988_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6998" *) _06504_;
  assign _05989_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7008" *) _06505_;
  assign _05990_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7018" *) _06506_;
  assign _05991_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7028" *) _06507_;
  assign _05992_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7038" *) _06508_;
  assign _05993_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7048" *) _06509_;
  assign _05994_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7058" *) _06510_;
  assign _05995_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7068" *) _06511_;
  assign _05996_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7078" *) _06512_;
  assign _05997_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7088" *) _06513_;
  assign _05998_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7098" *) _06514_;
  assign _05999_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7108" *) _06515_;
  assign _06000_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7118" *) _06516_;
  assign _06001_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7128" *) _06517_;
  assign _06002_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7138" *) _06518_;
  assign _06003_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7148" *) _06519_;
  assign _06004_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7158" *) _06520_;
  assign _06005_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7168" *) _06521_;
  assign _06006_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7178" *) _06522_;
  assign _06007_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7188" *) _06523_;
  assign _06008_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7198" *) _06524_;
  assign _06009_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7208" *) _06525_;
  assign _06010_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7218" *) _06526_;
  assign _06011_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7228" *) _06527_;
  assign _06012_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7238" *) _06528_;
  assign _06013_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7248" *) _06529_;
  assign _06014_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7258" *) _06530_;
  assign _06015_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7268" *) _06531_;
  assign _06016_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7278" *) _06532_;
  assign _06017_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7288" *) _06533_;
  assign _06018_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7298" *) _06534_;
  assign _06019_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7308" *) _06535_;
  assign _06020_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7318" *) _06536_;
  assign _06021_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7328" *) _06409_;
  assign _06022_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7338" *) _06410_;
  assign _06023_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7348" *) _06411_;
  assign _06024_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7358" *) _06412_;
  assign _06025_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7368" *) _06413_;
  assign _06026_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7378" *) _06414_;
  assign _06027_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7388" *) _06415_;
  assign _06028_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7398" *) _06416_;
  assign _06029_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7408" *) _06417_;
  assign _06030_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7418" *) _06418_;
  assign _06031_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7428" *) _06419_;
  assign _06032_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7438" *) _06420_;
  assign _06033_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7448" *) _06421_;
  assign _06034_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7458" *) _06422_;
  assign _06035_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7468" *) _06423_;
  assign _06036_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7478" *) _06424_;
  assign _06037_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7488" *) _06425_;
  assign _06038_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7498" *) _06426_;
  assign _06039_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7508" *) _06427_;
  assign _06040_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7518" *) _06428_;
  assign _06041_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7528" *) _06429_;
  assign _06042_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7538" *) _06430_;
  assign _06043_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7548" *) _06431_;
  assign _06044_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7558" *) _06432_;
  assign _06045_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7568" *) _06433_;
  assign _06046_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7578" *) _06434_;
  assign _06047_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7588" *) _06435_;
  assign _06048_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7598" *) _06436_;
  assign _06049_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7608" *) _06437_;
  assign _06050_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7618" *) _06438_;
  assign _06051_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7628" *) _06439_;
  assign _06052_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7638" *) _06440_;
  assign _06053_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7648" *) _06441_;
  assign _06054_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7658" *) _06442_;
  assign _06055_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7668" *) _06443_;
  assign _06056_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7678" *) _06444_;
  assign _06057_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7688" *) _06445_;
  assign _06058_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7698" *) _06446_;
  assign _06059_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7708" *) _06447_;
  assign _06060_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7718" *) _06448_;
  assign _06061_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7728" *) _06449_;
  assign _06062_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7738" *) _06450_;
  assign _06063_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7748" *) _06451_;
  assign _06064_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7758" *) _06452_;
  assign _06065_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7768" *) _06453_;
  assign _06066_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7778" *) _06454_;
  assign _06067_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7788" *) _06455_;
  assign _06068_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7798" *) _06456_;
  assign _06069_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7808" *) _06457_;
  assign _06070_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7818" *) _06458_;
  assign _06071_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7828" *) _06459_;
  assign _06072_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7838" *) _06460_;
  assign _06073_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7848" *) _06461_;
  assign _06074_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7858" *) _06462_;
  assign _06075_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7868" *) _06463_;
  assign _06076_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7878" *) _06464_;
  assign _06077_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7888" *) _06465_;
  assign _06078_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7898" *) _06466_;
  assign _06079_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7908" *) _06467_;
  assign _06080_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7918" *) _06468_;
  assign _06081_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7928" *) _06469_;
  assign _06082_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7938" *) _06470_;
  assign _06083_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7948" *) _06471_;
  assign _06084_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7958" *) _06472_;
  assign _06085_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7968" *) _06473_;
  assign _06086_ = wt_pre_sel[1] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7978" *) _06474_;
  assign _06087_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8014" *) cfg_is_fp16_d1[68];
  assign _06088_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8044" *) _06475_;
  assign _06089_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8054" *) _06476_;
  assign _06090_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8064" *) _06477_;
  assign _06091_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8074" *) _06478_;
  assign _06092_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8084" *) _06479_;
  assign _06093_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8094" *) _06480_;
  assign _06094_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8104" *) _06481_;
  assign _06095_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8114" *) _06482_;
  assign _06096_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8124" *) _06483_;
  assign _06097_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8134" *) _06484_;
  assign _06098_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8144" *) _06485_;
  assign _06099_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8154" *) _06486_;
  assign _06100_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8164" *) _06487_;
  assign _06101_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8174" *) _06488_;
  assign _06102_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8184" *) _06489_;
  assign _06103_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8194" *) _06490_;
  assign _06104_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8204" *) _06491_;
  assign _06105_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8214" *) _06492_;
  assign _06106_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8224" *) _06493_;
  assign _06107_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8234" *) _06494_;
  assign _06108_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8244" *) _06495_;
  assign _06109_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8254" *) _06496_;
  assign _06110_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8264" *) _06497_;
  assign _06111_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8274" *) _06498_;
  assign _06112_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8284" *) _06499_;
  assign _06113_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8294" *) _06500_;
  assign _06114_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8304" *) _06501_;
  assign _06115_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8314" *) _06502_;
  assign _06116_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8324" *) _06503_;
  assign _06117_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8334" *) _06504_;
  assign _06118_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8344" *) _06505_;
  assign _06119_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8354" *) _06506_;
  assign _06120_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8364" *) _06507_;
  assign _06121_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8374" *) _06508_;
  assign _06122_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8384" *) _06509_;
  assign _06123_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8394" *) _06510_;
  assign _06124_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8404" *) _06511_;
  assign _06125_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8414" *) _06512_;
  assign _06126_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8424" *) _06513_;
  assign _06127_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8434" *) _06514_;
  assign _06128_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8444" *) _06515_;
  assign _06129_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8454" *) _06516_;
  assign _06130_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8464" *) _06517_;
  assign _06131_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8474" *) _06518_;
  assign _06132_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8484" *) _06519_;
  assign _06133_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8494" *) _06520_;
  assign _06134_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8504" *) _06521_;
  assign _06135_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8514" *) _06522_;
  assign _06136_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8524" *) _06523_;
  assign _06137_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8534" *) _06524_;
  assign _06138_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8544" *) _06525_;
  assign _06139_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8554" *) _06526_;
  assign _06140_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8564" *) _06527_;
  assign _06141_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8574" *) _06528_;
  assign _06142_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8584" *) _06529_;
  assign _06143_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8594" *) _06530_;
  assign _06144_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8604" *) _06531_;
  assign _06145_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8614" *) _06532_;
  assign _06146_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8624" *) _06533_;
  assign _06147_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8634" *) _06534_;
  assign _06148_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8644" *) _06535_;
  assign _06149_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8654" *) _06536_;
  assign _06150_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8664" *) _06409_;
  assign _06151_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8674" *) _06410_;
  assign _06152_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8684" *) _06411_;
  assign _06153_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8694" *) _06412_;
  assign _06154_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8704" *) _06413_;
  assign _06155_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8714" *) _06414_;
  assign _06156_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8724" *) _06415_;
  assign _06157_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8734" *) _06416_;
  assign _06158_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8744" *) _06417_;
  assign _06159_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8754" *) _06418_;
  assign _06160_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8764" *) _06419_;
  assign _06161_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8774" *) _06420_;
  assign _06162_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8784" *) _06421_;
  assign _06163_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8794" *) _06422_;
  assign _06164_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8804" *) _06423_;
  assign _06165_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8814" *) _06424_;
  assign _06166_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8824" *) _06425_;
  assign _06167_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8834" *) _06426_;
  assign _06168_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8844" *) _06427_;
  assign _06169_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8854" *) _06428_;
  assign _06170_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8864" *) _06429_;
  assign _06171_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8874" *) _06430_;
  assign _06172_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8884" *) _06431_;
  assign _06173_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8894" *) _06432_;
  assign _06174_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8904" *) _06433_;
  assign _06175_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8914" *) _06434_;
  assign _06176_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8924" *) _06435_;
  assign _06177_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8934" *) _06436_;
  assign _06178_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8944" *) _06437_;
  assign _06179_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8954" *) _06438_;
  assign _06180_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8964" *) _06439_;
  assign _06181_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8974" *) _06440_;
  assign _06182_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8984" *) _06441_;
  assign _06183_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8994" *) _06442_;
  assign _06184_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9004" *) _06443_;
  assign _06185_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9014" *) _06444_;
  assign _06186_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9024" *) _06445_;
  assign _06187_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9034" *) _06446_;
  assign _06188_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9044" *) _06447_;
  assign _06189_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9054" *) _06448_;
  assign _06190_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9064" *) _06449_;
  assign _06191_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9074" *) _06450_;
  assign _06192_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9084" *) _06451_;
  assign _06193_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9094" *) _06452_;
  assign _06194_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9104" *) _06453_;
  assign _06195_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9114" *) _06454_;
  assign _06196_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9124" *) _06455_;
  assign _06197_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9134" *) _06456_;
  assign _06198_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9144" *) _06457_;
  assign _06199_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9154" *) _06458_;
  assign _06200_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9164" *) _06459_;
  assign _06201_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9174" *) _06460_;
  assign _06202_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9184" *) _06461_;
  assign _06203_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9194" *) _06462_;
  assign _06204_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9204" *) _06463_;
  assign _06205_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9214" *) _06464_;
  assign _06206_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9224" *) _06465_;
  assign _06207_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9234" *) _06466_;
  assign _06208_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9244" *) _06467_;
  assign _06209_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9254" *) _06468_;
  assign _06210_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9264" *) _06469_;
  assign _06211_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9274" *) _06470_;
  assign _06212_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9284" *) _06471_;
  assign _06213_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9294" *) _06472_;
  assign _06214_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9304" *) _06473_;
  assign _06215_ = wt_pre_sel[2] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9314" *) _06474_;
  assign _06216_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9350" *) cfg_is_fp16_d1[69];
  assign _06217_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9380" *) _06475_;
  assign _06218_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9390" *) _06476_;
  assign _06219_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9400" *) _06477_;
  assign _06220_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9410" *) _06478_;
  assign _06221_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9420" *) _06479_;
  assign _06222_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9430" *) _06480_;
  assign _06223_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9440" *) _06481_;
  assign _06224_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9450" *) _06482_;
  assign _06225_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9460" *) _06483_;
  assign _06226_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9470" *) _06484_;
  assign _06227_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9480" *) _06485_;
  assign _06228_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9490" *) _06486_;
  assign _06229_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9500" *) _06487_;
  assign _06230_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9510" *) _06488_;
  assign _06231_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9520" *) _06489_;
  assign _06232_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9530" *) _06490_;
  assign _06233_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9540" *) _06491_;
  assign _06234_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9550" *) _06492_;
  assign _06235_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9560" *) _06493_;
  assign _06236_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9570" *) _06494_;
  assign _06237_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9580" *) _06495_;
  assign _06238_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9590" *) _06496_;
  assign _06239_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9600" *) _06497_;
  assign _06240_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9610" *) _06498_;
  assign _06241_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9620" *) _06499_;
  assign _06242_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9630" *) _06500_;
  assign _06243_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9640" *) _06501_;
  assign _06244_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9650" *) _06502_;
  assign _06245_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9660" *) _06503_;
  assign _06246_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9670" *) _06504_;
  assign _06247_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9680" *) _06505_;
  assign _06248_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9690" *) _06506_;
  assign _06249_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9700" *) _06507_;
  assign _06250_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9710" *) _06508_;
  assign _06251_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9720" *) _06509_;
  assign _06252_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9730" *) _06510_;
  assign _06253_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9740" *) _06511_;
  assign _06254_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9750" *) _06512_;
  assign _06255_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9760" *) _06513_;
  assign _06256_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9770" *) _06514_;
  assign _06257_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9780" *) _06515_;
  assign _06258_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9790" *) _06516_;
  assign _06259_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9800" *) _06517_;
  assign _06260_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9810" *) _06518_;
  assign _06261_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9820" *) _06519_;
  assign _06262_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9830" *) _06520_;
  assign _06263_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9840" *) _06521_;
  assign _06264_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9850" *) _06522_;
  assign _06265_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9860" *) _06523_;
  assign _06266_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9870" *) _06524_;
  assign _06267_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9880" *) _06525_;
  assign _06268_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9890" *) _06526_;
  assign _06269_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9900" *) _06527_;
  assign _06270_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9910" *) _06528_;
  assign _06271_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9920" *) _06529_;
  assign _06272_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9930" *) _06530_;
  assign _06273_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9940" *) _06531_;
  assign _06274_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9950" *) _06532_;
  assign _06275_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9960" *) _06533_;
  assign _06276_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9970" *) _06534_;
  assign _06277_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9980" *) _06535_;
  assign _06278_ = wt_pre_sel[3] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9990" *) _06536_;
  assign _06407_ = ~ (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29041" *) dat_has_nan;
  assign _06408_ = ~ (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3968" *) wt_has_nan;
  assign _06409_ = wt_pre_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10000" *) wt_pre_nan[31];
  assign _06410_ = wt_pre_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10010" *) wt_pre_nan[31];
  assign _06411_ = wt_pre_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10020" *) wt_pre_nan[32];
  assign _06412_ = wt_pre_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10030" *) wt_pre_nan[32];
  assign _06413_ = wt_pre_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10040" *) wt_pre_nan[33];
  assign _06414_ = wt_pre_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10050" *) wt_pre_nan[33];
  assign _06415_ = wt_pre_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10060" *) wt_pre_nan[34];
  assign _06416_ = wt_pre_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10070" *) wt_pre_nan[34];
  assign _06417_ = wt_pre_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10080" *) wt_pre_nan[35];
  assign _06418_ = wt_pre_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10090" *) wt_pre_nan[35];
  assign _06419_ = wt_pre_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10100" *) wt_pre_nan[36];
  assign _06420_ = wt_pre_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10110" *) wt_pre_nan[36];
  assign _06421_ = wt_pre_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10120" *) wt_pre_nan[37];
  assign _06422_ = wt_pre_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10130" *) wt_pre_nan[37];
  assign _06423_ = wt_pre_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10140" *) wt_pre_nan[38];
  assign _06424_ = wt_pre_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10150" *) wt_pre_nan[38];
  assign _06425_ = wt_pre_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10160" *) wt_pre_nan[39];
  assign _06426_ = wt_pre_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10170" *) wt_pre_nan[39];
  assign _06427_ = wt_pre_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10180" *) wt_pre_nan[40];
  assign _06428_ = wt_pre_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10190" *) wt_pre_nan[40];
  assign _06429_ = wt_pre_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10200" *) wt_pre_nan[41];
  assign _06430_ = wt_pre_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10210" *) wt_pre_nan[41];
  assign _06431_ = wt_pre_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10220" *) wt_pre_nan[42];
  assign _06432_ = wt_pre_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10230" *) wt_pre_nan[42];
  assign _06433_ = wt_pre_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10240" *) wt_pre_nan[43];
  assign _06434_ = wt_pre_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10250" *) wt_pre_nan[43];
  assign _06435_ = wt_pre_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10260" *) wt_pre_nan[44];
  assign _06436_ = wt_pre_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10270" *) wt_pre_nan[44];
  assign _06437_ = wt_pre_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10280" *) wt_pre_nan[45];
  assign _06438_ = wt_pre_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10290" *) wt_pre_nan[45];
  assign _06439_ = wt_pre_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10300" *) wt_pre_nan[46];
  assign _06440_ = wt_pre_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10310" *) wt_pre_nan[46];
  assign _06441_ = wt_pre_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10320" *) wt_pre_nan[47];
  assign _06442_ = wt_pre_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10330" *) wt_pre_nan[47];
  assign _06443_ = wt_pre_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10340" *) wt_pre_nan[48];
  assign _06444_ = wt_pre_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10350" *) wt_pre_nan[48];
  assign _06445_ = wt_pre_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10360" *) wt_pre_nan[49];
  assign _06446_ = wt_pre_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10370" *) wt_pre_nan[49];
  assign _06447_ = wt_pre_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10380" *) wt_pre_nan[50];
  assign _06448_ = wt_pre_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10390" *) wt_pre_nan[50];
  assign _06449_ = wt_pre_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10400" *) wt_pre_nan[51];
  assign _06450_ = wt_pre_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10410" *) wt_pre_nan[51];
  assign _06451_ = wt_pre_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10420" *) wt_pre_nan[52];
  assign _06452_ = wt_pre_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10430" *) wt_pre_nan[52];
  assign _06453_ = wt_pre_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10440" *) wt_pre_nan[53];
  assign _06454_ = wt_pre_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10450" *) wt_pre_nan[53];
  assign _06455_ = wt_pre_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10460" *) wt_pre_nan[54];
  assign _06456_ = wt_pre_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10470" *) wt_pre_nan[54];
  assign _06457_ = wt_pre_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10480" *) wt_pre_nan[55];
  assign _06458_ = wt_pre_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10490" *) wt_pre_nan[55];
  assign _06459_ = wt_pre_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10500" *) wt_pre_nan[56];
  assign _06460_ = wt_pre_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10510" *) wt_pre_nan[56];
  assign _06461_ = wt_pre_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10520" *) wt_pre_nan[57];
  assign _06462_ = wt_pre_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10530" *) wt_pre_nan[57];
  assign _06463_ = wt_pre_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10540" *) wt_pre_nan[58];
  assign _06464_ = wt_pre_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10550" *) wt_pre_nan[58];
  assign _06465_ = wt_pre_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10560" *) wt_pre_nan[59];
  assign _06466_ = wt_pre_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10570" *) wt_pre_nan[59];
  assign _06467_ = wt_pre_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10580" *) wt_pre_nan[60];
  assign _06468_ = wt_pre_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10590" *) wt_pre_nan[60];
  assign _06469_ = wt_pre_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10600" *) wt_pre_nan[61];
  assign _06470_ = wt_pre_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10610" *) wt_pre_nan[61];
  assign _06471_ = wt_pre_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10620" *) wt_pre_nan[62];
  assign _06472_ = wt_pre_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10630" *) wt_pre_nan[62];
  assign _06473_ = wt_pre_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10640" *) wt_pre_nan[63];
  assign _06474_ = wt_pre_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10650" *) wt_pre_nan[63];
  assign _06475_ = wt_pre_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10716" *) wt_pre_nan[0];
  assign _06476_ = wt_pre_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10726" *) wt_pre_nan[0];
  assign _06477_ = wt_pre_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10736" *) wt_pre_nan[1];
  assign _06478_ = wt_pre_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10746" *) wt_pre_nan[1];
  assign _06479_ = wt_pre_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10756" *) wt_pre_nan[2];
  assign _06480_ = wt_pre_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10766" *) wt_pre_nan[2];
  assign _06481_ = wt_pre_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10776" *) wt_pre_nan[3];
  assign _06482_ = wt_pre_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10786" *) wt_pre_nan[3];
  assign _06483_ = wt_pre_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10796" *) wt_pre_nan[4];
  assign _06484_ = wt_pre_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10806" *) wt_pre_nan[4];
  assign _06485_ = wt_pre_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10816" *) wt_pre_nan[5];
  assign _06486_ = wt_pre_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10826" *) wt_pre_nan[5];
  assign _06487_ = wt_pre_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10836" *) wt_pre_nan[6];
  assign _06488_ = wt_pre_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10846" *) wt_pre_nan[6];
  assign _06489_ = wt_pre_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10856" *) wt_pre_nan[7];
  assign _06490_ = wt_pre_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10866" *) wt_pre_nan[7];
  assign _06491_ = wt_pre_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10876" *) wt_pre_nan[8];
  assign _06492_ = wt_pre_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10886" *) wt_pre_nan[8];
  assign _06493_ = wt_pre_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10896" *) wt_pre_nan[9];
  assign _06494_ = wt_pre_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10906" *) wt_pre_nan[9];
  assign _06495_ = wt_pre_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10916" *) wt_pre_nan[10];
  assign _06496_ = wt_pre_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10926" *) wt_pre_nan[10];
  assign _06497_ = wt_pre_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10936" *) wt_pre_nan[11];
  assign _06498_ = wt_pre_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10946" *) wt_pre_nan[11];
  assign _06499_ = wt_pre_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10956" *) wt_pre_nan[12];
  assign _06500_ = wt_pre_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10966" *) wt_pre_nan[12];
  assign _06501_ = wt_pre_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10976" *) wt_pre_nan[13];
  assign _06502_ = wt_pre_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10986" *) wt_pre_nan[13];
  assign _06503_ = wt_pre_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10996" *) wt_pre_nan[14];
  assign _06504_ = wt_pre_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11006" *) wt_pre_nan[14];
  assign _06505_ = wt_pre_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11016" *) wt_pre_nan[15];
  assign _06506_ = wt_pre_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11026" *) wt_pre_nan[15];
  assign _06507_ = wt_pre_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11036" *) wt_pre_nan[16];
  assign _06508_ = wt_pre_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11046" *) wt_pre_nan[16];
  assign _06509_ = wt_pre_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11056" *) wt_pre_nan[17];
  assign _06510_ = wt_pre_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11066" *) wt_pre_nan[17];
  assign _06511_ = wt_pre_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11076" *) wt_pre_nan[18];
  assign _06512_ = wt_pre_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11086" *) wt_pre_nan[18];
  assign _06513_ = wt_pre_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11096" *) wt_pre_nan[19];
  assign _06514_ = wt_pre_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11106" *) wt_pre_nan[19];
  assign _06515_ = wt_pre_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11116" *) wt_pre_nan[20];
  assign _06516_ = wt_pre_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11126" *) wt_pre_nan[20];
  assign _06517_ = wt_pre_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11136" *) wt_pre_nan[21];
  assign _06518_ = wt_pre_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11146" *) wt_pre_nan[21];
  assign _06519_ = wt_pre_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11156" *) wt_pre_nan[22];
  assign _06520_ = wt_pre_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11166" *) wt_pre_nan[22];
  assign _06521_ = wt_pre_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11176" *) wt_pre_nan[23];
  assign _06522_ = wt_pre_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11186" *) wt_pre_nan[23];
  assign _06523_ = wt_pre_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11196" *) wt_pre_nan[24];
  assign _06524_ = wt_pre_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11206" *) wt_pre_nan[24];
  assign _06525_ = wt_pre_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11216" *) wt_pre_nan[25];
  assign _06526_ = wt_pre_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11226" *) wt_pre_nan[25];
  assign _06527_ = wt_pre_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11236" *) wt_pre_nan[26];
  assign _06528_ = wt_pre_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11246" *) wt_pre_nan[26];
  assign _06529_ = wt_pre_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11256" *) wt_pre_nan[27];
  assign _06530_ = wt_pre_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11266" *) wt_pre_nan[27];
  assign _06531_ = wt_pre_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11276" *) wt_pre_nan[28];
  assign _06532_ = wt_pre_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11286" *) wt_pre_nan[28];
  assign _06533_ = wt_pre_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11296" *) wt_pre_nan[29];
  assign _06534_ = wt_pre_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11306" *) wt_pre_nan[29];
  assign _06535_ = wt_pre_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11316" *) wt_pre_nan[30];
  assign _06536_ = wt_pre_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11326" *) wt_pre_nan[30];
  assign _06537_ = wt0_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16049" *) wt0_sd_nan[0];
  assign _06538_ = wt0_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16059" *) wt0_sd_nan[0];
  assign _06539_ = wt0_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16069" *) wt0_sd_nan[1];
  assign _06540_ = wt0_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16079" *) wt0_sd_nan[1];
  assign _06541_ = wt0_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16089" *) wt0_sd_nan[2];
  assign _06542_ = wt0_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16099" *) wt0_sd_nan[2];
  assign _06543_ = wt0_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16109" *) wt0_sd_nan[3];
  assign _06544_ = wt0_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16119" *) wt0_sd_nan[3];
  assign _06545_ = wt0_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16129" *) wt0_sd_nan[4];
  assign _06546_ = wt0_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16139" *) wt0_sd_nan[4];
  assign _06547_ = wt0_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16149" *) wt0_sd_nan[5];
  assign _06548_ = wt0_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16159" *) wt0_sd_nan[5];
  assign _06549_ = wt0_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16169" *) wt0_sd_nan[6];
  assign _06550_ = wt0_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16179" *) wt0_sd_nan[6];
  assign _06551_ = wt0_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16189" *) wt0_sd_nan[7];
  assign _06552_ = wt0_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16199" *) wt0_sd_nan[7];
  assign _06553_ = wt0_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16209" *) wt0_sd_nan[8];
  assign _06554_ = wt0_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16219" *) wt0_sd_nan[8];
  assign _06555_ = wt0_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16229" *) wt0_sd_nan[9];
  assign _06556_ = wt0_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16239" *) wt0_sd_nan[9];
  assign _06557_ = wt0_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16249" *) wt0_sd_nan[10];
  assign _06558_ = wt0_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16259" *) wt0_sd_nan[10];
  assign _06559_ = wt0_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16269" *) wt0_sd_nan[11];
  assign _06560_ = wt0_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16279" *) wt0_sd_nan[11];
  assign _06561_ = wt0_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16289" *) wt0_sd_nan[12];
  assign _06562_ = wt0_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16299" *) wt0_sd_nan[12];
  assign _06563_ = wt0_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16309" *) wt0_sd_nan[13];
  assign _06564_ = wt0_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16319" *) wt0_sd_nan[13];
  assign _06565_ = wt0_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16329" *) wt0_sd_nan[14];
  assign _06566_ = wt0_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16339" *) wt0_sd_nan[14];
  assign _06567_ = wt0_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16349" *) wt0_sd_nan[15];
  assign _06568_ = wt0_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16359" *) wt0_sd_nan[15];
  assign _06569_ = wt0_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16369" *) wt0_sd_nan[16];
  assign _06570_ = wt0_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16379" *) wt0_sd_nan[16];
  assign _06571_ = wt0_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16389" *) wt0_sd_nan[17];
  assign _06572_ = wt0_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16399" *) wt0_sd_nan[17];
  assign _06573_ = wt0_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16409" *) wt0_sd_nan[18];
  assign _06574_ = wt0_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16419" *) wt0_sd_nan[18];
  assign _06575_ = wt0_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16429" *) wt0_sd_nan[19];
  assign _06576_ = wt0_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16439" *) wt0_sd_nan[19];
  assign _06577_ = wt0_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16449" *) wt0_sd_nan[20];
  assign _06578_ = wt0_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16459" *) wt0_sd_nan[20];
  assign _06579_ = wt0_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16469" *) wt0_sd_nan[21];
  assign _06580_ = wt0_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16479" *) wt0_sd_nan[21];
  assign _06581_ = wt0_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16489" *) wt0_sd_nan[22];
  assign _06582_ = wt0_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16499" *) wt0_sd_nan[22];
  assign _06583_ = wt0_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16509" *) wt0_sd_nan[23];
  assign _06584_ = wt0_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16519" *) wt0_sd_nan[23];
  assign _06585_ = wt0_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16529" *) wt0_sd_nan[24];
  assign _06586_ = wt0_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16539" *) wt0_sd_nan[24];
  assign _06587_ = wt0_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16549" *) wt0_sd_nan[25];
  assign _06588_ = wt0_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16559" *) wt0_sd_nan[25];
  assign _06589_ = wt0_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16569" *) wt0_sd_nan[26];
  assign _06590_ = wt0_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16579" *) wt0_sd_nan[26];
  assign _06591_ = wt0_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16589" *) wt0_sd_nan[27];
  assign _06592_ = wt0_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16599" *) wt0_sd_nan[27];
  assign _06593_ = wt0_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16609" *) wt0_sd_nan[28];
  assign _06594_ = wt0_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16619" *) wt0_sd_nan[28];
  assign _06595_ = wt0_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16629" *) wt0_sd_nan[29];
  assign _06596_ = wt0_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16639" *) wt0_sd_nan[29];
  assign _06597_ = wt0_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16649" *) wt0_sd_nan[30];
  assign _06598_ = wt0_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16659" *) wt0_sd_nan[30];
  assign _06599_ = wt0_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16669" *) wt0_sd_nan[31];
  assign _06600_ = wt0_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16679" *) wt0_sd_nan[31];
  assign _06601_ = wt0_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16689" *) wt0_sd_nan[32];
  assign _06602_ = wt0_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16699" *) wt0_sd_nan[32];
  assign _06603_ = wt0_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16709" *) wt0_sd_nan[33];
  assign _06604_ = wt0_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16719" *) wt0_sd_nan[33];
  assign _06605_ = wt0_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16729" *) wt0_sd_nan[34];
  assign _06606_ = wt0_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16739" *) wt0_sd_nan[34];
  assign _06607_ = wt0_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16749" *) wt0_sd_nan[35];
  assign _06608_ = wt0_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16759" *) wt0_sd_nan[35];
  assign _06609_ = wt0_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16769" *) wt0_sd_nan[36];
  assign _06610_ = wt0_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16779" *) wt0_sd_nan[36];
  assign _06611_ = wt0_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16789" *) wt0_sd_nan[37];
  assign _06612_ = wt0_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16799" *) wt0_sd_nan[37];
  assign _06613_ = wt0_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16809" *) wt0_sd_nan[38];
  assign _06614_ = wt0_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16819" *) wt0_sd_nan[38];
  assign _06615_ = wt0_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16829" *) wt0_sd_nan[39];
  assign _06616_ = wt0_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16839" *) wt0_sd_nan[39];
  assign _06617_ = wt0_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16849" *) wt0_sd_nan[40];
  assign _06618_ = wt0_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16859" *) wt0_sd_nan[40];
  assign _06619_ = wt0_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16869" *) wt0_sd_nan[41];
  assign _06620_ = wt0_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16879" *) wt0_sd_nan[41];
  assign _06621_ = wt0_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16889" *) wt0_sd_nan[42];
  assign _06622_ = wt0_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16899" *) wt0_sd_nan[42];
  assign _06623_ = wt0_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16909" *) wt0_sd_nan[43];
  assign _06624_ = wt0_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16919" *) wt0_sd_nan[43];
  assign _06625_ = wt0_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16929" *) wt0_sd_nan[44];
  assign _06626_ = wt0_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16939" *) wt0_sd_nan[44];
  assign _06627_ = wt0_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16949" *) wt0_sd_nan[45];
  assign _06628_ = wt0_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16959" *) wt0_sd_nan[45];
  assign _06629_ = wt0_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16969" *) wt0_sd_nan[46];
  assign _06630_ = wt0_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16979" *) wt0_sd_nan[46];
  assign _06631_ = wt0_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16989" *) wt0_sd_nan[47];
  assign _06632_ = wt0_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16999" *) wt0_sd_nan[47];
  assign _06633_ = wt0_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17009" *) wt0_sd_nan[48];
  assign _06634_ = wt0_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17019" *) wt0_sd_nan[48];
  assign _06635_ = wt0_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17029" *) wt0_sd_nan[49];
  assign _06636_ = wt0_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17039" *) wt0_sd_nan[49];
  assign _06637_ = wt0_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17049" *) wt0_sd_nan[50];
  assign _06638_ = wt0_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17059" *) wt0_sd_nan[50];
  assign _06639_ = wt0_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17069" *) wt0_sd_nan[51];
  assign _06640_ = wt0_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17079" *) wt0_sd_nan[51];
  assign _06641_ = wt0_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17089" *) wt0_sd_nan[52];
  assign _06642_ = wt0_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17099" *) wt0_sd_nan[52];
  assign _06643_ = wt0_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17109" *) wt0_sd_nan[53];
  assign _06644_ = wt0_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17119" *) wt0_sd_nan[53];
  assign _06645_ = wt0_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17129" *) wt0_sd_nan[54];
  assign _06646_ = wt0_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17139" *) wt0_sd_nan[54];
  assign _06647_ = wt0_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17149" *) wt0_sd_nan[55];
  assign _06648_ = wt0_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17159" *) wt0_sd_nan[55];
  assign _06649_ = wt0_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17169" *) wt0_sd_nan[56];
  assign _06650_ = wt0_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17179" *) wt0_sd_nan[56];
  assign _06651_ = wt0_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17189" *) wt0_sd_nan[57];
  assign _06652_ = wt0_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17199" *) wt0_sd_nan[57];
  assign _06653_ = wt0_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17209" *) wt0_sd_nan[58];
  assign _06654_ = wt0_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17219" *) wt0_sd_nan[58];
  assign _06655_ = wt0_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17229" *) wt0_sd_nan[59];
  assign _06656_ = wt0_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17239" *) wt0_sd_nan[59];
  assign _06657_ = wt0_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17249" *) wt0_sd_nan[60];
  assign _06658_ = wt0_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17259" *) wt0_sd_nan[60];
  assign _06659_ = wt0_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17269" *) wt0_sd_nan[61];
  assign _06660_ = wt0_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17279" *) wt0_sd_nan[61];
  assign _06661_ = wt0_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17289" *) wt0_sd_nan[62];
  assign _06662_ = wt0_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17299" *) wt0_sd_nan[62];
  assign _06663_ = wt0_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17309" *) wt0_sd_nan[63];
  assign _06664_ = wt0_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17319" *) wt0_sd_nan[63];
  assign _06665_ = wt1_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17373" *) wt1_sd_nan[0];
  assign _06666_ = wt1_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17383" *) wt1_sd_nan[0];
  assign _06667_ = wt1_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17393" *) wt1_sd_nan[1];
  assign _06668_ = wt1_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17403" *) wt1_sd_nan[1];
  assign _06669_ = wt1_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17413" *) wt1_sd_nan[2];
  assign _06670_ = wt1_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17423" *) wt1_sd_nan[2];
  assign _06671_ = wt1_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17433" *) wt1_sd_nan[3];
  assign _06672_ = wt1_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17443" *) wt1_sd_nan[3];
  assign _06673_ = wt1_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17453" *) wt1_sd_nan[4];
  assign _06674_ = wt1_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17463" *) wt1_sd_nan[4];
  assign _06675_ = wt1_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17473" *) wt1_sd_nan[5];
  assign _06676_ = wt1_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17483" *) wt1_sd_nan[5];
  assign _06677_ = wt1_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17493" *) wt1_sd_nan[6];
  assign _06678_ = wt1_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17503" *) wt1_sd_nan[6];
  assign _06679_ = wt1_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17513" *) wt1_sd_nan[7];
  assign _06680_ = wt1_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17523" *) wt1_sd_nan[7];
  assign _06681_ = wt1_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17533" *) wt1_sd_nan[8];
  assign _06682_ = wt1_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17543" *) wt1_sd_nan[8];
  assign _06683_ = wt1_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17553" *) wt1_sd_nan[9];
  assign _06684_ = wt1_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17563" *) wt1_sd_nan[9];
  assign _06685_ = wt1_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17573" *) wt1_sd_nan[10];
  assign _06686_ = wt1_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17583" *) wt1_sd_nan[10];
  assign _06687_ = wt1_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17593" *) wt1_sd_nan[11];
  assign _06688_ = wt1_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17603" *) wt1_sd_nan[11];
  assign _06689_ = wt1_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17613" *) wt1_sd_nan[12];
  assign _06690_ = wt1_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17623" *) wt1_sd_nan[12];
  assign _06691_ = wt1_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17633" *) wt1_sd_nan[13];
  assign _06692_ = wt1_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17643" *) wt1_sd_nan[13];
  assign _06693_ = wt1_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17653" *) wt1_sd_nan[14];
  assign _06694_ = wt1_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17663" *) wt1_sd_nan[14];
  assign _06695_ = wt1_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17673" *) wt1_sd_nan[15];
  assign _06696_ = wt1_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17683" *) wt1_sd_nan[15];
  assign _06697_ = wt1_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17693" *) wt1_sd_nan[16];
  assign _06698_ = wt1_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17703" *) wt1_sd_nan[16];
  assign _06699_ = wt1_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17713" *) wt1_sd_nan[17];
  assign _06700_ = wt1_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17723" *) wt1_sd_nan[17];
  assign _06701_ = wt1_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17733" *) wt1_sd_nan[18];
  assign _06702_ = wt1_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17743" *) wt1_sd_nan[18];
  assign _06703_ = wt1_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17753" *) wt1_sd_nan[19];
  assign _06704_ = wt1_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17763" *) wt1_sd_nan[19];
  assign _06705_ = wt1_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17773" *) wt1_sd_nan[20];
  assign _06706_ = wt1_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17783" *) wt1_sd_nan[20];
  assign _06707_ = wt1_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17793" *) wt1_sd_nan[21];
  assign _06708_ = wt1_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17803" *) wt1_sd_nan[21];
  assign _06709_ = wt1_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17813" *) wt1_sd_nan[22];
  assign _06710_ = wt1_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17823" *) wt1_sd_nan[22];
  assign _06711_ = wt1_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17833" *) wt1_sd_nan[23];
  assign _06712_ = wt1_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17843" *) wt1_sd_nan[23];
  assign _06713_ = wt1_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17853" *) wt1_sd_nan[24];
  assign _06714_ = wt1_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17863" *) wt1_sd_nan[24];
  assign _06715_ = wt1_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17873" *) wt1_sd_nan[25];
  assign _06716_ = wt1_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17883" *) wt1_sd_nan[25];
  assign _06717_ = wt1_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17893" *) wt1_sd_nan[26];
  assign _06718_ = wt1_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17903" *) wt1_sd_nan[26];
  assign _06719_ = wt1_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17913" *) wt1_sd_nan[27];
  assign _06720_ = wt1_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17923" *) wt1_sd_nan[27];
  assign _06721_ = wt1_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17933" *) wt1_sd_nan[28];
  assign _06722_ = wt1_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17943" *) wt1_sd_nan[28];
  assign _06723_ = wt1_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17953" *) wt1_sd_nan[29];
  assign _06724_ = wt1_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17963" *) wt1_sd_nan[29];
  assign _06725_ = wt1_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17973" *) wt1_sd_nan[30];
  assign _06726_ = wt1_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17983" *) wt1_sd_nan[30];
  assign _06727_ = wt1_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17993" *) wt1_sd_nan[31];
  assign _06728_ = wt1_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18003" *) wt1_sd_nan[31];
  assign _06729_ = wt1_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18013" *) wt1_sd_nan[32];
  assign _06730_ = wt1_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18023" *) wt1_sd_nan[32];
  assign _06731_ = wt1_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18033" *) wt1_sd_nan[33];
  assign _06732_ = wt1_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18043" *) wt1_sd_nan[33];
  assign _06733_ = wt1_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18053" *) wt1_sd_nan[34];
  assign _06734_ = wt1_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18063" *) wt1_sd_nan[34];
  assign _06735_ = wt1_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18073" *) wt1_sd_nan[35];
  assign _06736_ = wt1_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18083" *) wt1_sd_nan[35];
  assign _06737_ = wt1_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18093" *) wt1_sd_nan[36];
  assign _06738_ = wt1_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18103" *) wt1_sd_nan[36];
  assign _06739_ = wt1_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18113" *) wt1_sd_nan[37];
  assign _06740_ = wt1_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18123" *) wt1_sd_nan[37];
  assign _06741_ = wt1_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18133" *) wt1_sd_nan[38];
  assign _06742_ = wt1_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18143" *) wt1_sd_nan[38];
  assign _06743_ = wt1_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18153" *) wt1_sd_nan[39];
  assign _06744_ = wt1_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18163" *) wt1_sd_nan[39];
  assign _06745_ = wt1_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18173" *) wt1_sd_nan[40];
  assign _06746_ = wt1_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18183" *) wt1_sd_nan[40];
  assign _06747_ = wt1_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18193" *) wt1_sd_nan[41];
  assign _06748_ = wt1_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18203" *) wt1_sd_nan[41];
  assign _06749_ = wt1_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18213" *) wt1_sd_nan[42];
  assign _06750_ = wt1_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18223" *) wt1_sd_nan[42];
  assign _06751_ = wt1_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18233" *) wt1_sd_nan[43];
  assign _06752_ = wt1_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18243" *) wt1_sd_nan[43];
  assign _06753_ = wt1_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18253" *) wt1_sd_nan[44];
  assign _06754_ = wt1_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18263" *) wt1_sd_nan[44];
  assign _06755_ = wt1_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18273" *) wt1_sd_nan[45];
  assign _06756_ = wt1_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18283" *) wt1_sd_nan[45];
  assign _06757_ = wt1_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18293" *) wt1_sd_nan[46];
  assign _06758_ = wt1_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18303" *) wt1_sd_nan[46];
  assign _06759_ = wt1_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18313" *) wt1_sd_nan[47];
  assign _06760_ = wt1_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18323" *) wt1_sd_nan[47];
  assign _06761_ = wt1_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18333" *) wt1_sd_nan[48];
  assign _06762_ = wt1_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18343" *) wt1_sd_nan[48];
  assign _06763_ = wt1_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18353" *) wt1_sd_nan[49];
  assign _06764_ = wt1_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18363" *) wt1_sd_nan[49];
  assign _06765_ = wt1_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18373" *) wt1_sd_nan[50];
  assign _06766_ = wt1_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18383" *) wt1_sd_nan[50];
  assign _06767_ = wt1_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18393" *) wt1_sd_nan[51];
  assign _06768_ = wt1_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18403" *) wt1_sd_nan[51];
  assign _06769_ = wt1_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18413" *) wt1_sd_nan[52];
  assign _06770_ = wt1_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18423" *) wt1_sd_nan[52];
  assign _06771_ = wt1_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18433" *) wt1_sd_nan[53];
  assign _06772_ = wt1_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18443" *) wt1_sd_nan[53];
  assign _06773_ = wt1_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18453" *) wt1_sd_nan[54];
  assign _06774_ = wt1_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18463" *) wt1_sd_nan[54];
  assign _06775_ = wt1_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18473" *) wt1_sd_nan[55];
  assign _06776_ = wt1_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18483" *) wt1_sd_nan[55];
  assign _06777_ = wt1_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18493" *) wt1_sd_nan[56];
  assign _06778_ = wt1_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18503" *) wt1_sd_nan[56];
  assign _06779_ = wt1_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18513" *) wt1_sd_nan[57];
  assign _06780_ = wt1_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18523" *) wt1_sd_nan[57];
  assign _06781_ = wt1_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18533" *) wt1_sd_nan[58];
  assign _06782_ = wt1_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18543" *) wt1_sd_nan[58];
  assign _06783_ = wt1_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18553" *) wt1_sd_nan[59];
  assign _06784_ = wt1_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18563" *) wt1_sd_nan[59];
  assign _06785_ = wt1_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18573" *) wt1_sd_nan[60];
  assign _06786_ = wt1_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18583" *) wt1_sd_nan[60];
  assign _06787_ = wt1_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18593" *) wt1_sd_nan[61];
  assign _06788_ = wt1_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18603" *) wt1_sd_nan[61];
  assign _06789_ = wt1_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18613" *) wt1_sd_nan[62];
  assign _06790_ = wt1_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18623" *) wt1_sd_nan[62];
  assign _06791_ = wt1_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18633" *) wt1_sd_nan[63];
  assign _06792_ = wt1_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18643" *) wt1_sd_nan[63];
  assign _06793_ = wt2_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18697" *) wt2_sd_nan[0];
  assign _06794_ = wt2_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18707" *) wt2_sd_nan[0];
  assign _06795_ = wt2_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18717" *) wt2_sd_nan[1];
  assign _06796_ = wt2_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18727" *) wt2_sd_nan[1];
  assign _06797_ = wt2_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18737" *) wt2_sd_nan[2];
  assign _06798_ = wt2_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18747" *) wt2_sd_nan[2];
  assign _06799_ = wt2_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18757" *) wt2_sd_nan[3];
  assign _06800_ = wt2_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18767" *) wt2_sd_nan[3];
  assign _06801_ = wt2_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18777" *) wt2_sd_nan[4];
  assign _06802_ = wt2_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18787" *) wt2_sd_nan[4];
  assign _06803_ = wt2_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18797" *) wt2_sd_nan[5];
  assign _06804_ = wt2_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18807" *) wt2_sd_nan[5];
  assign _06805_ = wt2_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18817" *) wt2_sd_nan[6];
  assign _06806_ = wt2_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18827" *) wt2_sd_nan[6];
  assign _06807_ = wt2_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18837" *) wt2_sd_nan[7];
  assign _06808_ = wt2_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18847" *) wt2_sd_nan[7];
  assign _06809_ = wt2_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18857" *) wt2_sd_nan[8];
  assign _06810_ = wt2_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18867" *) wt2_sd_nan[8];
  assign _06811_ = wt2_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18877" *) wt2_sd_nan[9];
  assign _06812_ = wt2_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18887" *) wt2_sd_nan[9];
  assign _06813_ = wt2_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18897" *) wt2_sd_nan[10];
  assign _06814_ = wt2_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18907" *) wt2_sd_nan[10];
  assign _06815_ = wt2_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18917" *) wt2_sd_nan[11];
  assign _06816_ = wt2_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18927" *) wt2_sd_nan[11];
  assign _06817_ = wt2_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18937" *) wt2_sd_nan[12];
  assign _06818_ = wt2_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18947" *) wt2_sd_nan[12];
  assign _06819_ = wt2_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18957" *) wt2_sd_nan[13];
  assign _06820_ = wt2_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18967" *) wt2_sd_nan[13];
  assign _06821_ = wt2_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18977" *) wt2_sd_nan[14];
  assign _06822_ = wt2_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18987" *) wt2_sd_nan[14];
  assign _06823_ = wt2_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18997" *) wt2_sd_nan[15];
  assign _06824_ = wt2_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19007" *) wt2_sd_nan[15];
  assign _06825_ = wt2_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19017" *) wt2_sd_nan[16];
  assign _06826_ = wt2_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19027" *) wt2_sd_nan[16];
  assign _06827_ = wt2_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19037" *) wt2_sd_nan[17];
  assign _06828_ = wt2_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19047" *) wt2_sd_nan[17];
  assign _06829_ = wt2_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19057" *) wt2_sd_nan[18];
  assign _06830_ = wt2_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19067" *) wt2_sd_nan[18];
  assign _06831_ = wt2_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19077" *) wt2_sd_nan[19];
  assign _06832_ = wt2_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19087" *) wt2_sd_nan[19];
  assign _06833_ = wt2_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19097" *) wt2_sd_nan[20];
  assign _06834_ = wt2_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19107" *) wt2_sd_nan[20];
  assign _06835_ = wt2_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19117" *) wt2_sd_nan[21];
  assign _06836_ = wt2_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19127" *) wt2_sd_nan[21];
  assign _06837_ = wt2_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19137" *) wt2_sd_nan[22];
  assign _06838_ = wt2_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19147" *) wt2_sd_nan[22];
  assign _06839_ = wt2_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19157" *) wt2_sd_nan[23];
  assign _06840_ = wt2_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19167" *) wt2_sd_nan[23];
  assign _06841_ = wt2_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19177" *) wt2_sd_nan[24];
  assign _06842_ = wt2_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19187" *) wt2_sd_nan[24];
  assign _06843_ = wt2_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19197" *) wt2_sd_nan[25];
  assign _06844_ = wt2_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19207" *) wt2_sd_nan[25];
  assign _06845_ = wt2_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19217" *) wt2_sd_nan[26];
  assign _06846_ = wt2_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19227" *) wt2_sd_nan[26];
  assign _06847_ = wt2_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19237" *) wt2_sd_nan[27];
  assign _06848_ = wt2_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19247" *) wt2_sd_nan[27];
  assign _06849_ = wt2_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19257" *) wt2_sd_nan[28];
  assign _06850_ = wt2_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19267" *) wt2_sd_nan[28];
  assign _06851_ = wt2_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19277" *) wt2_sd_nan[29];
  assign _06852_ = wt2_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19287" *) wt2_sd_nan[29];
  assign _06853_ = wt2_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19297" *) wt2_sd_nan[30];
  assign _06854_ = wt2_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19307" *) wt2_sd_nan[30];
  assign _06855_ = wt2_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19317" *) wt2_sd_nan[31];
  assign _06856_ = wt2_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19327" *) wt2_sd_nan[31];
  assign _06857_ = wt2_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19337" *) wt2_sd_nan[32];
  assign _06858_ = wt2_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19347" *) wt2_sd_nan[32];
  assign _06859_ = wt2_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19357" *) wt2_sd_nan[33];
  assign _06860_ = wt2_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19367" *) wt2_sd_nan[33];
  assign _06861_ = wt2_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19377" *) wt2_sd_nan[34];
  assign _06862_ = wt2_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19387" *) wt2_sd_nan[34];
  assign _06863_ = wt2_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19397" *) wt2_sd_nan[35];
  assign _06864_ = wt2_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19407" *) wt2_sd_nan[35];
  assign _06865_ = wt2_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19417" *) wt2_sd_nan[36];
  assign _06866_ = wt2_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19427" *) wt2_sd_nan[36];
  assign _06867_ = wt2_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19437" *) wt2_sd_nan[37];
  assign _06868_ = wt2_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19447" *) wt2_sd_nan[37];
  assign _06869_ = wt2_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19457" *) wt2_sd_nan[38];
  assign _06870_ = wt2_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19467" *) wt2_sd_nan[38];
  assign _06871_ = wt2_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19477" *) wt2_sd_nan[39];
  assign _06872_ = wt2_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19487" *) wt2_sd_nan[39];
  assign _06873_ = wt2_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19497" *) wt2_sd_nan[40];
  assign _06874_ = wt2_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19507" *) wt2_sd_nan[40];
  assign _06875_ = wt2_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19517" *) wt2_sd_nan[41];
  assign _06876_ = wt2_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19527" *) wt2_sd_nan[41];
  assign _06877_ = wt2_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19537" *) wt2_sd_nan[42];
  assign _06878_ = wt2_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19547" *) wt2_sd_nan[42];
  assign _06879_ = wt2_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19557" *) wt2_sd_nan[43];
  assign _06880_ = wt2_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19567" *) wt2_sd_nan[43];
  assign _06881_ = wt2_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19577" *) wt2_sd_nan[44];
  assign _06882_ = wt2_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19587" *) wt2_sd_nan[44];
  assign _06883_ = wt2_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19597" *) wt2_sd_nan[45];
  assign _06884_ = wt2_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19607" *) wt2_sd_nan[45];
  assign _06885_ = wt2_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19617" *) wt2_sd_nan[46];
  assign _06886_ = wt2_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19627" *) wt2_sd_nan[46];
  assign _06887_ = wt2_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19637" *) wt2_sd_nan[47];
  assign _06888_ = wt2_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19647" *) wt2_sd_nan[47];
  assign _06889_ = wt2_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19657" *) wt2_sd_nan[48];
  assign _06890_ = wt2_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19667" *) wt2_sd_nan[48];
  assign _06891_ = wt2_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19677" *) wt2_sd_nan[49];
  assign _06892_ = wt2_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19687" *) wt2_sd_nan[49];
  assign _06893_ = wt2_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19697" *) wt2_sd_nan[50];
  assign _06894_ = wt2_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19707" *) wt2_sd_nan[50];
  assign _06895_ = wt2_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19717" *) wt2_sd_nan[51];
  assign _06896_ = wt2_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19727" *) wt2_sd_nan[51];
  assign _06897_ = wt2_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19737" *) wt2_sd_nan[52];
  assign _06898_ = wt2_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19747" *) wt2_sd_nan[52];
  assign _06899_ = wt2_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19757" *) wt2_sd_nan[53];
  assign _06900_ = wt2_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19767" *) wt2_sd_nan[53];
  assign _06901_ = wt2_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19777" *) wt2_sd_nan[54];
  assign _06902_ = wt2_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19787" *) wt2_sd_nan[54];
  assign _06903_ = wt2_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19797" *) wt2_sd_nan[55];
  assign _06904_ = wt2_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19807" *) wt2_sd_nan[55];
  assign _06905_ = wt2_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19817" *) wt2_sd_nan[56];
  assign _06906_ = wt2_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19827" *) wt2_sd_nan[56];
  assign _06907_ = wt2_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19837" *) wt2_sd_nan[57];
  assign _06908_ = wt2_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19847" *) wt2_sd_nan[57];
  assign _06909_ = wt2_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19857" *) wt2_sd_nan[58];
  assign _06910_ = wt2_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19867" *) wt2_sd_nan[58];
  assign _06911_ = wt2_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19877" *) wt2_sd_nan[59];
  assign _06912_ = wt2_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19887" *) wt2_sd_nan[59];
  assign _06913_ = wt2_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19897" *) wt2_sd_nan[60];
  assign _06914_ = wt2_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19907" *) wt2_sd_nan[60];
  assign _06915_ = wt2_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19917" *) wt2_sd_nan[61];
  assign _06916_ = wt2_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19927" *) wt2_sd_nan[61];
  assign _06917_ = wt2_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19937" *) wt2_sd_nan[62];
  assign _06918_ = wt2_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19947" *) wt2_sd_nan[62];
  assign _06919_ = wt2_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19957" *) wt2_sd_nan[63];
  assign _06920_ = wt2_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19967" *) wt2_sd_nan[63];
  assign _06921_ = wt3_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20021" *) wt3_sd_nan[0];
  assign _06922_ = wt3_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20031" *) wt3_sd_nan[0];
  assign _06923_ = wt3_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20041" *) wt3_sd_nan[1];
  assign _06924_ = wt3_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20051" *) wt3_sd_nan[1];
  assign _06925_ = wt3_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20061" *) wt3_sd_nan[2];
  assign _06926_ = wt3_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20071" *) wt3_sd_nan[2];
  assign _06927_ = wt3_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20081" *) wt3_sd_nan[3];
  assign _06928_ = wt3_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20091" *) wt3_sd_nan[3];
  assign _06929_ = wt3_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20101" *) wt3_sd_nan[4];
  assign _06930_ = wt3_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20111" *) wt3_sd_nan[4];
  assign _06931_ = wt3_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20121" *) wt3_sd_nan[5];
  assign _06932_ = wt3_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20131" *) wt3_sd_nan[5];
  assign _06933_ = wt3_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20141" *) wt3_sd_nan[6];
  assign _06934_ = wt3_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20151" *) wt3_sd_nan[6];
  assign _06935_ = wt3_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20161" *) wt3_sd_nan[7];
  assign _06936_ = wt3_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20171" *) wt3_sd_nan[7];
  assign _06937_ = wt3_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20181" *) wt3_sd_nan[8];
  assign _06938_ = wt3_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20191" *) wt3_sd_nan[8];
  assign _06939_ = wt3_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20201" *) wt3_sd_nan[9];
  assign _06940_ = wt3_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20211" *) wt3_sd_nan[9];
  assign _06941_ = wt3_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20221" *) wt3_sd_nan[10];
  assign _06942_ = wt3_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20231" *) wt3_sd_nan[10];
  assign _06943_ = wt3_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20241" *) wt3_sd_nan[11];
  assign _06944_ = wt3_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20251" *) wt3_sd_nan[11];
  assign _06945_ = wt3_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20261" *) wt3_sd_nan[12];
  assign _06946_ = wt3_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20271" *) wt3_sd_nan[12];
  assign _06947_ = wt3_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20281" *) wt3_sd_nan[13];
  assign _06948_ = wt3_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20291" *) wt3_sd_nan[13];
  assign _06949_ = wt3_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20301" *) wt3_sd_nan[14];
  assign _06950_ = wt3_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20311" *) wt3_sd_nan[14];
  assign _06951_ = wt3_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20321" *) wt3_sd_nan[15];
  assign _06952_ = wt3_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20331" *) wt3_sd_nan[15];
  assign _06953_ = wt3_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20341" *) wt3_sd_nan[16];
  assign _06954_ = wt3_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20351" *) wt3_sd_nan[16];
  assign _06955_ = wt3_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20361" *) wt3_sd_nan[17];
  assign _06956_ = wt3_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20371" *) wt3_sd_nan[17];
  assign _06957_ = wt3_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20381" *) wt3_sd_nan[18];
  assign _06958_ = wt3_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20391" *) wt3_sd_nan[18];
  assign _06959_ = wt3_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20401" *) wt3_sd_nan[19];
  assign _06960_ = wt3_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20411" *) wt3_sd_nan[19];
  assign _06961_ = wt3_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20421" *) wt3_sd_nan[20];
  assign _06962_ = wt3_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20431" *) wt3_sd_nan[20];
  assign _06963_ = wt3_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20441" *) wt3_sd_nan[21];
  assign _06964_ = wt3_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20451" *) wt3_sd_nan[21];
  assign _06965_ = wt3_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20461" *) wt3_sd_nan[22];
  assign _06966_ = wt3_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20471" *) wt3_sd_nan[22];
  assign _06967_ = wt3_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20481" *) wt3_sd_nan[23];
  assign _06968_ = wt3_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20491" *) wt3_sd_nan[23];
  assign _06969_ = wt3_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20501" *) wt3_sd_nan[24];
  assign _06970_ = wt3_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20511" *) wt3_sd_nan[24];
  assign _06971_ = wt3_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20521" *) wt3_sd_nan[25];
  assign _06972_ = wt3_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20531" *) wt3_sd_nan[25];
  assign _06973_ = wt3_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20541" *) wt3_sd_nan[26];
  assign _06974_ = wt3_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20551" *) wt3_sd_nan[26];
  assign _06975_ = wt3_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20561" *) wt3_sd_nan[27];
  assign _06976_ = wt3_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20571" *) wt3_sd_nan[27];
  assign _06977_ = wt3_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20581" *) wt3_sd_nan[28];
  assign _06978_ = wt3_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20591" *) wt3_sd_nan[28];
  assign _06979_ = wt3_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20601" *) wt3_sd_nan[29];
  assign _06980_ = wt3_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20611" *) wt3_sd_nan[29];
  assign _06981_ = wt3_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20621" *) wt3_sd_nan[30];
  assign _06982_ = wt3_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20631" *) wt3_sd_nan[30];
  assign _06983_ = wt3_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20641" *) wt3_sd_nan[31];
  assign _06984_ = wt3_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20651" *) wt3_sd_nan[31];
  assign _06985_ = wt3_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20661" *) wt3_sd_nan[32];
  assign _06986_ = wt3_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20671" *) wt3_sd_nan[32];
  assign _06987_ = wt3_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20681" *) wt3_sd_nan[33];
  assign _06988_ = wt3_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20691" *) wt3_sd_nan[33];
  assign _06989_ = wt3_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20701" *) wt3_sd_nan[34];
  assign _06990_ = wt3_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20711" *) wt3_sd_nan[34];
  assign _06991_ = wt3_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20721" *) wt3_sd_nan[35];
  assign _06992_ = wt3_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20731" *) wt3_sd_nan[35];
  assign _06993_ = wt3_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20741" *) wt3_sd_nan[36];
  assign _06994_ = wt3_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20751" *) wt3_sd_nan[36];
  assign _06995_ = wt3_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20761" *) wt3_sd_nan[37];
  assign _06996_ = wt3_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20771" *) wt3_sd_nan[37];
  assign _06997_ = wt3_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20781" *) wt3_sd_nan[38];
  assign _06998_ = wt3_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20791" *) wt3_sd_nan[38];
  assign _06999_ = wt3_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20801" *) wt3_sd_nan[39];
  assign _07000_ = wt3_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20811" *) wt3_sd_nan[39];
  assign _07001_ = wt3_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20821" *) wt3_sd_nan[40];
  assign _07002_ = wt3_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20831" *) wt3_sd_nan[40];
  assign _07003_ = wt3_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20841" *) wt3_sd_nan[41];
  assign _07004_ = wt3_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20851" *) wt3_sd_nan[41];
  assign _07005_ = wt3_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20861" *) wt3_sd_nan[42];
  assign _07006_ = wt3_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20871" *) wt3_sd_nan[42];
  assign _07007_ = wt3_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20881" *) wt3_sd_nan[43];
  assign _07008_ = wt3_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20891" *) wt3_sd_nan[43];
  assign _07009_ = wt3_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20901" *) wt3_sd_nan[44];
  assign _07010_ = wt3_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20911" *) wt3_sd_nan[44];
  assign _07011_ = wt3_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20921" *) wt3_sd_nan[45];
  assign _07012_ = wt3_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20931" *) wt3_sd_nan[45];
  assign _07013_ = wt3_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20941" *) wt3_sd_nan[46];
  assign _07014_ = wt3_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20951" *) wt3_sd_nan[46];
  assign _07015_ = wt3_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20961" *) wt3_sd_nan[47];
  assign _07016_ = wt3_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20971" *) wt3_sd_nan[47];
  assign _07017_ = wt3_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20981" *) wt3_sd_nan[48];
  assign _07018_ = wt3_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20991" *) wt3_sd_nan[48];
  assign _07019_ = wt3_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21001" *) wt3_sd_nan[49];
  assign _07020_ = wt3_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21011" *) wt3_sd_nan[49];
  assign _07021_ = wt3_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21021" *) wt3_sd_nan[50];
  assign _07022_ = wt3_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21031" *) wt3_sd_nan[50];
  assign _07023_ = wt3_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21041" *) wt3_sd_nan[51];
  assign _07024_ = wt3_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21051" *) wt3_sd_nan[51];
  assign _07025_ = wt3_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21061" *) wt3_sd_nan[52];
  assign _07026_ = wt3_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21071" *) wt3_sd_nan[52];
  assign _07027_ = wt3_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21081" *) wt3_sd_nan[53];
  assign _07028_ = wt3_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21091" *) wt3_sd_nan[53];
  assign _07029_ = wt3_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21101" *) wt3_sd_nan[54];
  assign _07030_ = wt3_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21111" *) wt3_sd_nan[54];
  assign _07031_ = wt3_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21121" *) wt3_sd_nan[55];
  assign _07032_ = wt3_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21131" *) wt3_sd_nan[55];
  assign _07033_ = wt3_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21141" *) wt3_sd_nan[56];
  assign _07034_ = wt3_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21151" *) wt3_sd_nan[56];
  assign _07035_ = wt3_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21161" *) wt3_sd_nan[57];
  assign _07036_ = wt3_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21171" *) wt3_sd_nan[57];
  assign _07037_ = wt3_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21181" *) wt3_sd_nan[58];
  assign _07038_ = wt3_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21191" *) wt3_sd_nan[58];
  assign _07039_ = wt3_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21201" *) wt3_sd_nan[59];
  assign _07040_ = wt3_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21211" *) wt3_sd_nan[59];
  assign _07041_ = wt3_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21221" *) wt3_sd_nan[60];
  assign _07042_ = wt3_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21231" *) wt3_sd_nan[60];
  assign _07043_ = wt3_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21241" *) wt3_sd_nan[61];
  assign _07044_ = wt3_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21251" *) wt3_sd_nan[61];
  assign _07045_ = wt3_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21261" *) wt3_sd_nan[62];
  assign _07046_ = wt3_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21271" *) wt3_sd_nan[62];
  assign _07047_ = wt3_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21281" *) wt3_sd_nan[63];
  assign _07048_ = wt3_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21291" *) wt3_sd_nan[63];
  assign _07049_ = wt4_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21345" *) wt4_sd_nan[0];
  assign _07050_ = wt4_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21355" *) wt4_sd_nan[0];
  assign _07051_ = wt4_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21365" *) wt4_sd_nan[1];
  assign _07052_ = wt4_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21375" *) wt4_sd_nan[1];
  assign _07053_ = wt4_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21385" *) wt4_sd_nan[2];
  assign _07054_ = wt4_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21395" *) wt4_sd_nan[2];
  assign _07055_ = wt4_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21405" *) wt4_sd_nan[3];
  assign _07056_ = wt4_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21415" *) wt4_sd_nan[3];
  assign _07057_ = wt4_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21425" *) wt4_sd_nan[4];
  assign _07058_ = wt4_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21435" *) wt4_sd_nan[4];
  assign _07059_ = wt4_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21445" *) wt4_sd_nan[5];
  assign _07060_ = wt4_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21455" *) wt4_sd_nan[5];
  assign _07061_ = wt4_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21465" *) wt4_sd_nan[6];
  assign _07062_ = wt4_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21475" *) wt4_sd_nan[6];
  assign _07063_ = wt4_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21485" *) wt4_sd_nan[7];
  assign _07064_ = wt4_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21495" *) wt4_sd_nan[7];
  assign _07065_ = wt4_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21505" *) wt4_sd_nan[8];
  assign _07066_ = wt4_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21515" *) wt4_sd_nan[8];
  assign _07067_ = wt4_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21525" *) wt4_sd_nan[9];
  assign _07068_ = wt4_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21535" *) wt4_sd_nan[9];
  assign _07069_ = wt4_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21545" *) wt4_sd_nan[10];
  assign _07070_ = wt4_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21555" *) wt4_sd_nan[10];
  assign _07071_ = wt4_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21565" *) wt4_sd_nan[11];
  assign _07072_ = wt4_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21575" *) wt4_sd_nan[11];
  assign _07073_ = wt4_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21585" *) wt4_sd_nan[12];
  assign _07074_ = wt4_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21595" *) wt4_sd_nan[12];
  assign _07075_ = wt4_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21605" *) wt4_sd_nan[13];
  assign _07076_ = wt4_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21615" *) wt4_sd_nan[13];
  assign _07077_ = wt4_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21625" *) wt4_sd_nan[14];
  assign _07078_ = wt4_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21635" *) wt4_sd_nan[14];
  assign _07079_ = wt4_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21645" *) wt4_sd_nan[15];
  assign _07080_ = wt4_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21655" *) wt4_sd_nan[15];
  assign _07081_ = wt4_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21665" *) wt4_sd_nan[16];
  assign _07082_ = wt4_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21675" *) wt4_sd_nan[16];
  assign _07083_ = wt4_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21685" *) wt4_sd_nan[17];
  assign _07084_ = wt4_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21695" *) wt4_sd_nan[17];
  assign _07085_ = wt4_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21705" *) wt4_sd_nan[18];
  assign _07086_ = wt4_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21715" *) wt4_sd_nan[18];
  assign _07087_ = wt4_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21725" *) wt4_sd_nan[19];
  assign _07088_ = wt4_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21735" *) wt4_sd_nan[19];
  assign _07089_ = wt4_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21745" *) wt4_sd_nan[20];
  assign _07090_ = wt4_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21755" *) wt4_sd_nan[20];
  assign _07091_ = wt4_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21765" *) wt4_sd_nan[21];
  assign _07092_ = wt4_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21775" *) wt4_sd_nan[21];
  assign _07093_ = wt4_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21785" *) wt4_sd_nan[22];
  assign _07094_ = wt4_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21795" *) wt4_sd_nan[22];
  assign _07095_ = wt4_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21805" *) wt4_sd_nan[23];
  assign _07096_ = wt4_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21815" *) wt4_sd_nan[23];
  assign _07097_ = wt4_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21825" *) wt4_sd_nan[24];
  assign _07098_ = wt4_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21835" *) wt4_sd_nan[24];
  assign _07099_ = wt4_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21845" *) wt4_sd_nan[25];
  assign _07100_ = wt4_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21855" *) wt4_sd_nan[25];
  assign _07101_ = wt4_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21865" *) wt4_sd_nan[26];
  assign _07102_ = wt4_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21875" *) wt4_sd_nan[26];
  assign _07103_ = wt4_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21885" *) wt4_sd_nan[27];
  assign _07104_ = wt4_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21895" *) wt4_sd_nan[27];
  assign _07105_ = wt4_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21905" *) wt4_sd_nan[28];
  assign _07106_ = wt4_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21915" *) wt4_sd_nan[28];
  assign _07107_ = wt4_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21925" *) wt4_sd_nan[29];
  assign _07108_ = wt4_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21935" *) wt4_sd_nan[29];
  assign _07109_ = wt4_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21945" *) wt4_sd_nan[30];
  assign _07110_ = wt4_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21955" *) wt4_sd_nan[30];
  assign _07111_ = wt4_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21965" *) wt4_sd_nan[31];
  assign _07112_ = wt4_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21975" *) wt4_sd_nan[31];
  assign _07113_ = wt4_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21985" *) wt4_sd_nan[32];
  assign _07114_ = wt4_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21995" *) wt4_sd_nan[32];
  assign _07115_ = wt4_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22005" *) wt4_sd_nan[33];
  assign _07116_ = wt4_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22015" *) wt4_sd_nan[33];
  assign _07117_ = wt4_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22025" *) wt4_sd_nan[34];
  assign _07118_ = wt4_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22035" *) wt4_sd_nan[34];
  assign _07119_ = wt4_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22045" *) wt4_sd_nan[35];
  assign _07120_ = wt4_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22055" *) wt4_sd_nan[35];
  assign _07121_ = wt4_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22065" *) wt4_sd_nan[36];
  assign _07122_ = wt4_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22075" *) wt4_sd_nan[36];
  assign _07123_ = wt4_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22085" *) wt4_sd_nan[37];
  assign _07124_ = wt4_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22095" *) wt4_sd_nan[37];
  assign _07125_ = wt4_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22105" *) wt4_sd_nan[38];
  assign _07126_ = wt4_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22115" *) wt4_sd_nan[38];
  assign _07127_ = wt4_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22125" *) wt4_sd_nan[39];
  assign _07128_ = wt4_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22135" *) wt4_sd_nan[39];
  assign _07129_ = wt4_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22145" *) wt4_sd_nan[40];
  assign _07130_ = wt4_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22155" *) wt4_sd_nan[40];
  assign _07131_ = wt4_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22165" *) wt4_sd_nan[41];
  assign _07132_ = wt4_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22175" *) wt4_sd_nan[41];
  assign _07133_ = wt4_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22185" *) wt4_sd_nan[42];
  assign _07134_ = wt4_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22195" *) wt4_sd_nan[42];
  assign _07135_ = wt4_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22205" *) wt4_sd_nan[43];
  assign _07136_ = wt4_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22215" *) wt4_sd_nan[43];
  assign _07137_ = wt4_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22225" *) wt4_sd_nan[44];
  assign _07138_ = wt4_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22235" *) wt4_sd_nan[44];
  assign _07139_ = wt4_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22245" *) wt4_sd_nan[45];
  assign _07140_ = wt4_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22255" *) wt4_sd_nan[45];
  assign _07141_ = wt4_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22265" *) wt4_sd_nan[46];
  assign _07142_ = wt4_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22275" *) wt4_sd_nan[46];
  assign _07143_ = wt4_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22285" *) wt4_sd_nan[47];
  assign _07144_ = wt4_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22295" *) wt4_sd_nan[47];
  assign _07145_ = wt4_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22305" *) wt4_sd_nan[48];
  assign _07146_ = wt4_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22315" *) wt4_sd_nan[48];
  assign _07147_ = wt4_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22325" *) wt4_sd_nan[49];
  assign _07148_ = wt4_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22335" *) wt4_sd_nan[49];
  assign _07149_ = wt4_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22345" *) wt4_sd_nan[50];
  assign _07150_ = wt4_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22355" *) wt4_sd_nan[50];
  assign _07151_ = wt4_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22365" *) wt4_sd_nan[51];
  assign _07152_ = wt4_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22375" *) wt4_sd_nan[51];
  assign _07153_ = wt4_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22385" *) wt4_sd_nan[52];
  assign _07154_ = wt4_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22395" *) wt4_sd_nan[52];
  assign _07155_ = wt4_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22405" *) wt4_sd_nan[53];
  assign _07156_ = wt4_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22415" *) wt4_sd_nan[53];
  assign _07157_ = wt4_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22425" *) wt4_sd_nan[54];
  assign _07158_ = wt4_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22435" *) wt4_sd_nan[54];
  assign _07159_ = wt4_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22445" *) wt4_sd_nan[55];
  assign _07160_ = wt4_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22455" *) wt4_sd_nan[55];
  assign _07161_ = wt4_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22465" *) wt4_sd_nan[56];
  assign _07162_ = wt4_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22475" *) wt4_sd_nan[56];
  assign _07163_ = wt4_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22485" *) wt4_sd_nan[57];
  assign _07164_ = wt4_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22495" *) wt4_sd_nan[57];
  assign _07165_ = wt4_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22505" *) wt4_sd_nan[58];
  assign _07166_ = wt4_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22515" *) wt4_sd_nan[58];
  assign _07167_ = wt4_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22525" *) wt4_sd_nan[59];
  assign _07168_ = wt4_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22535" *) wt4_sd_nan[59];
  assign _07169_ = wt4_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22545" *) wt4_sd_nan[60];
  assign _07170_ = wt4_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22555" *) wt4_sd_nan[60];
  assign _07171_ = wt4_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22565" *) wt4_sd_nan[61];
  assign _07172_ = wt4_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22575" *) wt4_sd_nan[61];
  assign _07173_ = wt4_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22585" *) wt4_sd_nan[62];
  assign _07174_ = wt4_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22595" *) wt4_sd_nan[62];
  assign _07175_ = wt4_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22605" *) wt4_sd_nan[63];
  assign _07176_ = wt4_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22615" *) wt4_sd_nan[63];
  assign _07177_ = wt5_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22669" *) wt5_sd_nan[0];
  assign _07178_ = wt5_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22679" *) wt5_sd_nan[0];
  assign _07179_ = wt5_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22689" *) wt5_sd_nan[1];
  assign _07180_ = wt5_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22699" *) wt5_sd_nan[1];
  assign _07181_ = wt5_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22709" *) wt5_sd_nan[2];
  assign _07182_ = wt5_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22719" *) wt5_sd_nan[2];
  assign _07183_ = wt5_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22729" *) wt5_sd_nan[3];
  assign _07184_ = wt5_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22739" *) wt5_sd_nan[3];
  assign _07185_ = wt5_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22749" *) wt5_sd_nan[4];
  assign _07186_ = wt5_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22759" *) wt5_sd_nan[4];
  assign _07187_ = wt5_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22769" *) wt5_sd_nan[5];
  assign _07188_ = wt5_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22779" *) wt5_sd_nan[5];
  assign _07189_ = wt5_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22789" *) wt5_sd_nan[6];
  assign _07190_ = wt5_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22799" *) wt5_sd_nan[6];
  assign _07191_ = wt5_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22809" *) wt5_sd_nan[7];
  assign _07192_ = wt5_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22819" *) wt5_sd_nan[7];
  assign _07193_ = wt5_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22829" *) wt5_sd_nan[8];
  assign _07194_ = wt5_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22839" *) wt5_sd_nan[8];
  assign _07195_ = wt5_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22849" *) wt5_sd_nan[9];
  assign _07196_ = wt5_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22859" *) wt5_sd_nan[9];
  assign _07197_ = wt5_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22869" *) wt5_sd_nan[10];
  assign _07198_ = wt5_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22879" *) wt5_sd_nan[10];
  assign _07199_ = wt5_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22889" *) wt5_sd_nan[11];
  assign _07200_ = wt5_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22899" *) wt5_sd_nan[11];
  assign _07201_ = wt5_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22909" *) wt5_sd_nan[12];
  assign _07202_ = wt5_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22919" *) wt5_sd_nan[12];
  assign _07203_ = wt5_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22929" *) wt5_sd_nan[13];
  assign _07204_ = wt5_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22939" *) wt5_sd_nan[13];
  assign _07205_ = wt5_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22949" *) wt5_sd_nan[14];
  assign _07206_ = wt5_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22959" *) wt5_sd_nan[14];
  assign _07207_ = wt5_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22969" *) wt5_sd_nan[15];
  assign _07208_ = wt5_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22979" *) wt5_sd_nan[15];
  assign _07209_ = wt5_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22989" *) wt5_sd_nan[16];
  assign _07210_ = wt5_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22999" *) wt5_sd_nan[16];
  assign _07211_ = wt5_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23009" *) wt5_sd_nan[17];
  assign _07212_ = wt5_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23019" *) wt5_sd_nan[17];
  assign _07213_ = wt5_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23029" *) wt5_sd_nan[18];
  assign _07214_ = wt5_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23039" *) wt5_sd_nan[18];
  assign _07215_ = wt5_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23049" *) wt5_sd_nan[19];
  assign _07216_ = wt5_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23059" *) wt5_sd_nan[19];
  assign _07217_ = wt5_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23069" *) wt5_sd_nan[20];
  assign _07218_ = wt5_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23079" *) wt5_sd_nan[20];
  assign _07219_ = wt5_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23089" *) wt5_sd_nan[21];
  assign _07220_ = wt5_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23099" *) wt5_sd_nan[21];
  assign _07221_ = wt5_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23109" *) wt5_sd_nan[22];
  assign _07222_ = wt5_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23119" *) wt5_sd_nan[22];
  assign _07223_ = wt5_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23129" *) wt5_sd_nan[23];
  assign _07224_ = wt5_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23139" *) wt5_sd_nan[23];
  assign _07225_ = wt5_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23149" *) wt5_sd_nan[24];
  assign _07226_ = wt5_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23159" *) wt5_sd_nan[24];
  assign _07227_ = wt5_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23169" *) wt5_sd_nan[25];
  assign _07228_ = wt5_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23179" *) wt5_sd_nan[25];
  assign _07229_ = wt5_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23189" *) wt5_sd_nan[26];
  assign _07230_ = wt5_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23199" *) wt5_sd_nan[26];
  assign _07231_ = wt5_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23209" *) wt5_sd_nan[27];
  assign _07232_ = wt5_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23219" *) wt5_sd_nan[27];
  assign _07233_ = wt5_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23229" *) wt5_sd_nan[28];
  assign _07234_ = wt5_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23239" *) wt5_sd_nan[28];
  assign _07235_ = wt5_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23249" *) wt5_sd_nan[29];
  assign _07236_ = wt5_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23259" *) wt5_sd_nan[29];
  assign _07237_ = wt5_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23269" *) wt5_sd_nan[30];
  assign _07238_ = wt5_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23279" *) wt5_sd_nan[30];
  assign _07239_ = wt5_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23289" *) wt5_sd_nan[31];
  assign _07240_ = wt5_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23299" *) wt5_sd_nan[31];
  assign _07241_ = wt5_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23309" *) wt5_sd_nan[32];
  assign _07242_ = wt5_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23319" *) wt5_sd_nan[32];
  assign _07243_ = wt5_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23329" *) wt5_sd_nan[33];
  assign _07244_ = wt5_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23339" *) wt5_sd_nan[33];
  assign _07245_ = wt5_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23349" *) wt5_sd_nan[34];
  assign _07246_ = wt5_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23359" *) wt5_sd_nan[34];
  assign _07247_ = wt5_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23369" *) wt5_sd_nan[35];
  assign _07248_ = wt5_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23379" *) wt5_sd_nan[35];
  assign _07249_ = wt5_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23389" *) wt5_sd_nan[36];
  assign _07250_ = wt5_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23399" *) wt5_sd_nan[36];
  assign _07251_ = wt5_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23409" *) wt5_sd_nan[37];
  assign _07252_ = wt5_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23419" *) wt5_sd_nan[37];
  assign _07253_ = wt5_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23429" *) wt5_sd_nan[38];
  assign _07254_ = wt5_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23439" *) wt5_sd_nan[38];
  assign _07255_ = wt5_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23449" *) wt5_sd_nan[39];
  assign _07256_ = wt5_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23459" *) wt5_sd_nan[39];
  assign _07257_ = wt5_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23469" *) wt5_sd_nan[40];
  assign _07258_ = wt5_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23479" *) wt5_sd_nan[40];
  assign _07259_ = wt5_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23489" *) wt5_sd_nan[41];
  assign _07260_ = wt5_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23499" *) wt5_sd_nan[41];
  assign _07261_ = wt5_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23509" *) wt5_sd_nan[42];
  assign _07262_ = wt5_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23519" *) wt5_sd_nan[42];
  assign _07263_ = wt5_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23529" *) wt5_sd_nan[43];
  assign _07264_ = wt5_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23539" *) wt5_sd_nan[43];
  assign _07265_ = wt5_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23549" *) wt5_sd_nan[44];
  assign _07266_ = wt5_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23559" *) wt5_sd_nan[44];
  assign _07267_ = wt5_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23569" *) wt5_sd_nan[45];
  assign _07268_ = wt5_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23579" *) wt5_sd_nan[45];
  assign _07269_ = wt5_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23589" *) wt5_sd_nan[46];
  assign _07270_ = wt5_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23599" *) wt5_sd_nan[46];
  assign _07271_ = wt5_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23609" *) wt5_sd_nan[47];
  assign _07272_ = wt5_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23619" *) wt5_sd_nan[47];
  assign _07273_ = wt5_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23629" *) wt5_sd_nan[48];
  assign _07274_ = wt5_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23639" *) wt5_sd_nan[48];
  assign _07275_ = wt5_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23649" *) wt5_sd_nan[49];
  assign _07276_ = wt5_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23659" *) wt5_sd_nan[49];
  assign _07277_ = wt5_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23669" *) wt5_sd_nan[50];
  assign _07278_ = wt5_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23679" *) wt5_sd_nan[50];
  assign _07279_ = wt5_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23689" *) wt5_sd_nan[51];
  assign _07280_ = wt5_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23699" *) wt5_sd_nan[51];
  assign _07281_ = wt5_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23709" *) wt5_sd_nan[52];
  assign _07282_ = wt5_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23719" *) wt5_sd_nan[52];
  assign _07283_ = wt5_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23729" *) wt5_sd_nan[53];
  assign _07284_ = wt5_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23739" *) wt5_sd_nan[53];
  assign _07285_ = wt5_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23749" *) wt5_sd_nan[54];
  assign _07286_ = wt5_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23759" *) wt5_sd_nan[54];
  assign _07287_ = wt5_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23769" *) wt5_sd_nan[55];
  assign _07288_ = wt5_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23779" *) wt5_sd_nan[55];
  assign _07289_ = wt5_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23789" *) wt5_sd_nan[56];
  assign _07290_ = wt5_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23799" *) wt5_sd_nan[56];
  assign _07291_ = wt5_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23809" *) wt5_sd_nan[57];
  assign _07292_ = wt5_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23819" *) wt5_sd_nan[57];
  assign _07293_ = wt5_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23829" *) wt5_sd_nan[58];
  assign _07294_ = wt5_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23839" *) wt5_sd_nan[58];
  assign _07295_ = wt5_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23849" *) wt5_sd_nan[59];
  assign _07296_ = wt5_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23859" *) wt5_sd_nan[59];
  assign _07297_ = wt5_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23869" *) wt5_sd_nan[60];
  assign _07298_ = wt5_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23879" *) wt5_sd_nan[60];
  assign _07299_ = wt5_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23889" *) wt5_sd_nan[61];
  assign _07300_ = wt5_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23899" *) wt5_sd_nan[61];
  assign _07301_ = wt5_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23909" *) wt5_sd_nan[62];
  assign _07302_ = wt5_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23919" *) wt5_sd_nan[62];
  assign _07303_ = wt5_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23929" *) wt5_sd_nan[63];
  assign _07304_ = wt5_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23939" *) wt5_sd_nan[63];
  assign _07305_ = wt6_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23993" *) wt6_sd_nan[0];
  assign _07306_ = wt6_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24003" *) wt6_sd_nan[0];
  assign _07307_ = wt6_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24013" *) wt6_sd_nan[1];
  assign _07308_ = wt6_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24023" *) wt6_sd_nan[1];
  assign _07309_ = wt6_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24033" *) wt6_sd_nan[2];
  assign _07310_ = wt6_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24043" *) wt6_sd_nan[2];
  assign _07311_ = wt6_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24053" *) wt6_sd_nan[3];
  assign _07312_ = wt6_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24063" *) wt6_sd_nan[3];
  assign _07313_ = wt6_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24073" *) wt6_sd_nan[4];
  assign _07314_ = wt6_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24083" *) wt6_sd_nan[4];
  assign _07315_ = wt6_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24093" *) wt6_sd_nan[5];
  assign _07316_ = wt6_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24103" *) wt6_sd_nan[5];
  assign _07317_ = wt6_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24113" *) wt6_sd_nan[6];
  assign _07318_ = wt6_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24123" *) wt6_sd_nan[6];
  assign _07319_ = wt6_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24133" *) wt6_sd_nan[7];
  assign _07320_ = wt6_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24143" *) wt6_sd_nan[7];
  assign _07321_ = wt6_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24153" *) wt6_sd_nan[8];
  assign _07322_ = wt6_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24163" *) wt6_sd_nan[8];
  assign _07323_ = wt6_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24173" *) wt6_sd_nan[9];
  assign _07324_ = wt6_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24183" *) wt6_sd_nan[9];
  assign _07325_ = wt6_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24193" *) wt6_sd_nan[10];
  assign _07326_ = wt6_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24203" *) wt6_sd_nan[10];
  assign _07327_ = wt6_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24213" *) wt6_sd_nan[11];
  assign _07328_ = wt6_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24223" *) wt6_sd_nan[11];
  assign _07329_ = wt6_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24233" *) wt6_sd_nan[12];
  assign _07330_ = wt6_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24243" *) wt6_sd_nan[12];
  assign _07331_ = wt6_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24253" *) wt6_sd_nan[13];
  assign _07332_ = wt6_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24263" *) wt6_sd_nan[13];
  assign _07333_ = wt6_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24273" *) wt6_sd_nan[14];
  assign _07334_ = wt6_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24283" *) wt6_sd_nan[14];
  assign _07335_ = wt6_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24293" *) wt6_sd_nan[15];
  assign _07336_ = wt6_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24303" *) wt6_sd_nan[15];
  assign _07337_ = wt6_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24313" *) wt6_sd_nan[16];
  assign _07338_ = wt6_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24323" *) wt6_sd_nan[16];
  assign _07339_ = wt6_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24333" *) wt6_sd_nan[17];
  assign _07340_ = wt6_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24343" *) wt6_sd_nan[17];
  assign _07341_ = wt6_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24353" *) wt6_sd_nan[18];
  assign _07342_ = wt6_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24363" *) wt6_sd_nan[18];
  assign _07343_ = wt6_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24373" *) wt6_sd_nan[19];
  assign _07344_ = wt6_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24383" *) wt6_sd_nan[19];
  assign _07345_ = wt6_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24393" *) wt6_sd_nan[20];
  assign _07346_ = wt6_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24403" *) wt6_sd_nan[20];
  assign _07347_ = wt6_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24413" *) wt6_sd_nan[21];
  assign _07348_ = wt6_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24423" *) wt6_sd_nan[21];
  assign _07349_ = wt6_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24433" *) wt6_sd_nan[22];
  assign _07350_ = wt6_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24443" *) wt6_sd_nan[22];
  assign _07351_ = wt6_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24453" *) wt6_sd_nan[23];
  assign _07352_ = wt6_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24463" *) wt6_sd_nan[23];
  assign _07353_ = wt6_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24473" *) wt6_sd_nan[24];
  assign _07354_ = wt6_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24483" *) wt6_sd_nan[24];
  assign _07355_ = wt6_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24493" *) wt6_sd_nan[25];
  assign _07356_ = wt6_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24503" *) wt6_sd_nan[25];
  assign _07357_ = wt6_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24513" *) wt6_sd_nan[26];
  assign _07358_ = wt6_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24523" *) wt6_sd_nan[26];
  assign _07359_ = wt6_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24533" *) wt6_sd_nan[27];
  assign _07360_ = wt6_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24543" *) wt6_sd_nan[27];
  assign _07361_ = wt6_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24553" *) wt6_sd_nan[28];
  assign _07362_ = wt6_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24563" *) wt6_sd_nan[28];
  assign _07363_ = wt6_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24573" *) wt6_sd_nan[29];
  assign _07364_ = wt6_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24583" *) wt6_sd_nan[29];
  assign _07365_ = wt6_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24593" *) wt6_sd_nan[30];
  assign _07366_ = wt6_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24603" *) wt6_sd_nan[30];
  assign _07367_ = wt6_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24613" *) wt6_sd_nan[31];
  assign _07368_ = wt6_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24623" *) wt6_sd_nan[31];
  assign _07369_ = wt6_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24633" *) wt6_sd_nan[32];
  assign _07370_ = wt6_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24643" *) wt6_sd_nan[32];
  assign _07371_ = wt6_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24653" *) wt6_sd_nan[33];
  assign _07372_ = wt6_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24663" *) wt6_sd_nan[33];
  assign _07373_ = wt6_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24673" *) wt6_sd_nan[34];
  assign _07374_ = wt6_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24683" *) wt6_sd_nan[34];
  assign _07375_ = wt6_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24693" *) wt6_sd_nan[35];
  assign _07376_ = wt6_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24703" *) wt6_sd_nan[35];
  assign _07377_ = wt6_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24713" *) wt6_sd_nan[36];
  assign _07378_ = wt6_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24723" *) wt6_sd_nan[36];
  assign _07379_ = wt6_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24733" *) wt6_sd_nan[37];
  assign _07380_ = wt6_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24743" *) wt6_sd_nan[37];
  assign _07381_ = wt6_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24753" *) wt6_sd_nan[38];
  assign _07382_ = wt6_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24763" *) wt6_sd_nan[38];
  assign _07383_ = wt6_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24773" *) wt6_sd_nan[39];
  assign _07384_ = wt6_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24783" *) wt6_sd_nan[39];
  assign _07385_ = wt6_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24793" *) wt6_sd_nan[40];
  assign _07386_ = wt6_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24803" *) wt6_sd_nan[40];
  assign _07387_ = wt6_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24813" *) wt6_sd_nan[41];
  assign _07388_ = wt6_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24823" *) wt6_sd_nan[41];
  assign _07389_ = wt6_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24833" *) wt6_sd_nan[42];
  assign _07390_ = wt6_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24843" *) wt6_sd_nan[42];
  assign _07391_ = wt6_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24853" *) wt6_sd_nan[43];
  assign _07392_ = wt6_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24863" *) wt6_sd_nan[43];
  assign _07393_ = wt6_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24873" *) wt6_sd_nan[44];
  assign _07394_ = wt6_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24883" *) wt6_sd_nan[44];
  assign _07395_ = wt6_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24893" *) wt6_sd_nan[45];
  assign _07396_ = wt6_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24903" *) wt6_sd_nan[45];
  assign _07397_ = wt6_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24913" *) wt6_sd_nan[46];
  assign _07398_ = wt6_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24923" *) wt6_sd_nan[46];
  assign _07399_ = wt6_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24933" *) wt6_sd_nan[47];
  assign _07400_ = wt6_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24943" *) wt6_sd_nan[47];
  assign _07401_ = wt6_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24953" *) wt6_sd_nan[48];
  assign _07402_ = wt6_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24963" *) wt6_sd_nan[48];
  assign _07403_ = wt6_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24973" *) wt6_sd_nan[49];
  assign _07404_ = wt6_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24983" *) wt6_sd_nan[49];
  assign _07405_ = wt6_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24993" *) wt6_sd_nan[50];
  assign _07406_ = wt6_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25003" *) wt6_sd_nan[50];
  assign _07407_ = wt6_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25013" *) wt6_sd_nan[51];
  assign _07408_ = wt6_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25023" *) wt6_sd_nan[51];
  assign _07409_ = wt6_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25033" *) wt6_sd_nan[52];
  assign _07410_ = wt6_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25043" *) wt6_sd_nan[52];
  assign _07411_ = wt6_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25053" *) wt6_sd_nan[53];
  assign _07412_ = wt6_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25063" *) wt6_sd_nan[53];
  assign _07413_ = wt6_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25073" *) wt6_sd_nan[54];
  assign _07414_ = wt6_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25083" *) wt6_sd_nan[54];
  assign _07415_ = wt6_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25093" *) wt6_sd_nan[55];
  assign _07416_ = wt6_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25103" *) wt6_sd_nan[55];
  assign _07417_ = wt6_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25113" *) wt6_sd_nan[56];
  assign _07418_ = wt6_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25123" *) wt6_sd_nan[56];
  assign _07419_ = wt6_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25133" *) wt6_sd_nan[57];
  assign _07420_ = wt6_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25143" *) wt6_sd_nan[57];
  assign _07421_ = wt6_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25153" *) wt6_sd_nan[58];
  assign _07422_ = wt6_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25163" *) wt6_sd_nan[58];
  assign _07423_ = wt6_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25173" *) wt6_sd_nan[59];
  assign _07424_ = wt6_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25183" *) wt6_sd_nan[59];
  assign _07425_ = wt6_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25193" *) wt6_sd_nan[60];
  assign _07426_ = wt6_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25203" *) wt6_sd_nan[60];
  assign _07427_ = wt6_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25213" *) wt6_sd_nan[61];
  assign _07428_ = wt6_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25223" *) wt6_sd_nan[61];
  assign _07429_ = wt6_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25233" *) wt6_sd_nan[62];
  assign _07430_ = wt6_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25243" *) wt6_sd_nan[62];
  assign _07431_ = wt6_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25253" *) wt6_sd_nan[63];
  assign _07432_ = wt6_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25263" *) wt6_sd_nan[63];
  assign _07433_ = wt7_sd_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25317" *) wt7_sd_nan[0];
  assign _07434_ = wt7_sd_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25327" *) wt7_sd_nan[0];
  assign _07435_ = wt7_sd_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25337" *) wt7_sd_nan[1];
  assign _07436_ = wt7_sd_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25347" *) wt7_sd_nan[1];
  assign _07437_ = wt7_sd_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25357" *) wt7_sd_nan[2];
  assign _07438_ = wt7_sd_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25367" *) wt7_sd_nan[2];
  assign _07439_ = wt7_sd_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25377" *) wt7_sd_nan[3];
  assign _07440_ = wt7_sd_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25387" *) wt7_sd_nan[3];
  assign _07441_ = wt7_sd_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25397" *) wt7_sd_nan[4];
  assign _07442_ = wt7_sd_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25407" *) wt7_sd_nan[4];
  assign _07443_ = wt7_sd_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25417" *) wt7_sd_nan[5];
  assign _07444_ = wt7_sd_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25427" *) wt7_sd_nan[5];
  assign _07445_ = wt7_sd_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25437" *) wt7_sd_nan[6];
  assign _07446_ = wt7_sd_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25447" *) wt7_sd_nan[6];
  assign _07447_ = wt7_sd_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25457" *) wt7_sd_nan[7];
  assign _07448_ = wt7_sd_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25467" *) wt7_sd_nan[7];
  assign _07449_ = wt7_sd_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25477" *) wt7_sd_nan[8];
  assign _07450_ = wt7_sd_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25487" *) wt7_sd_nan[8];
  assign _07451_ = wt7_sd_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25497" *) wt7_sd_nan[9];
  assign _07452_ = wt7_sd_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25507" *) wt7_sd_nan[9];
  assign _07453_ = wt7_sd_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25517" *) wt7_sd_nan[10];
  assign _07454_ = wt7_sd_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25527" *) wt7_sd_nan[10];
  assign _07455_ = wt7_sd_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25537" *) wt7_sd_nan[11];
  assign _07456_ = wt7_sd_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25547" *) wt7_sd_nan[11];
  assign _07457_ = wt7_sd_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25557" *) wt7_sd_nan[12];
  assign _07458_ = wt7_sd_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25567" *) wt7_sd_nan[12];
  assign _07459_ = wt7_sd_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25577" *) wt7_sd_nan[13];
  assign _07460_ = wt7_sd_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25587" *) wt7_sd_nan[13];
  assign _07461_ = wt7_sd_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25597" *) wt7_sd_nan[14];
  assign _07462_ = wt7_sd_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25607" *) wt7_sd_nan[14];
  assign _07463_ = wt7_sd_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25617" *) wt7_sd_nan[15];
  assign _07464_ = wt7_sd_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25627" *) wt7_sd_nan[15];
  assign _07465_ = wt7_sd_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25637" *) wt7_sd_nan[16];
  assign _07466_ = wt7_sd_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25647" *) wt7_sd_nan[16];
  assign _07467_ = wt7_sd_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25657" *) wt7_sd_nan[17];
  assign _07468_ = wt7_sd_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25667" *) wt7_sd_nan[17];
  assign _07469_ = wt7_sd_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25677" *) wt7_sd_nan[18];
  assign _07470_ = wt7_sd_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25687" *) wt7_sd_nan[18];
  assign _07471_ = wt7_sd_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25697" *) wt7_sd_nan[19];
  assign _07472_ = wt7_sd_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25707" *) wt7_sd_nan[19];
  assign _07473_ = wt7_sd_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25717" *) wt7_sd_nan[20];
  assign _07474_ = wt7_sd_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25727" *) wt7_sd_nan[20];
  assign _07475_ = wt7_sd_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25737" *) wt7_sd_nan[21];
  assign _07476_ = wt7_sd_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25747" *) wt7_sd_nan[21];
  assign _07477_ = wt7_sd_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25757" *) wt7_sd_nan[22];
  assign _07478_ = wt7_sd_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25767" *) wt7_sd_nan[22];
  assign _07479_ = wt7_sd_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25777" *) wt7_sd_nan[23];
  assign _07480_ = wt7_sd_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25787" *) wt7_sd_nan[23];
  assign _07481_ = wt7_sd_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25797" *) wt7_sd_nan[24];
  assign _07482_ = wt7_sd_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25807" *) wt7_sd_nan[24];
  assign _07483_ = wt7_sd_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25817" *) wt7_sd_nan[25];
  assign _07484_ = wt7_sd_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25827" *) wt7_sd_nan[25];
  assign _07485_ = wt7_sd_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25837" *) wt7_sd_nan[26];
  assign _07486_ = wt7_sd_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25847" *) wt7_sd_nan[26];
  assign _07487_ = wt7_sd_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25857" *) wt7_sd_nan[27];
  assign _07488_ = wt7_sd_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25867" *) wt7_sd_nan[27];
  assign _07489_ = wt7_sd_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25877" *) wt7_sd_nan[28];
  assign _07490_ = wt7_sd_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25887" *) wt7_sd_nan[28];
  assign _07491_ = wt7_sd_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25897" *) wt7_sd_nan[29];
  assign _07492_ = wt7_sd_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25907" *) wt7_sd_nan[29];
  assign _07493_ = wt7_sd_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25917" *) wt7_sd_nan[30];
  assign _07494_ = wt7_sd_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25927" *) wt7_sd_nan[30];
  assign _07495_ = wt7_sd_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25937" *) wt7_sd_nan[31];
  assign _07496_ = wt7_sd_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25947" *) wt7_sd_nan[31];
  assign _07497_ = wt7_sd_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25957" *) wt7_sd_nan[32];
  assign _07498_ = wt7_sd_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25967" *) wt7_sd_nan[32];
  assign _07499_ = wt7_sd_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25977" *) wt7_sd_nan[33];
  assign _07500_ = wt7_sd_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25987" *) wt7_sd_nan[33];
  assign _07501_ = wt7_sd_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25997" *) wt7_sd_nan[34];
  assign _07502_ = wt7_sd_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26007" *) wt7_sd_nan[34];
  assign _07503_ = wt7_sd_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26017" *) wt7_sd_nan[35];
  assign _07504_ = wt7_sd_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26027" *) wt7_sd_nan[35];
  assign _07505_ = wt7_sd_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26037" *) wt7_sd_nan[36];
  assign _07506_ = wt7_sd_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26047" *) wt7_sd_nan[36];
  assign _07507_ = wt7_sd_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26057" *) wt7_sd_nan[37];
  assign _07508_ = wt7_sd_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26067" *) wt7_sd_nan[37];
  assign _07509_ = wt7_sd_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26077" *) wt7_sd_nan[38];
  assign _07510_ = wt7_sd_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26087" *) wt7_sd_nan[38];
  assign _07511_ = wt7_sd_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26097" *) wt7_sd_nan[39];
  assign _07512_ = wt7_sd_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26107" *) wt7_sd_nan[39];
  assign _07513_ = wt7_sd_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26117" *) wt7_sd_nan[40];
  assign _07514_ = wt7_sd_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26127" *) wt7_sd_nan[40];
  assign _07515_ = wt7_sd_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26137" *) wt7_sd_nan[41];
  assign _07516_ = wt7_sd_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26147" *) wt7_sd_nan[41];
  assign _07517_ = wt7_sd_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26157" *) wt7_sd_nan[42];
  assign _07518_ = wt7_sd_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26167" *) wt7_sd_nan[42];
  assign _07519_ = wt7_sd_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26177" *) wt7_sd_nan[43];
  assign _07520_ = wt7_sd_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26187" *) wt7_sd_nan[43];
  assign _07521_ = wt7_sd_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26197" *) wt7_sd_nan[44];
  assign _07522_ = wt7_sd_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26207" *) wt7_sd_nan[44];
  assign _07523_ = wt7_sd_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26217" *) wt7_sd_nan[45];
  assign _07524_ = wt7_sd_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26227" *) wt7_sd_nan[45];
  assign _07525_ = wt7_sd_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26237" *) wt7_sd_nan[46];
  assign _07526_ = wt7_sd_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26247" *) wt7_sd_nan[46];
  assign _07527_ = wt7_sd_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26257" *) wt7_sd_nan[47];
  assign _07528_ = wt7_sd_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26267" *) wt7_sd_nan[47];
  assign _07529_ = wt7_sd_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26277" *) wt7_sd_nan[48];
  assign _07530_ = wt7_sd_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26287" *) wt7_sd_nan[48];
  assign _07531_ = wt7_sd_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26297" *) wt7_sd_nan[49];
  assign _07532_ = wt7_sd_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26307" *) wt7_sd_nan[49];
  assign _07533_ = wt7_sd_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26317" *) wt7_sd_nan[50];
  assign _07534_ = wt7_sd_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26327" *) wt7_sd_nan[50];
  assign _07535_ = wt7_sd_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26337" *) wt7_sd_nan[51];
  assign _07536_ = wt7_sd_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26347" *) wt7_sd_nan[51];
  assign _07537_ = wt7_sd_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26357" *) wt7_sd_nan[52];
  assign _07538_ = wt7_sd_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26367" *) wt7_sd_nan[52];
  assign _07539_ = wt7_sd_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26377" *) wt7_sd_nan[53];
  assign _07540_ = wt7_sd_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26387" *) wt7_sd_nan[53];
  assign _07541_ = wt7_sd_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26397" *) wt7_sd_nan[54];
  assign _07542_ = wt7_sd_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26407" *) wt7_sd_nan[54];
  assign _07543_ = wt7_sd_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26417" *) wt7_sd_nan[55];
  assign _07544_ = wt7_sd_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26427" *) wt7_sd_nan[55];
  assign _07545_ = wt7_sd_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26437" *) wt7_sd_nan[56];
  assign _07546_ = wt7_sd_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26447" *) wt7_sd_nan[56];
  assign _07547_ = wt7_sd_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26457" *) wt7_sd_nan[57];
  assign _07548_ = wt7_sd_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26467" *) wt7_sd_nan[57];
  assign _07549_ = wt7_sd_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26477" *) wt7_sd_nan[58];
  assign _07550_ = wt7_sd_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26487" *) wt7_sd_nan[58];
  assign _07551_ = wt7_sd_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26497" *) wt7_sd_nan[59];
  assign _07552_ = wt7_sd_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26507" *) wt7_sd_nan[59];
  assign _07553_ = wt7_sd_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26517" *) wt7_sd_nan[60];
  assign _07554_ = wt7_sd_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26527" *) wt7_sd_nan[60];
  assign _07555_ = wt7_sd_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26537" *) wt7_sd_nan[61];
  assign _07556_ = wt7_sd_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26547" *) wt7_sd_nan[61];
  assign _07557_ = wt7_sd_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26557" *) wt7_sd_nan[62];
  assign _07558_ = wt7_sd_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26567" *) wt7_sd_nan[62];
  assign _07559_ = wt7_sd_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26577" *) wt7_sd_nan[63];
  assign _07560_ = wt7_sd_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26587" *) wt7_sd_nan[63];
  assign _07561_ = { in_dat_data_fp16_63, in_dat_data_fp16_62, in_dat_data_fp16_61, in_dat_data_fp16_60, in_dat_data_fp16_59, in_dat_data_fp16_58, in_dat_data_fp16_57, in_dat_data_fp16_56, in_dat_data_fp16_55, in_dat_data_fp16_54, in_dat_data_fp16_53, in_dat_data_fp16_52, in_dat_data_fp16_51, in_dat_data_fp16_50, in_dat_data_fp16_49, in_dat_data_fp16_48, in_dat_data_fp16_47, in_dat_data_fp16_46, in_dat_data_fp16_45, in_dat_data_fp16_44, in_dat_data_fp16_43, in_dat_data_fp16_42, in_dat_data_fp16_41, in_dat_data_fp16_40, in_dat_data_fp16_39, in_dat_data_fp16_38, in_dat_data_fp16_37, in_dat_data_fp16_36, in_dat_data_fp16_35, in_dat_data_fp16_34, in_dat_data_fp16_33, in_dat_data_fp16_32, in_dat_data_fp16_31, in_dat_data_fp16_30, in_dat_data_fp16_29, in_dat_data_fp16_28, in_dat_data_fp16_27, in_dat_data_fp16_26, in_dat_data_fp16_25, in_dat_data_fp16_24, in_dat_data_fp16_23, in_dat_data_fp16_22, in_dat_data_fp16_21, in_dat_data_fp16_20, in_dat_data_fp16_19, in_dat_data_fp16_18, in_dat_data_fp16_17, in_dat_data_fp16_16, in_dat_data_fp16_15, in_dat_data_fp16_14, in_dat_data_fp16_13, in_dat_data_fp16_12, in_dat_data_fp16_11, in_dat_data_fp16_10, in_dat_data_fp16_9, in_dat_data_fp16_8, in_dat_data_fp16_7, in_dat_data_fp16_6, in_dat_data_fp16_5, in_dat_data_fp16_4, in_dat_data_fp16_3, in_dat_data_fp16_2, in_dat_data_fp16_1, in_dat_data_fp16_0 } | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29032" *) { in_dat_data_int8_63, in_dat_data_int8_62, in_dat_data_int8_61, in_dat_data_int8_60, in_dat_data_int8_59, in_dat_data_int8_58, in_dat_data_int8_57, in_dat_data_int8_56, in_dat_data_int8_55, in_dat_data_int8_54, in_dat_data_int8_53, in_dat_data_int8_52, in_dat_data_int8_51, in_dat_data_int8_50, in_dat_data_int8_49, in_dat_data_int8_48, in_dat_data_int8_47, in_dat_data_int8_46, in_dat_data_int8_45, in_dat_data_int8_44, in_dat_data_int8_43, in_dat_data_int8_42, in_dat_data_int8_41, in_dat_data_int8_40, in_dat_data_int8_39, in_dat_data_int8_38, in_dat_data_int8_37, in_dat_data_int8_36, in_dat_data_int8_35, in_dat_data_int8_34, in_dat_data_int8_33, in_dat_data_int8_32, in_dat_data_int8_31, in_dat_data_int8_30, in_dat_data_int8_29, in_dat_data_int8_28, in_dat_data_int8_27, in_dat_data_int8_26, in_dat_data_int8_25, in_dat_data_int8_24, in_dat_data_int8_23, in_dat_data_int8_22, in_dat_data_int8_21, in_dat_data_int8_20, in_dat_data_int8_19, in_dat_data_int8_18, in_dat_data_int8_17, in_dat_data_int8_16, in_dat_data_int8_15, in_dat_data_int8_14, in_dat_data_int8_13, in_dat_data_int8_12, in_dat_data_int8_11, in_dat_data_int8_10, in_dat_data_int8_9, in_dat_data_int8_8, in_dat_data_int8_7, in_dat_data_int8_6, in_dat_data_int8_5, in_dat_data_int8_4, in_dat_data_int8_3, in_dat_data_int8_2, in_dat_data_int8_1, in_dat_data_int8_0 };
  assign dat_pre_data_w = _07561_ | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29032" *) { in_dat_data_int16_63, in_dat_data_int16_62, in_dat_data_int16_61, in_dat_data_int16_60, in_dat_data_int16_59, in_dat_data_int16_58, in_dat_data_int16_57, in_dat_data_int16_56, in_dat_data_int16_55, in_dat_data_int16_54, in_dat_data_int16_53, in_dat_data_int16_52, in_dat_data_int16_51, in_dat_data_int16_50, in_dat_data_int16_49, in_dat_data_int16_48, in_dat_data_int16_47, in_dat_data_int16_46, in_dat_data_int16_45, in_dat_data_int16_44, in_dat_data_int16_43, in_dat_data_int16_42, in_dat_data_int16_41, in_dat_data_int16_40, in_dat_data_int16_39, in_dat_data_int16_38, in_dat_data_int16_37, in_dat_data_int16_36, in_dat_data_int16_35, in_dat_data_int16_34, in_dat_data_int16_33, in_dat_data_int16_32, in_dat_data_int16_31, in_dat_data_int16_30, in_dat_data_int16_29, in_dat_data_int16_28, in_dat_data_int16_27, in_dat_data_int16_26, in_dat_data_int16_25, in_dat_data_int16_24, in_dat_data_int16_23, in_dat_data_int16_22, in_dat_data_int16_21, in_dat_data_int16_20, in_dat_data_int16_19, in_dat_data_int16_18, in_dat_data_int16_17, in_dat_data_int16_16, in_dat_data_int16_15, in_dat_data_int16_14, in_dat_data_int16_13, in_dat_data_int16_12, in_dat_data_int16_11, in_dat_data_int16_10, in_dat_data_int16_9, in_dat_data_int16_8, in_dat_data_int16_7, in_dat_data_int16_6, in_dat_data_int16_5, in_dat_data_int16_4, in_dat_data_int16_3, in_dat_data_int16_2, in_dat_data_int16_1, in_dat_data_int16_0 };
  assign _07562_ = dat_pre_nz_w[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29086" *) in_dat_nan[0];
  assign _07563_ = dat_pre_nz_w[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29096" *) in_dat_nan[0];
  assign _07564_ = dat_pre_nz_w[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29106" *) in_dat_nan[1];
  assign _07565_ = dat_pre_nz_w[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29116" *) in_dat_nan[1];
  assign _07566_ = dat_pre_nz_w[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29126" *) in_dat_nan[2];
  assign _07567_ = dat_pre_nz_w[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29136" *) in_dat_nan[2];
  assign _07568_ = dat_pre_nz_w[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29146" *) in_dat_nan[3];
  assign _07569_ = dat_pre_nz_w[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29156" *) in_dat_nan[3];
  assign _07570_ = dat_pre_nz_w[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29166" *) in_dat_nan[4];
  assign _07571_ = dat_pre_nz_w[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29176" *) in_dat_nan[4];
  assign _07572_ = dat_pre_nz_w[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29186" *) in_dat_nan[5];
  assign _07573_ = dat_pre_nz_w[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29196" *) in_dat_nan[5];
  assign _07574_ = dat_pre_nz_w[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29206" *) in_dat_nan[6];
  assign _07575_ = dat_pre_nz_w[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29216" *) in_dat_nan[6];
  assign _07576_ = dat_pre_nz_w[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29226" *) in_dat_nan[7];
  assign _07577_ = dat_pre_nz_w[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29236" *) in_dat_nan[7];
  assign _07578_ = dat_pre_nz_w[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29246" *) in_dat_nan[8];
  assign _07579_ = dat_pre_nz_w[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29256" *) in_dat_nan[8];
  assign _07580_ = dat_pre_nz_w[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29266" *) in_dat_nan[9];
  assign _07581_ = dat_pre_nz_w[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29276" *) in_dat_nan[9];
  assign _07582_ = dat_pre_nz_w[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29286" *) in_dat_nan[10];
  assign _07583_ = dat_pre_nz_w[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29296" *) in_dat_nan[10];
  assign _07584_ = dat_pre_nz_w[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29306" *) in_dat_nan[11];
  assign _07585_ = dat_pre_nz_w[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29316" *) in_dat_nan[11];
  assign _07586_ = dat_pre_nz_w[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29326" *) in_dat_nan[12];
  assign _07587_ = dat_pre_nz_w[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29336" *) in_dat_nan[12];
  assign _07588_ = dat_pre_nz_w[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29346" *) in_dat_nan[13];
  assign _07589_ = dat_pre_nz_w[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29356" *) in_dat_nan[13];
  assign _07590_ = dat_pre_nz_w[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29366" *) in_dat_nan[14];
  assign _07591_ = dat_pre_nz_w[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29376" *) in_dat_nan[14];
  assign _07592_ = dat_pre_nz_w[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29386" *) in_dat_nan[15];
  assign _07593_ = dat_pre_nz_w[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29396" *) in_dat_nan[15];
  assign _07594_ = dat_pre_nz_w[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29406" *) in_dat_nan[16];
  assign _07595_ = dat_pre_nz_w[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29416" *) in_dat_nan[16];
  assign _07596_ = dat_pre_nz_w[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29426" *) in_dat_nan[17];
  assign _07597_ = dat_pre_nz_w[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29436" *) in_dat_nan[17];
  assign _07598_ = dat_pre_nz_w[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29446" *) in_dat_nan[18];
  assign _07599_ = dat_pre_nz_w[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29456" *) in_dat_nan[18];
  assign _07600_ = dat_pre_nz_w[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29466" *) in_dat_nan[19];
  assign _07601_ = dat_pre_nz_w[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29476" *) in_dat_nan[19];
  assign _07602_ = dat_pre_nz_w[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29486" *) in_dat_nan[20];
  assign _07603_ = dat_pre_nz_w[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29496" *) in_dat_nan[20];
  assign _07604_ = dat_pre_nz_w[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29506" *) in_dat_nan[21];
  assign _07605_ = dat_pre_nz_w[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29516" *) in_dat_nan[21];
  assign _07606_ = dat_pre_nz_w[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29526" *) in_dat_nan[22];
  assign _07607_ = dat_pre_nz_w[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29536" *) in_dat_nan[22];
  assign _07608_ = dat_pre_nz_w[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29546" *) in_dat_nan[23];
  assign _07609_ = dat_pre_nz_w[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29556" *) in_dat_nan[23];
  assign _07610_ = dat_pre_nz_w[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29566" *) in_dat_nan[24];
  assign _07611_ = dat_pre_nz_w[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29576" *) in_dat_nan[24];
  assign _07612_ = dat_pre_nz_w[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29586" *) in_dat_nan[25];
  assign _07613_ = dat_pre_nz_w[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29596" *) in_dat_nan[25];
  assign _07614_ = dat_pre_nz_w[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29606" *) in_dat_nan[26];
  assign _07615_ = dat_pre_nz_w[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29616" *) in_dat_nan[26];
  assign _07616_ = dat_pre_nz_w[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29626" *) in_dat_nan[27];
  assign _07617_ = dat_pre_nz_w[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29636" *) in_dat_nan[27];
  assign _07618_ = dat_pre_nz_w[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29646" *) in_dat_nan[28];
  assign _07619_ = dat_pre_nz_w[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29656" *) in_dat_nan[28];
  assign _07620_ = dat_pre_nz_w[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29666" *) in_dat_nan[29];
  assign _07621_ = dat_pre_nz_w[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29676" *) in_dat_nan[29];
  assign _07622_ = dat_pre_nz_w[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29686" *) in_dat_nan[30];
  assign _07623_ = dat_pre_nz_w[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29696" *) in_dat_nan[30];
  assign _07624_ = dat_pre_nz_w[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29706" *) in_dat_nan[31];
  assign _07625_ = dat_pre_nz_w[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29716" *) in_dat_nan[31];
  assign _07626_ = dat_pre_nz_w[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29726" *) in_dat_nan[32];
  assign _07627_ = dat_pre_nz_w[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29736" *) in_dat_nan[32];
  assign _07628_ = dat_pre_nz_w[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29746" *) in_dat_nan[33];
  assign _07629_ = dat_pre_nz_w[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29756" *) in_dat_nan[33];
  assign _07630_ = dat_pre_nz_w[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29766" *) in_dat_nan[34];
  assign _07631_ = dat_pre_nz_w[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29776" *) in_dat_nan[34];
  assign _07632_ = dat_pre_nz_w[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29786" *) in_dat_nan[35];
  assign _07633_ = dat_pre_nz_w[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29796" *) in_dat_nan[35];
  assign _07634_ = dat_pre_nz_w[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29806" *) in_dat_nan[36];
  assign _07635_ = dat_pre_nz_w[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29816" *) in_dat_nan[36];
  assign _07636_ = dat_pre_nz_w[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29826" *) in_dat_nan[37];
  assign _07637_ = dat_pre_nz_w[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29836" *) in_dat_nan[37];
  assign _07638_ = dat_pre_nz_w[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29846" *) in_dat_nan[38];
  assign _07639_ = dat_pre_nz_w[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29856" *) in_dat_nan[38];
  assign _07640_ = dat_pre_nz_w[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29866" *) in_dat_nan[39];
  assign _07641_ = dat_pre_nz_w[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29876" *) in_dat_nan[39];
  assign _07642_ = dat_pre_nz_w[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29886" *) in_dat_nan[40];
  assign _07643_ = dat_pre_nz_w[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29896" *) in_dat_nan[40];
  assign _07644_ = dat_pre_nz_w[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29906" *) in_dat_nan[41];
  assign _07645_ = dat_pre_nz_w[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29916" *) in_dat_nan[41];
  assign _07646_ = dat_pre_nz_w[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29926" *) in_dat_nan[42];
  assign _07647_ = dat_pre_nz_w[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29936" *) in_dat_nan[42];
  assign _07648_ = dat_pre_nz_w[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29946" *) in_dat_nan[43];
  assign _07649_ = dat_pre_nz_w[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29956" *) in_dat_nan[43];
  assign _07650_ = dat_pre_nz_w[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29966" *) in_dat_nan[44];
  assign _07651_ = dat_pre_nz_w[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29976" *) in_dat_nan[44];
  assign _07652_ = dat_pre_nz_w[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29986" *) in_dat_nan[45];
  assign _07653_ = dat_pre_nz_w[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29996" *) in_dat_nan[45];
  assign _07654_ = dat_pre_nz_w[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30006" *) in_dat_nan[46];
  assign _07655_ = dat_pre_nz_w[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30016" *) in_dat_nan[46];
  assign _07656_ = dat_pre_nz_w[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30026" *) in_dat_nan[47];
  assign _07657_ = dat_pre_nz_w[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30036" *) in_dat_nan[47];
  assign _07658_ = dat_pre_nz_w[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30046" *) in_dat_nan[48];
  assign _07659_ = dat_pre_nz_w[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30056" *) in_dat_nan[48];
  assign _07660_ = dat_pre_nz_w[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30066" *) in_dat_nan[49];
  assign _07661_ = dat_pre_nz_w[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30076" *) in_dat_nan[49];
  assign _07662_ = dat_pre_nz_w[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30086" *) in_dat_nan[50];
  assign _07663_ = dat_pre_nz_w[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30096" *) in_dat_nan[50];
  assign _07664_ = dat_pre_nz_w[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30106" *) in_dat_nan[51];
  assign _07665_ = dat_pre_nz_w[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30116" *) in_dat_nan[51];
  assign _07666_ = dat_pre_nz_w[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30126" *) in_dat_nan[52];
  assign _07667_ = dat_pre_nz_w[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30136" *) in_dat_nan[52];
  assign _07668_ = dat_pre_nz_w[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30146" *) in_dat_nan[53];
  assign _07669_ = dat_pre_nz_w[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30156" *) in_dat_nan[53];
  assign _07670_ = dat_pre_nz_w[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30166" *) in_dat_nan[54];
  assign _07671_ = dat_pre_nz_w[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30176" *) in_dat_nan[54];
  assign _07672_ = dat_pre_nz_w[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30186" *) in_dat_nan[55];
  assign _07673_ = dat_pre_nz_w[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30196" *) in_dat_nan[55];
  assign _07674_ = dat_pre_nz_w[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30206" *) in_dat_nan[56];
  assign _07675_ = dat_pre_nz_w[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30216" *) in_dat_nan[56];
  assign _07676_ = dat_pre_nz_w[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30226" *) in_dat_nan[57];
  assign _07677_ = dat_pre_nz_w[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30236" *) in_dat_nan[57];
  assign _07678_ = dat_pre_nz_w[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30246" *) in_dat_nan[58];
  assign _07679_ = dat_pre_nz_w[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30256" *) in_dat_nan[58];
  assign _07680_ = dat_pre_nz_w[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30266" *) in_dat_nan[59];
  assign _07681_ = dat_pre_nz_w[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30276" *) in_dat_nan[59];
  assign _07682_ = dat_pre_nz_w[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30286" *) in_dat_nan[60];
  assign _07683_ = dat_pre_nz_w[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30296" *) in_dat_nan[60];
  assign _07684_ = dat_pre_nz_w[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30306" *) in_dat_nan[61];
  assign _07685_ = dat_pre_nz_w[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30316" *) in_dat_nan[61];
  assign _07686_ = dat_pre_nz_w[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30326" *) in_dat_nan[62];
  assign _07687_ = dat_pre_nz_w[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30336" *) in_dat_nan[62];
  assign _07688_ = dat_pre_nz_w[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30346" *) in_dat_nan[63];
  assign _07689_ = dat_pre_nz_w[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30356" *) in_dat_nan[63];
  assign _07690_ = dat_pre_nz[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30674" *) dat_pre_nan[0];
  assign _07691_ = dat_pre_nz[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30684" *) dat_pre_nan[0];
  assign _07692_ = dat_pre_nz[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30694" *) dat_pre_nan[1];
  assign _07693_ = dat_pre_nz[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30704" *) dat_pre_nan[1];
  assign _07694_ = dat_pre_nz[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30714" *) dat_pre_nan[2];
  assign _07695_ = dat_pre_nz[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30724" *) dat_pre_nan[2];
  assign _07696_ = dat_pre_nz[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30734" *) dat_pre_nan[3];
  assign _07697_ = dat_pre_nz[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30744" *) dat_pre_nan[3];
  assign _07698_ = dat_pre_nz[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30754" *) dat_pre_nan[4];
  assign _07699_ = dat_pre_nz[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30764" *) dat_pre_nan[4];
  assign _07700_ = dat_pre_nz[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30774" *) dat_pre_nan[5];
  assign _07701_ = dat_pre_nz[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30784" *) dat_pre_nan[5];
  assign _07702_ = dat_pre_nz[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30794" *) dat_pre_nan[6];
  assign _07703_ = dat_pre_nz[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30804" *) dat_pre_nan[6];
  assign _07704_ = dat_pre_nz[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30814" *) dat_pre_nan[7];
  assign _07705_ = dat_pre_nz[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30824" *) dat_pre_nan[7];
  assign _07706_ = dat_pre_nz[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30834" *) dat_pre_nan[8];
  assign _07707_ = dat_pre_nz[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30844" *) dat_pre_nan[8];
  assign _07708_ = dat_pre_nz[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30854" *) dat_pre_nan[9];
  assign _07709_ = dat_pre_nz[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30864" *) dat_pre_nan[9];
  assign _07710_ = dat_pre_nz[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30874" *) dat_pre_nan[10];
  assign _07711_ = dat_pre_nz[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30884" *) dat_pre_nan[10];
  assign _07712_ = dat_pre_nz[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30894" *) dat_pre_nan[11];
  assign _07713_ = dat_pre_nz[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30904" *) dat_pre_nan[11];
  assign _07714_ = dat_pre_nz[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30914" *) dat_pre_nan[12];
  assign _07715_ = dat_pre_nz[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30924" *) dat_pre_nan[12];
  assign _07716_ = dat_pre_nz[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30934" *) dat_pre_nan[13];
  assign _07717_ = dat_pre_nz[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30944" *) dat_pre_nan[13];
  assign _07718_ = dat_pre_nz[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30954" *) dat_pre_nan[14];
  assign _07719_ = dat_pre_nz[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30964" *) dat_pre_nan[14];
  assign _07720_ = dat_pre_nz[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30974" *) dat_pre_nan[15];
  assign _07721_ = dat_pre_nz[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30984" *) dat_pre_nan[15];
  assign _07722_ = dat_pre_nz[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30994" *) dat_pre_nan[16];
  assign _07723_ = dat_pre_nz[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31004" *) dat_pre_nan[16];
  assign _07724_ = dat_pre_nz[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31014" *) dat_pre_nan[17];
  assign _07725_ = dat_pre_nz[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31024" *) dat_pre_nan[17];
  assign _07726_ = dat_pre_nz[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31034" *) dat_pre_nan[18];
  assign _07727_ = dat_pre_nz[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31044" *) dat_pre_nan[18];
  assign _07728_ = dat_pre_nz[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31054" *) dat_pre_nan[19];
  assign _07729_ = dat_pre_nz[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31064" *) dat_pre_nan[19];
  assign _07730_ = dat_pre_nz[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31074" *) dat_pre_nan[20];
  assign _07731_ = dat_pre_nz[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31084" *) dat_pre_nan[20];
  assign _07732_ = dat_pre_nz[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31094" *) dat_pre_nan[21];
  assign _07733_ = dat_pre_nz[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31104" *) dat_pre_nan[21];
  assign _07734_ = dat_pre_nz[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31114" *) dat_pre_nan[22];
  assign _07735_ = dat_pre_nz[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31124" *) dat_pre_nan[22];
  assign _07736_ = dat_pre_nz[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31134" *) dat_pre_nan[23];
  assign _07737_ = dat_pre_nz[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31144" *) dat_pre_nan[23];
  assign _07738_ = dat_pre_nz[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31154" *) dat_pre_nan[24];
  assign _07739_ = dat_pre_nz[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31164" *) dat_pre_nan[24];
  assign _07740_ = dat_pre_nz[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31174" *) dat_pre_nan[25];
  assign _07741_ = dat_pre_nz[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31184" *) dat_pre_nan[25];
  assign _07742_ = dat_pre_nz[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31194" *) dat_pre_nan[26];
  assign _07743_ = dat_pre_nz[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31204" *) dat_pre_nan[26];
  assign _07744_ = dat_pre_nz[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31214" *) dat_pre_nan[27];
  assign _07745_ = dat_pre_nz[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31224" *) dat_pre_nan[27];
  assign _07746_ = dat_pre_nz[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31234" *) dat_pre_nan[28];
  assign _07747_ = dat_pre_nz[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31244" *) dat_pre_nan[28];
  assign _07748_ = dat_pre_nz[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31254" *) dat_pre_nan[29];
  assign _07749_ = dat_pre_nz[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31264" *) dat_pre_nan[29];
  assign _07750_ = dat_pre_nz[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31274" *) dat_pre_nan[30];
  assign _07751_ = dat_pre_nz[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31284" *) dat_pre_nan[30];
  assign _07752_ = dat_pre_nz[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31294" *) dat_pre_nan[31];
  assign _07753_ = dat_pre_nz[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31304" *) dat_pre_nan[31];
  assign _07754_ = dat_pre_nz[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31314" *) dat_pre_nan[32];
  assign _07755_ = dat_pre_nz[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31324" *) dat_pre_nan[32];
  assign _07756_ = dat_pre_nz[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31334" *) dat_pre_nan[33];
  assign _07757_ = dat_pre_nz[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31344" *) dat_pre_nan[33];
  assign _07758_ = dat_pre_nz[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31354" *) dat_pre_nan[34];
  assign _07759_ = dat_pre_nz[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31364" *) dat_pre_nan[34];
  assign _07760_ = dat_pre_nz[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31374" *) dat_pre_nan[35];
  assign _07761_ = dat_pre_nz[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31384" *) dat_pre_nan[35];
  assign _07762_ = dat_pre_nz[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31394" *) dat_pre_nan[36];
  assign _07763_ = dat_pre_nz[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31404" *) dat_pre_nan[36];
  assign _07764_ = dat_pre_nz[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31414" *) dat_pre_nan[37];
  assign _07765_ = dat_pre_nz[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31424" *) dat_pre_nan[37];
  assign _07766_ = dat_pre_nz[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31434" *) dat_pre_nan[38];
  assign _07767_ = dat_pre_nz[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31444" *) dat_pre_nan[38];
  assign _07768_ = dat_pre_nz[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31454" *) dat_pre_nan[39];
  assign _07769_ = dat_pre_nz[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31464" *) dat_pre_nan[39];
  assign _07770_ = dat_pre_nz[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31474" *) dat_pre_nan[40];
  assign _07771_ = dat_pre_nz[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31484" *) dat_pre_nan[40];
  assign _07772_ = dat_pre_nz[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31494" *) dat_pre_nan[41];
  assign _07773_ = dat_pre_nz[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31504" *) dat_pre_nan[41];
  assign _07774_ = dat_pre_nz[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31514" *) dat_pre_nan[42];
  assign _07775_ = dat_pre_nz[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31524" *) dat_pre_nan[42];
  assign _07776_ = dat_pre_nz[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31534" *) dat_pre_nan[43];
  assign _07777_ = dat_pre_nz[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31544" *) dat_pre_nan[43];
  assign _07778_ = dat_pre_nz[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31554" *) dat_pre_nan[44];
  assign _07779_ = dat_pre_nz[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31564" *) dat_pre_nan[44];
  assign _07780_ = dat_pre_nz[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31574" *) dat_pre_nan[45];
  assign _07781_ = dat_pre_nz[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31584" *) dat_pre_nan[45];
  assign _07782_ = dat_pre_nz[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31594" *) dat_pre_nan[46];
  assign _07783_ = dat_pre_nz[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31604" *) dat_pre_nan[46];
  assign _07784_ = dat_pre_nz[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31614" *) dat_pre_nan[47];
  assign _07785_ = dat_pre_nz[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31624" *) dat_pre_nan[47];
  assign _07786_ = dat_pre_nz[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31634" *) dat_pre_nan[48];
  assign _07787_ = dat_pre_nz[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31644" *) dat_pre_nan[48];
  assign _07788_ = dat_pre_nz[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31654" *) dat_pre_nan[49];
  assign _07789_ = dat_pre_nz[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31664" *) dat_pre_nan[49];
  assign _07790_ = dat_pre_nz[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31674" *) dat_pre_nan[50];
  assign _07791_ = dat_pre_nz[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31684" *) dat_pre_nan[50];
  assign _07792_ = dat_pre_nz[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31694" *) dat_pre_nan[51];
  assign _07793_ = dat_pre_nz[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31704" *) dat_pre_nan[51];
  assign _07794_ = dat_pre_nz[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31714" *) dat_pre_nan[52];
  assign _07795_ = dat_pre_nz[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31724" *) dat_pre_nan[52];
  assign _07796_ = dat_pre_nz[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31734" *) dat_pre_nan[53];
  assign _07797_ = dat_pre_nz[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31744" *) dat_pre_nan[53];
  assign _07798_ = dat_pre_nz[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31754" *) dat_pre_nan[54];
  assign _07799_ = dat_pre_nz[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31764" *) dat_pre_nan[54];
  assign _07800_ = dat_pre_nz[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31774" *) dat_pre_nan[55];
  assign _07801_ = dat_pre_nz[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31784" *) dat_pre_nan[55];
  assign _07802_ = dat_pre_nz[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31794" *) dat_pre_nan[56];
  assign _07803_ = dat_pre_nz[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31804" *) dat_pre_nan[56];
  assign _07804_ = dat_pre_nz[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31814" *) dat_pre_nan[57];
  assign _07805_ = dat_pre_nz[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31824" *) dat_pre_nan[57];
  assign _07806_ = dat_pre_nz[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31834" *) dat_pre_nan[58];
  assign _07807_ = dat_pre_nz[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31844" *) dat_pre_nan[58];
  assign _07808_ = dat_pre_nz[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31854" *) dat_pre_nan[59];
  assign _07809_ = dat_pre_nz[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31864" *) dat_pre_nan[59];
  assign _07810_ = dat_pre_nz[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31874" *) dat_pre_nan[60];
  assign _07811_ = dat_pre_nz[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31884" *) dat_pre_nan[60];
  assign _07812_ = dat_pre_nz[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31894" *) dat_pre_nan[61];
  assign _07813_ = dat_pre_nz[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31904" *) dat_pre_nan[61];
  assign _07814_ = dat_pre_nz[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31914" *) dat_pre_nan[62];
  assign _07815_ = dat_pre_nz[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31924" *) dat_pre_nan[62];
  assign _07816_ = dat_pre_nz[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31934" *) dat_pre_nan[63];
  assign _07817_ = dat_pre_nz[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31944" *) dat_pre_nan[63];
  assign _07818_ = { in_wt_data_fp16_63, in_wt_data_fp16_62, in_wt_data_fp16_61, in_wt_data_fp16_60, in_wt_data_fp16_59, in_wt_data_fp16_58, in_wt_data_fp16_57, in_wt_data_fp16_56, in_wt_data_fp16_55, in_wt_data_fp16_54, in_wt_data_fp16_53, in_wt_data_fp16_52, in_wt_data_fp16_51, in_wt_data_fp16_50, in_wt_data_fp16_49, in_wt_data_fp16_48, in_wt_data_fp16_47, in_wt_data_fp16_46, in_wt_data_fp16_45, in_wt_data_fp16_44, in_wt_data_fp16_43, in_wt_data_fp16_42, in_wt_data_fp16_41, in_wt_data_fp16_40, in_wt_data_fp16_39, in_wt_data_fp16_38, in_wt_data_fp16_37, in_wt_data_fp16_36, in_wt_data_fp16_35, in_wt_data_fp16_34, in_wt_data_fp16_33, in_wt_data_fp16_32, in_wt_data_fp16_31, in_wt_data_fp16_30, in_wt_data_fp16_29, in_wt_data_fp16_28, in_wt_data_fp16_27, in_wt_data_fp16_26, in_wt_data_fp16_25, in_wt_data_fp16_24, in_wt_data_fp16_23, in_wt_data_fp16_22, in_wt_data_fp16_21, in_wt_data_fp16_20, in_wt_data_fp16_19, in_wt_data_fp16_18, in_wt_data_fp16_17, in_wt_data_fp16_16, in_wt_data_fp16_15, in_wt_data_fp16_14, in_wt_data_fp16_13, in_wt_data_fp16_12, in_wt_data_fp16_11, in_wt_data_fp16_10, in_wt_data_fp16_9, in_wt_data_fp16_8, in_wt_data_fp16_7, in_wt_data_fp16_6, in_wt_data_fp16_5, in_wt_data_fp16_4, in_wt_data_fp16_3, in_wt_data_fp16_2, in_wt_data_fp16_1, in_wt_data_fp16_0 } | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3959" *) { in_wt_data_int8_63, in_wt_data_int8_62, in_wt_data_int8_61, in_wt_data_int8_60, in_wt_data_int8_59, in_wt_data_int8_58, in_wt_data_int8_57, in_wt_data_int8_56, in_wt_data_int8_55, in_wt_data_int8_54, in_wt_data_int8_53, in_wt_data_int8_52, in_wt_data_int8_51, in_wt_data_int8_50, in_wt_data_int8_49, in_wt_data_int8_48, in_wt_data_int8_47, in_wt_data_int8_46, in_wt_data_int8_45, in_wt_data_int8_44, in_wt_data_int8_43, in_wt_data_int8_42, in_wt_data_int8_41, in_wt_data_int8_40, in_wt_data_int8_39, in_wt_data_int8_38, in_wt_data_int8_37, in_wt_data_int8_36, in_wt_data_int8_35, in_wt_data_int8_34, in_wt_data_int8_33, in_wt_data_int8_32, in_wt_data_int8_31, in_wt_data_int8_30, in_wt_data_int8_29, in_wt_data_int8_28, in_wt_data_int8_27, in_wt_data_int8_26, in_wt_data_int8_25, in_wt_data_int8_24, in_wt_data_int8_23, in_wt_data_int8_22, in_wt_data_int8_21, in_wt_data_int8_20, in_wt_data_int8_19, in_wt_data_int8_18, in_wt_data_int8_17, in_wt_data_int8_16, in_wt_data_int8_15, in_wt_data_int8_14, in_wt_data_int8_13, in_wt_data_int8_12, in_wt_data_int8_11, in_wt_data_int8_10, in_wt_data_int8_9, in_wt_data_int8_8, in_wt_data_int8_7, in_wt_data_int8_6, in_wt_data_int8_5, in_wt_data_int8_4, in_wt_data_int8_3, in_wt_data_int8_2, in_wt_data_int8_1, in_wt_data_int8_0 };
  assign wt_pre_data_w = _07818_ | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3959" *) { in_wt_data_int16_63, in_wt_data_int16_62, in_wt_data_int16_61, in_wt_data_int16_60, in_wt_data_int16_59, in_wt_data_int16_58, in_wt_data_int16_57, in_wt_data_int16_56, in_wt_data_int16_55, in_wt_data_int16_54, in_wt_data_int16_53, in_wt_data_int16_52, in_wt_data_int16_51, in_wt_data_int16_50, in_wt_data_int16_49, in_wt_data_int16_48, in_wt_data_int16_47, in_wt_data_int16_46, in_wt_data_int16_45, in_wt_data_int16_44, in_wt_data_int16_43, in_wt_data_int16_42, in_wt_data_int16_41, in_wt_data_int16_40, in_wt_data_int16_39, in_wt_data_int16_38, in_wt_data_int16_37, in_wt_data_int16_36, in_wt_data_int16_35, in_wt_data_int16_34, in_wt_data_int16_33, in_wt_data_int16_32, in_wt_data_int16_31, in_wt_data_int16_30, in_wt_data_int16_29, in_wt_data_int16_28, in_wt_data_int16_27, in_wt_data_int16_26, in_wt_data_int16_25, in_wt_data_int16_24, in_wt_data_int16_23, in_wt_data_int16_22, in_wt_data_int16_21, in_wt_data_int16_20, in_wt_data_int16_19, in_wt_data_int16_18, in_wt_data_int16_17, in_wt_data_int16_16, in_wt_data_int16_15, in_wt_data_int16_14, in_wt_data_int16_13, in_wt_data_int16_12, in_wt_data_int16_11, in_wt_data_int16_10, in_wt_data_int16_9, in_wt_data_int16_8, in_wt_data_int16_7, in_wt_data_int16_6, in_wt_data_int16_5, in_wt_data_int16_4, in_wt_data_int16_3, in_wt_data_int16_2, in_wt_data_int16_1, in_wt_data_int16_0 };
  assign _07819_ = wt_pre_nz_w[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4033" *) in_wt_nan[0];
  assign _07820_ = wt_pre_nz_w[1] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4043" *) in_wt_nan[0];
  assign _07821_ = wt_pre_nz_w[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4053" *) in_wt_nan[1];
  assign _07822_ = wt_pre_nz_w[3] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4063" *) in_wt_nan[1];
  assign _07823_ = wt_pre_nz_w[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4073" *) in_wt_nan[2];
  assign _07824_ = wt_pre_nz_w[5] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4083" *) in_wt_nan[2];
  assign _07825_ = wt_pre_nz_w[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4093" *) in_wt_nan[3];
  assign _07826_ = wt_pre_nz_w[7] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4103" *) in_wt_nan[3];
  assign _07827_ = wt_pre_nz_w[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4113" *) in_wt_nan[4];
  assign _07828_ = wt_pre_nz_w[9] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4123" *) in_wt_nan[4];
  assign _07829_ = wt_pre_nz_w[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4133" *) in_wt_nan[5];
  assign _07830_ = wt_pre_nz_w[11] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4143" *) in_wt_nan[5];
  assign _07831_ = wt_pre_nz_w[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4153" *) in_wt_nan[6];
  assign _07832_ = wt_pre_nz_w[13] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4163" *) in_wt_nan[6];
  assign _07833_ = wt_pre_nz_w[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4173" *) in_wt_nan[7];
  assign _07834_ = wt_pre_nz_w[15] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4183" *) in_wt_nan[7];
  assign _07835_ = wt_pre_nz_w[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4193" *) in_wt_nan[8];
  assign _07836_ = wt_pre_nz_w[17] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4203" *) in_wt_nan[8];
  assign _07837_ = wt_pre_nz_w[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4213" *) in_wt_nan[9];
  assign _07838_ = wt_pre_nz_w[19] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4223" *) in_wt_nan[9];
  assign _07839_ = wt_pre_nz_w[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4233" *) in_wt_nan[10];
  assign _07840_ = wt_pre_nz_w[21] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4243" *) in_wt_nan[10];
  assign _07841_ = wt_pre_nz_w[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4253" *) in_wt_nan[11];
  assign _07842_ = wt_pre_nz_w[23] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4263" *) in_wt_nan[11];
  assign _07843_ = wt_pre_nz_w[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4273" *) in_wt_nan[12];
  assign _07844_ = wt_pre_nz_w[25] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4283" *) in_wt_nan[12];
  assign _07845_ = wt_pre_nz_w[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4293" *) in_wt_nan[13];
  assign _07846_ = wt_pre_nz_w[27] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4303" *) in_wt_nan[13];
  assign _07847_ = wt_pre_nz_w[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4313" *) in_wt_nan[14];
  assign _07848_ = wt_pre_nz_w[29] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4323" *) in_wt_nan[14];
  assign _07849_ = wt_pre_nz_w[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4333" *) in_wt_nan[15];
  assign _07850_ = wt_pre_nz_w[31] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4343" *) in_wt_nan[15];
  assign _07851_ = wt_pre_nz_w[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4353" *) in_wt_nan[16];
  assign _07852_ = wt_pre_nz_w[33] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4363" *) in_wt_nan[16];
  assign _07853_ = wt_pre_nz_w[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4373" *) in_wt_nan[17];
  assign _07854_ = wt_pre_nz_w[35] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4383" *) in_wt_nan[17];
  assign _07855_ = wt_pre_nz_w[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4393" *) in_wt_nan[18];
  assign _07856_ = wt_pre_nz_w[37] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4403" *) in_wt_nan[18];
  assign _07857_ = wt_pre_nz_w[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4413" *) in_wt_nan[19];
  assign _07858_ = wt_pre_nz_w[39] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4423" *) in_wt_nan[19];
  assign _07859_ = wt_pre_nz_w[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4433" *) in_wt_nan[20];
  assign _07860_ = wt_pre_nz_w[41] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4443" *) in_wt_nan[20];
  assign _07861_ = wt_pre_nz_w[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4453" *) in_wt_nan[21];
  assign _07862_ = wt_pre_nz_w[43] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4463" *) in_wt_nan[21];
  assign _07863_ = wt_pre_nz_w[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4473" *) in_wt_nan[22];
  assign _07864_ = wt_pre_nz_w[45] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4483" *) in_wt_nan[22];
  assign _07865_ = wt_pre_nz_w[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4493" *) in_wt_nan[23];
  assign _07866_ = wt_pre_nz_w[47] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4503" *) in_wt_nan[23];
  assign _07867_ = wt_pre_nz_w[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4513" *) in_wt_nan[24];
  assign _07868_ = wt_pre_nz_w[49] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4523" *) in_wt_nan[24];
  assign _07869_ = wt_pre_nz_w[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4533" *) in_wt_nan[25];
  assign _07870_ = wt_pre_nz_w[51] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4543" *) in_wt_nan[25];
  assign _07871_ = wt_pre_nz_w[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4553" *) in_wt_nan[26];
  assign _07872_ = wt_pre_nz_w[53] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4563" *) in_wt_nan[26];
  assign _07873_ = wt_pre_nz_w[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4573" *) in_wt_nan[27];
  assign _07874_ = wt_pre_nz_w[55] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4583" *) in_wt_nan[27];
  assign _07875_ = wt_pre_nz_w[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4593" *) in_wt_nan[28];
  assign _07876_ = wt_pre_nz_w[57] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4603" *) in_wt_nan[28];
  assign _07877_ = wt_pre_nz_w[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4613" *) in_wt_nan[29];
  assign _07878_ = wt_pre_nz_w[59] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4623" *) in_wt_nan[29];
  assign _07879_ = wt_pre_nz_w[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4633" *) in_wt_nan[30];
  assign _07880_ = wt_pre_nz_w[61] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4643" *) in_wt_nan[30];
  assign _07881_ = wt_pre_nz_w[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4653" *) in_wt_nan[31];
  assign _07882_ = wt_pre_nz_w[63] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4663" *) in_wt_nan[31];
  assign _07883_ = wt_pre_nz_w[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4673" *) in_wt_nan[32];
  assign _07884_ = wt_pre_nz_w[65] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4683" *) in_wt_nan[32];
  assign _07885_ = wt_pre_nz_w[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4693" *) in_wt_nan[33];
  assign _07886_ = wt_pre_nz_w[67] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4703" *) in_wt_nan[33];
  assign _07887_ = wt_pre_nz_w[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4713" *) in_wt_nan[34];
  assign _07888_ = wt_pre_nz_w[69] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4723" *) in_wt_nan[34];
  assign _07889_ = wt_pre_nz_w[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4733" *) in_wt_nan[35];
  assign _07890_ = wt_pre_nz_w[71] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4743" *) in_wt_nan[35];
  assign _07891_ = wt_pre_nz_w[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4753" *) in_wt_nan[36];
  assign _07892_ = wt_pre_nz_w[73] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4763" *) in_wt_nan[36];
  assign _07893_ = wt_pre_nz_w[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4773" *) in_wt_nan[37];
  assign _07894_ = wt_pre_nz_w[75] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4783" *) in_wt_nan[37];
  assign _07895_ = wt_pre_nz_w[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4793" *) in_wt_nan[38];
  assign _07896_ = wt_pre_nz_w[77] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4803" *) in_wt_nan[38];
  assign _07897_ = wt_pre_nz_w[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4813" *) in_wt_nan[39];
  assign _07898_ = wt_pre_nz_w[79] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4823" *) in_wt_nan[39];
  assign _07899_ = wt_pre_nz_w[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4833" *) in_wt_nan[40];
  assign _07900_ = wt_pre_nz_w[81] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4843" *) in_wt_nan[40];
  assign _07901_ = wt_pre_nz_w[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4853" *) in_wt_nan[41];
  assign _07902_ = wt_pre_nz_w[83] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4863" *) in_wt_nan[41];
  assign _07903_ = wt_pre_nz_w[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4873" *) in_wt_nan[42];
  assign _07904_ = wt_pre_nz_w[85] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4883" *) in_wt_nan[42];
  assign _07905_ = wt_pre_nz_w[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4893" *) in_wt_nan[43];
  assign _07906_ = wt_pre_nz_w[87] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4903" *) in_wt_nan[43];
  assign _07907_ = wt_pre_nz_w[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4913" *) in_wt_nan[44];
  assign _07908_ = wt_pre_nz_w[89] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4923" *) in_wt_nan[44];
  assign _07909_ = wt_pre_nz_w[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4933" *) in_wt_nan[45];
  assign _07910_ = wt_pre_nz_w[91] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4943" *) in_wt_nan[45];
  assign _07911_ = wt_pre_nz_w[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4953" *) in_wt_nan[46];
  assign _07912_ = wt_pre_nz_w[93] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4963" *) in_wt_nan[46];
  assign _07913_ = wt_pre_nz_w[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4973" *) in_wt_nan[47];
  assign _07914_ = wt_pre_nz_w[95] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4983" *) in_wt_nan[47];
  assign _07915_ = wt_pre_nz_w[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4993" *) in_wt_nan[48];
  assign _07916_ = wt_pre_nz_w[97] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5003" *) in_wt_nan[48];
  assign _07917_ = wt_pre_nz_w[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5013" *) in_wt_nan[49];
  assign _07918_ = wt_pre_nz_w[99] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5023" *) in_wt_nan[49];
  assign _07919_ = wt_pre_nz_w[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5033" *) in_wt_nan[50];
  assign _07920_ = wt_pre_nz_w[101] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5043" *) in_wt_nan[50];
  assign _07921_ = wt_pre_nz_w[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5053" *) in_wt_nan[51];
  assign _07922_ = wt_pre_nz_w[103] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5063" *) in_wt_nan[51];
  assign _07923_ = wt_pre_nz_w[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5073" *) in_wt_nan[52];
  assign _07924_ = wt_pre_nz_w[105] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5083" *) in_wt_nan[52];
  assign _07925_ = wt_pre_nz_w[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5093" *) in_wt_nan[53];
  assign _07926_ = wt_pre_nz_w[107] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5103" *) in_wt_nan[53];
  assign _07927_ = wt_pre_nz_w[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5113" *) in_wt_nan[54];
  assign _07928_ = wt_pre_nz_w[109] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5123" *) in_wt_nan[54];
  assign _07929_ = wt_pre_nz_w[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5133" *) in_wt_nan[55];
  assign _07930_ = wt_pre_nz_w[111] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5143" *) in_wt_nan[55];
  assign _07931_ = wt_pre_nz_w[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5153" *) in_wt_nan[56];
  assign _07932_ = wt_pre_nz_w[113] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5163" *) in_wt_nan[56];
  assign _07933_ = wt_pre_nz_w[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5173" *) in_wt_nan[57];
  assign _07934_ = wt_pre_nz_w[115] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5183" *) in_wt_nan[57];
  assign _07935_ = wt_pre_nz_w[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5193" *) in_wt_nan[58];
  assign _07936_ = wt_pre_nz_w[117] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5203" *) in_wt_nan[58];
  assign _07937_ = wt_pre_nz_w[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5213" *) in_wt_nan[59];
  assign _07938_ = wt_pre_nz_w[119] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5223" *) in_wt_nan[59];
  assign _07939_ = wt_pre_nz_w[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5233" *) in_wt_nan[60];
  assign _07940_ = wt_pre_nz_w[121] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5243" *) in_wt_nan[60];
  assign _07941_ = wt_pre_nz_w[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5253" *) in_wt_nan[61];
  assign _07942_ = wt_pre_nz_w[123] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5263" *) in_wt_nan[61];
  assign _07943_ = wt_pre_nz_w[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5273" *) in_wt_nan[62];
  assign _07944_ = wt_pre_nz_w[125] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5283" *) in_wt_nan[62];
  assign _07945_ = wt_pre_nz_w[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5293" *) in_wt_nan[63];
  assign _07946_ = wt_pre_nz_w[127] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5303" *) in_wt_nan[63];
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[1023:1016] <= _00901_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[1015:1008] <= _00900_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[1007:1000] <= _00899_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[999:992] <= _01026_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[991:984] <= _01025_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[983:976] <= _01024_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[975:968] <= _01023_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[967:960] <= _01022_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[959:952] <= _01020_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[951:944] <= _01019_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[943:936] <= _01018_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[935:928] <= _01017_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[927:920] <= _01016_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[919:912] <= _01015_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[911:904] <= _01014_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[903:896] <= _01013_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[895:888] <= _01012_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[887:880] <= _01011_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[879:872] <= _01009_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[871:864] <= _01008_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[863:856] <= _01007_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[855:848] <= _01006_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[847:840] <= _01005_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[839:832] <= _01004_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[831:824] <= _01003_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[823:816] <= _01002_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[815:808] <= _01001_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[807:800] <= _01000_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[799:792] <= _00997_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[791:784] <= _00996_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[783:776] <= _00995_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[775:768] <= _00994_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[767:760] <= _00993_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[759:752] <= _00992_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[751:744] <= _00991_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[743:736] <= _00990_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[735:728] <= _00989_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[727:720] <= _00988_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[719:712] <= _00986_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[711:704] <= _00985_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[703:696] <= _00984_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[695:688] <= _00983_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[687:680] <= _00982_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[679:672] <= _00981_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[671:664] <= _00980_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[663:656] <= _00979_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[655:648] <= _00978_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[647:640] <= _00977_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[639:632] <= _00975_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[631:624] <= _00974_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[623:616] <= _00973_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[615:608] <= _00972_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[607:600] <= _00971_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[599:592] <= _00970_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[591:584] <= _00969_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[583:576] <= _00968_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[575:568] <= _00967_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[567:560] <= _00966_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[559:552] <= _00964_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[551:544] <= _00963_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[543:536] <= _00962_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[535:528] <= _00961_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[527:520] <= _00960_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[519:512] <= _00959_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[511:504] <= _00958_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[503:496] <= _00957_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[495:488] <= _00956_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[487:480] <= _00955_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[479:472] <= _00953_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[471:464] <= _00952_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[463:456] <= _00951_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[455:448] <= _00950_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[447:440] <= _00949_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[439:432] <= _00948_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[431:424] <= _00947_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[423:416] <= _00946_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[415:408] <= _00945_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[407:400] <= _00944_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[399:392] <= _00942_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[391:384] <= _00941_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[383:376] <= _00940_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[375:368] <= _00939_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[367:360] <= _00938_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[359:352] <= _00937_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[351:344] <= _00936_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[343:336] <= _00935_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[335:328] <= _00934_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[327:320] <= _00933_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[319:312] <= _00931_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[311:304] <= _00930_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[303:296] <= _00929_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[295:288] <= _00928_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[287:280] <= _00927_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[279:272] <= _00926_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[271:264] <= _00925_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[263:256] <= _00924_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[255:248] <= _00923_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[247:240] <= _00922_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[239:232] <= _00920_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[231:224] <= _00919_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[223:216] <= _00918_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[215:208] <= _00917_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[207:200] <= _00916_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[199:192] <= _00915_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[191:184] <= _00914_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[183:176] <= _00913_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[175:168] <= _00912_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[167:160] <= _00911_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[159:152] <= _00909_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[151:144] <= _00908_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[143:136] <= _00907_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[135:128] <= _00906_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[127:120] <= _00905_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[119:112] <= _00904_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[111:104] <= _00903_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[103:96] <= _00902_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[95:88] <= _01021_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[87:80] <= _01010_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[79:72] <= _00998_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[71:64] <= _00987_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[63:56] <= _00976_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[55:48] <= _00965_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[47:40] <= _00954_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[39:32] <= _00943_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[31:24] <= _00932_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[23:16] <= _00921_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[15:8] <= _00910_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg7[7:0] <= _00999_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg7 <= _01034_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg7 <= _01042_;
  reg [0:0] \dat_actv_pvld_reg7_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \dat_actv_pvld_reg7_reg[0]  <= 1'b0;
    else
      \dat_actv_pvld_reg7_reg[0]  <= dat_pre_pvld[0];
  assign dat_actv_pvld_reg7[0] = \dat_actv_pvld_reg7_reg[0] ;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[1023:1016] <= _00773_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[1015:1008] <= _00772_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[1007:1000] <= _00771_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[999:992] <= _00898_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[991:984] <= _00897_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[983:976] <= _00896_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[975:968] <= _00895_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[967:960] <= _00894_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[959:952] <= _00892_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[951:944] <= _00891_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[943:936] <= _00890_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[935:928] <= _00889_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[927:920] <= _00888_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[919:912] <= _00887_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[911:904] <= _00886_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[903:896] <= _00885_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[895:888] <= _00884_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[887:880] <= _00883_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[879:872] <= _00881_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[871:864] <= _00880_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[863:856] <= _00879_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[855:848] <= _00878_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[847:840] <= _00877_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[839:832] <= _00876_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[831:824] <= _00875_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[823:816] <= _00874_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[815:808] <= _00873_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[807:800] <= _00872_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[799:792] <= _00869_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[791:784] <= _00868_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[783:776] <= _00867_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[775:768] <= _00866_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[767:760] <= _00865_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[759:752] <= _00864_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[751:744] <= _00863_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[743:736] <= _00862_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[735:728] <= _00861_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[727:720] <= _00860_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[719:712] <= _00858_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[711:704] <= _00857_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[703:696] <= _00856_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[695:688] <= _00855_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[687:680] <= _00854_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[679:672] <= _00853_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[671:664] <= _00852_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[663:656] <= _00851_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[655:648] <= _00850_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[647:640] <= _00849_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[639:632] <= _00847_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[631:624] <= _00846_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[623:616] <= _00845_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[615:608] <= _00844_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[607:600] <= _00843_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[599:592] <= _00842_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[591:584] <= _00841_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[583:576] <= _00840_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[575:568] <= _00839_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[567:560] <= _00838_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[559:552] <= _00836_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[551:544] <= _00835_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[543:536] <= _00834_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[535:528] <= _00833_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[527:520] <= _00832_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[519:512] <= _00831_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[511:504] <= _00830_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[503:496] <= _00829_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[495:488] <= _00828_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[487:480] <= _00827_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[479:472] <= _00825_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[471:464] <= _00824_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[463:456] <= _00823_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[455:448] <= _00822_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[447:440] <= _00821_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[439:432] <= _00820_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[431:424] <= _00819_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[423:416] <= _00818_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[415:408] <= _00817_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[407:400] <= _00816_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[399:392] <= _00814_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[391:384] <= _00813_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[383:376] <= _00812_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[375:368] <= _00811_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[367:360] <= _00810_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[359:352] <= _00809_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[351:344] <= _00808_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[343:336] <= _00807_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[335:328] <= _00806_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[327:320] <= _00805_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[319:312] <= _00803_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[311:304] <= _00802_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[303:296] <= _00801_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[295:288] <= _00800_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[287:280] <= _00799_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[279:272] <= _00798_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[271:264] <= _00797_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[263:256] <= _00796_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[255:248] <= _00795_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[247:240] <= _00794_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[239:232] <= _00792_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[231:224] <= _00791_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[223:216] <= _00790_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[215:208] <= _00789_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[207:200] <= _00788_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[199:192] <= _00787_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[191:184] <= _00786_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[183:176] <= _00785_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[175:168] <= _00784_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[167:160] <= _00783_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[159:152] <= _00781_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[151:144] <= _00780_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[143:136] <= _00779_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[135:128] <= _00778_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[127:120] <= _00777_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[119:112] <= _00776_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[111:104] <= _00775_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[103:96] <= _00774_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[95:88] <= _00893_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[87:80] <= _00882_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[79:72] <= _00870_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[71:64] <= _00859_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[63:56] <= _00848_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[55:48] <= _00837_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[47:40] <= _00826_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[39:32] <= _00815_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[31:24] <= _00804_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[23:16] <= _00793_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[15:8] <= _00782_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg6[7:0] <= _00871_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg6 <= _01033_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg6 <= _01041_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[1023:1016] <= _00645_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[1015:1008] <= _00644_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[1007:1000] <= _00643_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[999:992] <= _00770_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[991:984] <= _00769_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[983:976] <= _00768_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[975:968] <= _00767_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[967:960] <= _00766_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[959:952] <= _00764_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[951:944] <= _00763_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[943:936] <= _00762_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[935:928] <= _00761_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[927:920] <= _00760_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[919:912] <= _00759_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[911:904] <= _00758_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[903:896] <= _00757_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[895:888] <= _00756_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[887:880] <= _00755_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[879:872] <= _00753_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[871:864] <= _00752_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[863:856] <= _00751_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[855:848] <= _00750_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[847:840] <= _00749_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[839:832] <= _00748_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[831:824] <= _00747_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[823:816] <= _00746_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[815:808] <= _00745_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[807:800] <= _00744_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[799:792] <= _00741_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[791:784] <= _00740_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[783:776] <= _00739_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[775:768] <= _00738_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[767:760] <= _00737_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[759:752] <= _00736_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[751:744] <= _00735_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[743:736] <= _00734_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[735:728] <= _00733_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[727:720] <= _00732_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[719:712] <= _00730_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[711:704] <= _00729_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[703:696] <= _00728_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[695:688] <= _00727_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[687:680] <= _00726_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[679:672] <= _00725_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[671:664] <= _00724_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[663:656] <= _00723_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[655:648] <= _00722_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[647:640] <= _00721_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[639:632] <= _00719_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[631:624] <= _00718_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[623:616] <= _00717_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[615:608] <= _00716_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[607:600] <= _00715_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[599:592] <= _00714_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[591:584] <= _00713_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[583:576] <= _00712_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[575:568] <= _00711_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[567:560] <= _00710_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[559:552] <= _00708_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[551:544] <= _00707_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[543:536] <= _00706_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[535:528] <= _00705_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[527:520] <= _00704_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[519:512] <= _00703_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[511:504] <= _00702_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[503:496] <= _00701_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[495:488] <= _00700_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[487:480] <= _00699_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[479:472] <= _00697_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[471:464] <= _00696_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[463:456] <= _00695_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[455:448] <= _00694_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[447:440] <= _00693_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[439:432] <= _00692_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[431:424] <= _00691_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[423:416] <= _00690_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[415:408] <= _00689_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[407:400] <= _00688_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[399:392] <= _00686_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[391:384] <= _00685_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[383:376] <= _00684_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[375:368] <= _00683_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[367:360] <= _00682_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[359:352] <= _00681_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[351:344] <= _00680_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[343:336] <= _00679_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[335:328] <= _00678_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[327:320] <= _00677_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[319:312] <= _00675_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[311:304] <= _00674_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[303:296] <= _00673_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[295:288] <= _00672_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[287:280] <= _00671_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[279:272] <= _00670_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[271:264] <= _00669_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[263:256] <= _00668_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[255:248] <= _00667_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[247:240] <= _00666_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[239:232] <= _00664_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[231:224] <= _00663_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[223:216] <= _00662_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[215:208] <= _00661_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[207:200] <= _00660_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[199:192] <= _00659_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[191:184] <= _00658_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[183:176] <= _00657_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[175:168] <= _00656_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[167:160] <= _00655_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[159:152] <= _00653_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[151:144] <= _00652_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[143:136] <= _00651_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[135:128] <= _00650_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[127:120] <= _00649_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[119:112] <= _00648_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[111:104] <= _00647_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[103:96] <= _00646_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[95:88] <= _00765_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[87:80] <= _00754_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[79:72] <= _00742_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[71:64] <= _00731_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[63:56] <= _00720_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[55:48] <= _00709_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[47:40] <= _00698_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[39:32] <= _00687_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[31:24] <= _00676_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[23:16] <= _00665_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[15:8] <= _00654_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg5[7:0] <= _00743_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg5 <= _01032_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg5 <= _01040_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[1023:1016] <= _00517_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[1015:1008] <= _00516_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[1007:1000] <= _00515_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[999:992] <= _00642_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[991:984] <= _00641_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[983:976] <= _00640_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[975:968] <= _00639_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[967:960] <= _00638_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[959:952] <= _00636_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[951:944] <= _00635_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[943:936] <= _00634_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[935:928] <= _00633_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[927:920] <= _00632_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[919:912] <= _00631_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[911:904] <= _00630_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[903:896] <= _00629_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[895:888] <= _00628_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[887:880] <= _00627_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[879:872] <= _00625_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[871:864] <= _00624_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[863:856] <= _00623_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[855:848] <= _00622_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[847:840] <= _00621_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[839:832] <= _00620_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[831:824] <= _00619_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[823:816] <= _00618_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[815:808] <= _00617_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[807:800] <= _00616_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[799:792] <= _00613_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[791:784] <= _00612_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[783:776] <= _00611_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[775:768] <= _00610_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[767:760] <= _00609_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[759:752] <= _00608_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[751:744] <= _00607_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[743:736] <= _00606_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[735:728] <= _00605_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[727:720] <= _00604_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[719:712] <= _00602_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[711:704] <= _00601_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[703:696] <= _00600_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[695:688] <= _00599_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[687:680] <= _00598_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[679:672] <= _00597_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[671:664] <= _00596_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[663:656] <= _00595_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[655:648] <= _00594_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[647:640] <= _00593_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[639:632] <= _00591_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[631:624] <= _00590_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[623:616] <= _00589_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[615:608] <= _00588_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[607:600] <= _00587_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[599:592] <= _00586_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[591:584] <= _00585_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[583:576] <= _00584_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[575:568] <= _00583_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[567:560] <= _00582_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[559:552] <= _00580_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[551:544] <= _00579_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[543:536] <= _00578_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[535:528] <= _00577_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[527:520] <= _00576_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[519:512] <= _00575_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[511:504] <= _00574_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[503:496] <= _00573_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[495:488] <= _00572_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[487:480] <= _00571_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[479:472] <= _00569_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[471:464] <= _00568_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[463:456] <= _00567_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[455:448] <= _00566_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[447:440] <= _00565_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[439:432] <= _00564_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[431:424] <= _00563_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[423:416] <= _00562_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[415:408] <= _00561_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[407:400] <= _00560_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[399:392] <= _00558_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[391:384] <= _00557_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[383:376] <= _00556_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[375:368] <= _00555_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[367:360] <= _00554_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[359:352] <= _00553_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[351:344] <= _00552_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[343:336] <= _00551_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[335:328] <= _00550_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[327:320] <= _00549_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[319:312] <= _00547_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[311:304] <= _00546_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[303:296] <= _00545_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[295:288] <= _00544_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[287:280] <= _00543_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[279:272] <= _00542_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[271:264] <= _00541_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[263:256] <= _00540_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[255:248] <= _00539_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[247:240] <= _00538_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[239:232] <= _00536_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[231:224] <= _00535_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[223:216] <= _00534_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[215:208] <= _00533_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[207:200] <= _00532_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[199:192] <= _00531_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[191:184] <= _00530_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[183:176] <= _00529_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[175:168] <= _00528_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[167:160] <= _00527_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[159:152] <= _00525_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[151:144] <= _00524_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[143:136] <= _00523_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[135:128] <= _00522_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[127:120] <= _00521_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[119:112] <= _00520_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[111:104] <= _00519_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[103:96] <= _00518_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[95:88] <= _00637_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[87:80] <= _00626_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[79:72] <= _00614_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[71:64] <= _00603_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[63:56] <= _00592_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[55:48] <= _00581_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[47:40] <= _00570_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[39:32] <= _00559_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[31:24] <= _00548_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[23:16] <= _00537_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[15:8] <= _00526_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg4[7:0] <= _00615_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg4 <= _01031_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg4 <= _01039_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[1023:1016] <= _00389_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[1015:1008] <= _00388_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[1007:1000] <= _00387_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[999:992] <= _00514_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[991:984] <= _00513_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[983:976] <= _00512_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[975:968] <= _00511_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[967:960] <= _00510_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[959:952] <= _00508_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[951:944] <= _00507_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[943:936] <= _00506_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[935:928] <= _00505_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[927:920] <= _00504_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[919:912] <= _00503_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[911:904] <= _00502_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[903:896] <= _00501_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[895:888] <= _00500_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[887:880] <= _00499_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[879:872] <= _00497_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[871:864] <= _00496_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[863:856] <= _00495_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[855:848] <= _00494_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[847:840] <= _00493_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[839:832] <= _00492_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[831:824] <= _00491_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[823:816] <= _00490_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[815:808] <= _00489_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[807:800] <= _00488_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[799:792] <= _00485_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[791:784] <= _00484_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[783:776] <= _00483_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[775:768] <= _00482_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[767:760] <= _00481_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[759:752] <= _00480_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[751:744] <= _00479_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[743:736] <= _00478_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[735:728] <= _00477_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[727:720] <= _00476_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[719:712] <= _00474_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[711:704] <= _00473_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[703:696] <= _00472_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[695:688] <= _00471_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[687:680] <= _00470_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[679:672] <= _00469_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[671:664] <= _00468_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[663:656] <= _00467_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[655:648] <= _00466_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[647:640] <= _00465_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[639:632] <= _00463_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[631:624] <= _00462_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[623:616] <= _00461_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[615:608] <= _00460_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[607:600] <= _00459_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[599:592] <= _00458_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[591:584] <= _00457_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[583:576] <= _00456_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[575:568] <= _00455_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[567:560] <= _00454_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[559:552] <= _00452_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[551:544] <= _00451_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[543:536] <= _00450_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[535:528] <= _00449_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[527:520] <= _00448_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[519:512] <= _00447_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[511:504] <= _00446_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[503:496] <= _00445_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[495:488] <= _00444_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[487:480] <= _00443_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[479:472] <= _00441_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[471:464] <= _00440_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[463:456] <= _00439_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[455:448] <= _00438_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[447:440] <= _00437_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[439:432] <= _00436_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[431:424] <= _00435_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[423:416] <= _00434_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[415:408] <= _00433_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[407:400] <= _00432_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[399:392] <= _00430_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[391:384] <= _00429_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[383:376] <= _00428_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[375:368] <= _00427_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[367:360] <= _00426_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[359:352] <= _00425_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[351:344] <= _00424_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[343:336] <= _00423_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[335:328] <= _00422_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[327:320] <= _00421_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[319:312] <= _00419_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[311:304] <= _00418_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[303:296] <= _00417_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[295:288] <= _00416_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[287:280] <= _00415_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[279:272] <= _00414_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[271:264] <= _00413_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[263:256] <= _00412_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[255:248] <= _00411_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[247:240] <= _00410_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[239:232] <= _00408_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[231:224] <= _00407_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[223:216] <= _00406_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[215:208] <= _00405_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[207:200] <= _00404_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[199:192] <= _00403_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[191:184] <= _00402_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[183:176] <= _00401_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[175:168] <= _00400_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[167:160] <= _00399_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[159:152] <= _00397_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[151:144] <= _00396_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[143:136] <= _00395_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[135:128] <= _00394_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[127:120] <= _00393_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[119:112] <= _00392_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[111:104] <= _00391_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[103:96] <= _00390_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[95:88] <= _00509_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[87:80] <= _00498_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[79:72] <= _00486_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[71:64] <= _00475_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[63:56] <= _00464_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[55:48] <= _00453_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[47:40] <= _00442_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[39:32] <= _00431_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[31:24] <= _00420_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[23:16] <= _00409_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[15:8] <= _00398_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg3[7:0] <= _00487_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg3 <= _01030_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg3 <= _01038_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[1023:1016] <= _00261_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[1015:1008] <= _00260_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[1007:1000] <= _00259_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[999:992] <= _00386_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[991:984] <= _00385_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[983:976] <= _00384_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[975:968] <= _00383_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[967:960] <= _00382_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[959:952] <= _00380_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[951:944] <= _00379_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[943:936] <= _00378_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[935:928] <= _00377_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[927:920] <= _00376_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[919:912] <= _00375_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[911:904] <= _00374_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[903:896] <= _00373_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[895:888] <= _00372_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[887:880] <= _00371_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[879:872] <= _00369_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[871:864] <= _00368_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[863:856] <= _00367_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[855:848] <= _00366_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[847:840] <= _00365_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[839:832] <= _00364_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[831:824] <= _00363_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[823:816] <= _00362_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[815:808] <= _00361_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[807:800] <= _00360_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[799:792] <= _00357_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[791:784] <= _00356_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[783:776] <= _00355_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[775:768] <= _00354_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[767:760] <= _00353_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[759:752] <= _00352_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[751:744] <= _00351_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[743:736] <= _00350_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[735:728] <= _00349_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[727:720] <= _00348_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[719:712] <= _00346_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[711:704] <= _00345_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[703:696] <= _00344_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[695:688] <= _00343_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[687:680] <= _00342_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[679:672] <= _00341_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[671:664] <= _00340_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[663:656] <= _00339_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[655:648] <= _00338_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[647:640] <= _00337_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[639:632] <= _00335_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[631:624] <= _00334_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[623:616] <= _00333_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[615:608] <= _00332_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[607:600] <= _00331_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[599:592] <= _00330_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[591:584] <= _00329_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[583:576] <= _00328_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[575:568] <= _00327_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[567:560] <= _00326_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[559:552] <= _00324_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[551:544] <= _00323_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[543:536] <= _00322_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[535:528] <= _00321_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[527:520] <= _00320_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[519:512] <= _00319_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[511:504] <= _00318_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[503:496] <= _00317_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[495:488] <= _00316_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[487:480] <= _00315_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[479:472] <= _00313_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[471:464] <= _00312_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[463:456] <= _00311_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[455:448] <= _00310_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[447:440] <= _00309_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[439:432] <= _00308_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[431:424] <= _00307_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[423:416] <= _00306_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[415:408] <= _00305_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[407:400] <= _00304_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[399:392] <= _00302_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[391:384] <= _00301_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[383:376] <= _00300_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[375:368] <= _00299_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[367:360] <= _00298_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[359:352] <= _00297_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[351:344] <= _00296_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[343:336] <= _00295_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[335:328] <= _00294_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[327:320] <= _00293_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[319:312] <= _00291_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[311:304] <= _00290_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[303:296] <= _00289_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[295:288] <= _00288_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[287:280] <= _00287_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[279:272] <= _00286_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[271:264] <= _00285_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[263:256] <= _00284_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[255:248] <= _00283_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[247:240] <= _00282_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[239:232] <= _00280_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[231:224] <= _00279_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[223:216] <= _00278_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[215:208] <= _00277_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[207:200] <= _00276_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[199:192] <= _00275_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[191:184] <= _00274_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[183:176] <= _00273_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[175:168] <= _00272_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[167:160] <= _00271_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[159:152] <= _00269_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[151:144] <= _00268_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[143:136] <= _00267_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[135:128] <= _00266_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[127:120] <= _00265_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[119:112] <= _00264_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[111:104] <= _00263_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[103:96] <= _00262_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[95:88] <= _00381_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[87:80] <= _00370_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[79:72] <= _00358_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[71:64] <= _00347_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[63:56] <= _00336_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[55:48] <= _00325_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[47:40] <= _00314_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[39:32] <= _00303_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[31:24] <= _00292_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[23:16] <= _00281_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[15:8] <= _00270_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg2[7:0] <= _00359_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg2 <= _01029_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg2 <= _01037_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[1023:1016] <= _00133_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[1015:1008] <= _00132_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[1007:1000] <= _00131_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[999:992] <= _00258_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[991:984] <= _00257_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[983:976] <= _00256_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[975:968] <= _00255_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[967:960] <= _00254_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[959:952] <= _00252_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[951:944] <= _00251_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[943:936] <= _00250_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[935:928] <= _00249_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[927:920] <= _00248_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[919:912] <= _00247_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[911:904] <= _00246_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[903:896] <= _00245_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[895:888] <= _00244_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[887:880] <= _00243_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[879:872] <= _00241_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[871:864] <= _00240_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[863:856] <= _00239_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[855:848] <= _00238_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[847:840] <= _00237_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[839:832] <= _00236_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[831:824] <= _00235_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[823:816] <= _00234_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[815:808] <= _00233_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[807:800] <= _00232_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[799:792] <= _00229_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[791:784] <= _00228_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[783:776] <= _00227_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[775:768] <= _00226_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[767:760] <= _00225_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[759:752] <= _00224_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[751:744] <= _00223_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[743:736] <= _00222_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[735:728] <= _00221_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[727:720] <= _00220_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[719:712] <= _00218_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[711:704] <= _00217_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[703:696] <= _00216_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[695:688] <= _00215_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[687:680] <= _00214_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[679:672] <= _00213_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[671:664] <= _00212_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[663:656] <= _00211_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[655:648] <= _00210_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[647:640] <= _00209_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[639:632] <= _00207_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[631:624] <= _00206_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[623:616] <= _00205_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[615:608] <= _00204_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[607:600] <= _00203_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[599:592] <= _00202_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[591:584] <= _00201_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[583:576] <= _00200_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[575:568] <= _00199_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[567:560] <= _00198_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[559:552] <= _00196_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[551:544] <= _00195_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[543:536] <= _00194_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[535:528] <= _00193_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[527:520] <= _00192_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[519:512] <= _00191_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[511:504] <= _00190_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[503:496] <= _00189_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[495:488] <= _00188_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[487:480] <= _00187_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[479:472] <= _00185_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[471:464] <= _00184_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[463:456] <= _00183_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[455:448] <= _00182_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[447:440] <= _00181_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[439:432] <= _00180_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[431:424] <= _00179_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[423:416] <= _00178_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[415:408] <= _00177_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[407:400] <= _00176_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[399:392] <= _00174_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[391:384] <= _00173_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[383:376] <= _00172_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[375:368] <= _00171_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[367:360] <= _00170_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[359:352] <= _00169_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[351:344] <= _00168_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[343:336] <= _00167_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[335:328] <= _00166_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[327:320] <= _00165_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[319:312] <= _00163_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[311:304] <= _00162_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[303:296] <= _00161_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[295:288] <= _00160_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[287:280] <= _00159_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[279:272] <= _00158_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[271:264] <= _00157_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[263:256] <= _00156_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[255:248] <= _00155_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[247:240] <= _00154_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[239:232] <= _00152_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[231:224] <= _00151_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[223:216] <= _00150_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[215:208] <= _00149_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[207:200] <= _00148_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[199:192] <= _00147_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[191:184] <= _00146_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[183:176] <= _00145_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[175:168] <= _00144_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[167:160] <= _00143_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[159:152] <= _00141_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[151:144] <= _00140_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[143:136] <= _00139_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[135:128] <= _00138_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[127:120] <= _00137_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[119:112] <= _00136_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[111:104] <= _00135_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[103:96] <= _00134_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[95:88] <= _00253_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[87:80] <= _00242_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[79:72] <= _00230_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[71:64] <= _00219_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[63:56] <= _00208_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[55:48] <= _00197_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[47:40] <= _00186_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[39:32] <= _00175_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[31:24] <= _00164_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[23:16] <= _00153_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[15:8] <= _00142_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg1[7:0] <= _00231_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg1 <= _01028_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg1 <= _01036_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[1023:1016] <= _00005_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[1015:1008] <= _00004_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[1007:1000] <= _00003_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[999:992] <= _00130_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[991:984] <= _00129_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[983:976] <= _00128_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[975:968] <= _00127_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[967:960] <= _00126_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[959:952] <= _00124_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[951:944] <= _00123_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[943:936] <= _00122_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[935:928] <= _00121_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[927:920] <= _00120_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[919:912] <= _00119_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[911:904] <= _00118_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[903:896] <= _00117_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[895:888] <= _00116_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[887:880] <= _00115_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[879:872] <= _00113_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[871:864] <= _00112_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[863:856] <= _00111_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[855:848] <= _00110_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[847:840] <= _00109_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[839:832] <= _00108_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[831:824] <= _00107_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[823:816] <= _00106_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[815:808] <= _00105_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[807:800] <= _00104_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[799:792] <= _00101_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[791:784] <= _00100_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[783:776] <= _00099_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[775:768] <= _00098_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[767:760] <= _00097_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[759:752] <= _00096_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[751:744] <= _00095_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[743:736] <= _00094_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[735:728] <= _00093_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[727:720] <= _00092_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[719:712] <= _00090_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[711:704] <= _00089_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[703:696] <= _00088_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[695:688] <= _00087_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[687:680] <= _00086_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[679:672] <= _00085_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[671:664] <= _00084_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[663:656] <= _00083_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[655:648] <= _00082_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[647:640] <= _00081_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[639:632] <= _00079_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[631:624] <= _00078_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[623:616] <= _00077_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[615:608] <= _00076_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[607:600] <= _00075_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[599:592] <= _00074_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[591:584] <= _00073_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[583:576] <= _00072_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[575:568] <= _00071_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[567:560] <= _00070_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[559:552] <= _00068_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[551:544] <= _00067_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[543:536] <= _00066_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[535:528] <= _00065_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[527:520] <= _00064_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[519:512] <= _00063_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[511:504] <= _00062_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[503:496] <= _00061_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[495:488] <= _00060_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[487:480] <= _00059_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[479:472] <= _00057_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[471:464] <= _00056_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[463:456] <= _00055_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[455:448] <= _00054_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[447:440] <= _00053_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[439:432] <= _00052_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[431:424] <= _00051_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[423:416] <= _00050_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[415:408] <= _00049_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[407:400] <= _00048_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[399:392] <= _00046_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[391:384] <= _00045_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[383:376] <= _00044_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[375:368] <= _00043_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[367:360] <= _00042_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[359:352] <= _00041_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[351:344] <= _00040_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[343:336] <= _00039_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[335:328] <= _00038_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[327:320] <= _00037_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[319:312] <= _00035_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[311:304] <= _00034_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[303:296] <= _00033_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[295:288] <= _00032_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[287:280] <= _00031_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[279:272] <= _00030_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[271:264] <= _00029_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[263:256] <= _00028_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[255:248] <= _00027_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[247:240] <= _00026_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[239:232] <= _00024_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[231:224] <= _00023_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[223:216] <= _00022_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[215:208] <= _00021_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[207:200] <= _00020_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[199:192] <= _00019_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[191:184] <= _00018_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[183:176] <= _00017_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[175:168] <= _00016_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[167:160] <= _00015_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[159:152] <= _00013_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[151:144] <= _00012_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[143:136] <= _00011_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[135:128] <= _00010_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[127:120] <= _00009_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[119:112] <= _00008_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[111:104] <= _00007_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[103:96] <= _00006_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[95:88] <= _00125_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[87:80] <= _00114_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[79:72] <= _00102_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[71:64] <= _00091_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[63:56] <= _00080_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[55:48] <= _00069_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[47:40] <= _00058_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[39:32] <= _00047_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[31:24] <= _00036_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[23:16] <= _00025_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[15:8] <= _00014_;
  always @(posedge nvdla_core_clk)
      dat_actv_data_reg0[7:0] <= _00103_;
  always @(posedge nvdla_core_clk)
      dat_actv_nan_reg0 <= _01027_;
  always @(posedge nvdla_core_clk)
      dat_actv_nz_reg0 <= _01035_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg7 <= _01178_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask7 <= _01186_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg6 <= _01177_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask6 <= _01185_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg5 <= _01176_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask5 <= _01184_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg4 <= _01175_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask4 <= _01183_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg3 <= _01174_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask3 <= _01182_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg2 <= _01173_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask2 <= _01181_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg1 <= _01172_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask1 <= _01180_;
  always @(posedge nvdla_core_clk)
      dat_pre_exp_reg0 <= _01171_;
  always @(posedge nvdla_core_clk)
      dat_pre_mask0 <= _01179_;
  reg [0:0] \dat_pre_stripe_end_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \dat_pre_stripe_end_reg[0]  <= 1'b0;
    else
      \dat_pre_stripe_end_reg[0]  <= _01189_[8];
  assign dat_pre_stripe_end[0] = \dat_pre_stripe_end_reg[0] ;
  reg [0:0] \dat_pre_stripe_st_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \dat_pre_stripe_st_reg[0]  <= 1'b0;
    else
      \dat_pre_stripe_st_reg[0]  <= _01190_[15];
  assign dat_pre_stripe_st[0] = \dat_pre_stripe_st_reg[0] ;
  always @(posedge nvdla_core_clk)
      dat_pre_data[1023:1016] <= _01045_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[1015:1008] <= _01044_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[1007:1000] <= _01043_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[999:992] <= _01170_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[991:984] <= _01169_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[983:976] <= _01168_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[975:968] <= _01167_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[967:960] <= _01166_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[959:952] <= _01164_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[951:944] <= _01163_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[943:936] <= _01162_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[935:928] <= _01161_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[927:920] <= _01160_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[919:912] <= _01159_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[911:904] <= _01158_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[903:896] <= _01157_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[895:888] <= _01156_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[887:880] <= _01155_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[879:872] <= _01153_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[871:864] <= _01152_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[863:856] <= _01151_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[855:848] <= _01150_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[847:840] <= _01149_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[839:832] <= _01148_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[831:824] <= _01147_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[823:816] <= _01146_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[815:808] <= _01145_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[807:800] <= _01144_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[799:792] <= _01141_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[791:784] <= _01140_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[783:776] <= _01139_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[775:768] <= _01138_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[767:760] <= _01137_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[759:752] <= _01136_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[751:744] <= _01135_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[743:736] <= _01134_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[735:728] <= _01133_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[727:720] <= _01132_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[719:712] <= _01130_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[711:704] <= _01129_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[703:696] <= _01128_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[695:688] <= _01127_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[687:680] <= _01126_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[679:672] <= _01125_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[671:664] <= _01124_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[663:656] <= _01123_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[655:648] <= _01122_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[647:640] <= _01121_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[639:632] <= _01119_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[631:624] <= _01118_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[623:616] <= _01117_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[615:608] <= _01116_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[607:600] <= _01115_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[599:592] <= _01114_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[591:584] <= _01113_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[583:576] <= _01112_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[575:568] <= _01111_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[567:560] <= _01110_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[559:552] <= _01108_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[551:544] <= _01107_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[543:536] <= _01106_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[535:528] <= _01105_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[527:520] <= _01104_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[519:512] <= _01103_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[511:504] <= _01102_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[503:496] <= _01101_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[495:488] <= _01100_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[487:480] <= _01099_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[479:472] <= _01097_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[471:464] <= _01096_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[463:456] <= _01095_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[455:448] <= _01094_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[447:440] <= _01093_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[439:432] <= _01092_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[431:424] <= _01091_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[423:416] <= _01090_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[415:408] <= _01089_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[407:400] <= _01088_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[399:392] <= _01086_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[391:384] <= _01085_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[383:376] <= _01084_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[375:368] <= _01083_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[367:360] <= _01082_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[359:352] <= _01081_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[351:344] <= _01080_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[343:336] <= _01079_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[335:328] <= _01078_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[327:320] <= _01077_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[319:312] <= _01075_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[311:304] <= _01074_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[303:296] <= _01073_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[295:288] <= _01072_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[287:280] <= _01071_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[279:272] <= _01070_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[271:264] <= _01069_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[263:256] <= _01068_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[255:248] <= _01067_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[247:240] <= _01066_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[239:232] <= _01064_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[231:224] <= _01063_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[223:216] <= _01062_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[215:208] <= _01061_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[207:200] <= _01060_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[199:192] <= _01059_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[191:184] <= _01058_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[183:176] <= _01057_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[175:168] <= _01056_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[167:160] <= _01055_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[159:152] <= _01053_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[151:144] <= _01052_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[143:136] <= _01051_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[135:128] <= _01050_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[127:120] <= _01049_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[119:112] <= _01048_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[111:104] <= _01047_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[103:96] <= _01046_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[95:88] <= _01165_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[87:80] <= _01154_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[79:72] <= _01142_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[71:64] <= _01131_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[63:56] <= _01120_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[55:48] <= _01109_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[47:40] <= _01098_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[39:32] <= _01087_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[31:24] <= _01076_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[23:16] <= _01065_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[15:8] <= _01054_;
  always @(posedge nvdla_core_clk)
      dat_pre_data[7:0] <= _01143_;
  always @(posedge nvdla_core_clk)
      dat_pre_nan <= _01187_;
  always @(posedge nvdla_core_clk)
      dat_pre_nz <= _01188_;
  reg [0:0] \dat_pre_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \dat_pre_pvld_reg[0]  <= 1'b0;
    else
      \dat_pre_pvld_reg[0]  <= in_dat_pvld;
  assign dat_pre_pvld[0] = \dat_pre_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_actv_stripe_end <= 1'b0;
    else
      dat_actv_stripe_end <= dat_pre_stripe_end[0];
  always @(posedge nvdla_core_clk)
      wt7_actv_data[1023:1016] <= _03027_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[1015:1008] <= _03026_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[1007:1000] <= _03025_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[999:992] <= _03152_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[991:984] <= _03151_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[983:976] <= _03150_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[975:968] <= _03149_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[967:960] <= _03148_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[959:952] <= _03146_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[951:944] <= _03145_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[943:936] <= _03144_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[935:928] <= _03143_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[927:920] <= _03142_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[919:912] <= _03141_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[911:904] <= _03140_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[903:896] <= _03139_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[895:888] <= _03138_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[887:880] <= _03137_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[879:872] <= _03135_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[871:864] <= _03134_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[863:856] <= _03133_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[855:848] <= _03132_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[847:840] <= _03131_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[839:832] <= _03130_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[831:824] <= _03129_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[823:816] <= _03128_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[815:808] <= _03127_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[807:800] <= _03126_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[799:792] <= _03123_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[791:784] <= _03122_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[783:776] <= _03121_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[775:768] <= _03120_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[767:760] <= _03119_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[759:752] <= _03118_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[751:744] <= _03117_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[743:736] <= _03116_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[735:728] <= _03115_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[727:720] <= _03114_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[719:712] <= _03112_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[711:704] <= _03111_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[703:696] <= _03110_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[695:688] <= _03109_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[687:680] <= _03108_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[679:672] <= _03107_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[671:664] <= _03106_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[663:656] <= _03105_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[655:648] <= _03104_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[647:640] <= _03103_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[639:632] <= _03101_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[631:624] <= _03100_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[623:616] <= _03099_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[615:608] <= _03098_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[607:600] <= _03097_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[599:592] <= _03096_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[591:584] <= _03095_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[583:576] <= _03094_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[575:568] <= _03093_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[567:560] <= _03092_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[559:552] <= _03090_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[551:544] <= _03089_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[543:536] <= _03088_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[535:528] <= _03087_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[527:520] <= _03086_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[519:512] <= _03085_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[511:504] <= _03084_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[503:496] <= _03083_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[495:488] <= _03082_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[487:480] <= _03081_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[479:472] <= _03079_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[471:464] <= _03078_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[463:456] <= _03077_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[455:448] <= _03076_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[447:440] <= _03075_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[439:432] <= _03074_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[431:424] <= _03073_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[423:416] <= _03072_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[415:408] <= _03071_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[407:400] <= _03070_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[399:392] <= _03068_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[391:384] <= _03067_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[383:376] <= _03066_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[375:368] <= _03065_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[367:360] <= _03064_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[359:352] <= _03063_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[351:344] <= _03062_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[343:336] <= _03061_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[335:328] <= _03060_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[327:320] <= _03059_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[319:312] <= _03057_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[311:304] <= _03056_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[303:296] <= _03055_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[295:288] <= _03054_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[287:280] <= _03053_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[279:272] <= _03052_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[271:264] <= _03051_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[263:256] <= _03050_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[255:248] <= _03049_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[247:240] <= _03048_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[239:232] <= _03046_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[231:224] <= _03045_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[223:216] <= _03044_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[215:208] <= _03043_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[207:200] <= _03042_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[199:192] <= _03041_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[191:184] <= _03040_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[183:176] <= _03039_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[175:168] <= _03038_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[167:160] <= _03037_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[159:152] <= _03035_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[151:144] <= _03034_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[143:136] <= _03033_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[135:128] <= _03032_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[127:120] <= _03031_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[119:112] <= _03030_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[111:104] <= _03029_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[103:96] <= _03028_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[95:88] <= _03147_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[87:80] <= _03136_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[79:72] <= _03124_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[71:64] <= _03113_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[63:56] <= _03102_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[55:48] <= _03091_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[47:40] <= _03080_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[39:32] <= _03069_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[31:24] <= _03058_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[23:16] <= _03047_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[15:8] <= _03036_;
  always @(posedge nvdla_core_clk)
      wt7_actv_data[7:0] <= _03125_;
  always @(posedge nvdla_core_clk)
      wt7_actv_nan <= _03153_;
  always @(posedge nvdla_core_clk)
      wt7_actv_nz <= _03154_;
  reg [0:0] \wt7_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt7_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt7_actv_pvld_reg[0]  <= wt7_actv_pvld_w;
  assign wt7_actv_pvld[0] = \wt7_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[1023:1016] <= _02765_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[1015:1008] <= _02764_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[1007:1000] <= _02763_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[999:992] <= _02890_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[991:984] <= _02889_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[983:976] <= _02888_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[975:968] <= _02887_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[967:960] <= _02886_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[959:952] <= _02884_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[951:944] <= _02883_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[943:936] <= _02882_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[935:928] <= _02881_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[927:920] <= _02880_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[919:912] <= _02879_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[911:904] <= _02878_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[903:896] <= _02877_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[895:888] <= _02876_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[887:880] <= _02875_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[879:872] <= _02873_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[871:864] <= _02872_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[863:856] <= _02871_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[855:848] <= _02870_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[847:840] <= _02869_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[839:832] <= _02868_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[831:824] <= _02867_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[823:816] <= _02866_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[815:808] <= _02865_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[807:800] <= _02864_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[799:792] <= _02861_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[791:784] <= _02860_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[783:776] <= _02859_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[775:768] <= _02858_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[767:760] <= _02857_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[759:752] <= _02856_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[751:744] <= _02855_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[743:736] <= _02854_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[735:728] <= _02853_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[727:720] <= _02852_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[719:712] <= _02850_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[711:704] <= _02849_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[703:696] <= _02848_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[695:688] <= _02847_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[687:680] <= _02846_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[679:672] <= _02845_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[671:664] <= _02844_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[663:656] <= _02843_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[655:648] <= _02842_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[647:640] <= _02841_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[639:632] <= _02839_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[631:624] <= _02838_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[623:616] <= _02837_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[615:608] <= _02836_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[607:600] <= _02835_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[599:592] <= _02834_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[591:584] <= _02833_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[583:576] <= _02832_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[575:568] <= _02831_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[567:560] <= _02830_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[559:552] <= _02828_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[551:544] <= _02827_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[543:536] <= _02826_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[535:528] <= _02825_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[527:520] <= _02824_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[519:512] <= _02823_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[511:504] <= _02822_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[503:496] <= _02821_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[495:488] <= _02820_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[487:480] <= _02819_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[479:472] <= _02817_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[471:464] <= _02816_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[463:456] <= _02815_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[455:448] <= _02814_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[447:440] <= _02813_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[439:432] <= _02812_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[431:424] <= _02811_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[423:416] <= _02810_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[415:408] <= _02809_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[407:400] <= _02808_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[399:392] <= _02806_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[391:384] <= _02805_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[383:376] <= _02804_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[375:368] <= _02803_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[367:360] <= _02802_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[359:352] <= _02801_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[351:344] <= _02800_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[343:336] <= _02799_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[335:328] <= _02798_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[327:320] <= _02797_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[319:312] <= _02795_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[311:304] <= _02794_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[303:296] <= _02793_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[295:288] <= _02792_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[287:280] <= _02791_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[279:272] <= _02790_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[271:264] <= _02789_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[263:256] <= _02788_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[255:248] <= _02787_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[247:240] <= _02786_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[239:232] <= _02784_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[231:224] <= _02783_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[223:216] <= _02782_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[215:208] <= _02781_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[207:200] <= _02780_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[199:192] <= _02779_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[191:184] <= _02778_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[183:176] <= _02777_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[175:168] <= _02776_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[167:160] <= _02775_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[159:152] <= _02773_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[151:144] <= _02772_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[143:136] <= _02771_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[135:128] <= _02770_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[127:120] <= _02769_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[119:112] <= _02768_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[111:104] <= _02767_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[103:96] <= _02766_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[95:88] <= _02885_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[87:80] <= _02874_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[79:72] <= _02862_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[71:64] <= _02851_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[63:56] <= _02840_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[55:48] <= _02829_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[47:40] <= _02818_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[39:32] <= _02807_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[31:24] <= _02796_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[23:16] <= _02785_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[15:8] <= _02774_;
  always @(posedge nvdla_core_clk)
      wt6_actv_data[7:0] <= _02863_;
  always @(posedge nvdla_core_clk)
      wt6_actv_nan <= _02891_;
  always @(posedge nvdla_core_clk)
      wt6_actv_nz <= _02892_;
  reg [0:0] \wt6_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt6_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt6_actv_pvld_reg[0]  <= wt6_actv_pvld_w;
  assign wt6_actv_pvld[0] = \wt6_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[1023:1016] <= _02503_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[1015:1008] <= _02502_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[1007:1000] <= _02501_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[999:992] <= _02628_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[991:984] <= _02627_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[983:976] <= _02626_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[975:968] <= _02625_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[967:960] <= _02624_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[959:952] <= _02622_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[951:944] <= _02621_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[943:936] <= _02620_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[935:928] <= _02619_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[927:920] <= _02618_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[919:912] <= _02617_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[911:904] <= _02616_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[903:896] <= _02615_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[895:888] <= _02614_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[887:880] <= _02613_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[879:872] <= _02611_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[871:864] <= _02610_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[863:856] <= _02609_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[855:848] <= _02608_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[847:840] <= _02607_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[839:832] <= _02606_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[831:824] <= _02605_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[823:816] <= _02604_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[815:808] <= _02603_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[807:800] <= _02602_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[799:792] <= _02599_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[791:784] <= _02598_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[783:776] <= _02597_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[775:768] <= _02596_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[767:760] <= _02595_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[759:752] <= _02594_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[751:744] <= _02593_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[743:736] <= _02592_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[735:728] <= _02591_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[727:720] <= _02590_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[719:712] <= _02588_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[711:704] <= _02587_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[703:696] <= _02586_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[695:688] <= _02585_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[687:680] <= _02584_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[679:672] <= _02583_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[671:664] <= _02582_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[663:656] <= _02581_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[655:648] <= _02580_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[647:640] <= _02579_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[639:632] <= _02577_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[631:624] <= _02576_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[623:616] <= _02575_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[615:608] <= _02574_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[607:600] <= _02573_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[599:592] <= _02572_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[591:584] <= _02571_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[583:576] <= _02570_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[575:568] <= _02569_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[567:560] <= _02568_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[559:552] <= _02566_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[551:544] <= _02565_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[543:536] <= _02564_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[535:528] <= _02563_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[527:520] <= _02562_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[519:512] <= _02561_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[511:504] <= _02560_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[503:496] <= _02559_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[495:488] <= _02558_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[487:480] <= _02557_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[479:472] <= _02555_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[471:464] <= _02554_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[463:456] <= _02553_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[455:448] <= _02552_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[447:440] <= _02551_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[439:432] <= _02550_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[431:424] <= _02549_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[423:416] <= _02548_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[415:408] <= _02547_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[407:400] <= _02546_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[399:392] <= _02544_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[391:384] <= _02543_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[383:376] <= _02542_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[375:368] <= _02541_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[367:360] <= _02540_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[359:352] <= _02539_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[351:344] <= _02538_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[343:336] <= _02537_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[335:328] <= _02536_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[327:320] <= _02535_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[319:312] <= _02533_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[311:304] <= _02532_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[303:296] <= _02531_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[295:288] <= _02530_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[287:280] <= _02529_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[279:272] <= _02528_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[271:264] <= _02527_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[263:256] <= _02526_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[255:248] <= _02525_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[247:240] <= _02524_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[239:232] <= _02522_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[231:224] <= _02521_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[223:216] <= _02520_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[215:208] <= _02519_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[207:200] <= _02518_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[199:192] <= _02517_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[191:184] <= _02516_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[183:176] <= _02515_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[175:168] <= _02514_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[167:160] <= _02513_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[159:152] <= _02511_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[151:144] <= _02510_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[143:136] <= _02509_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[135:128] <= _02508_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[127:120] <= _02507_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[119:112] <= _02506_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[111:104] <= _02505_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[103:96] <= _02504_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[95:88] <= _02623_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[87:80] <= _02612_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[79:72] <= _02600_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[71:64] <= _02589_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[63:56] <= _02578_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[55:48] <= _02567_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[47:40] <= _02556_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[39:32] <= _02545_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[31:24] <= _02534_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[23:16] <= _02523_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[15:8] <= _02512_;
  always @(posedge nvdla_core_clk)
      wt5_actv_data[7:0] <= _02601_;
  always @(posedge nvdla_core_clk)
      wt5_actv_nan <= _02629_;
  always @(posedge nvdla_core_clk)
      wt5_actv_nz <= _02630_;
  reg [0:0] \wt5_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt5_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt5_actv_pvld_reg[0]  <= wt5_actv_pvld_w;
  assign wt5_actv_pvld[0] = \wt5_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[1023:1016] <= _02241_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[1015:1008] <= _02240_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[1007:1000] <= _02239_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[999:992] <= _02366_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[991:984] <= _02365_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[983:976] <= _02364_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[975:968] <= _02363_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[967:960] <= _02362_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[959:952] <= _02360_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[951:944] <= _02359_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[943:936] <= _02358_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[935:928] <= _02357_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[927:920] <= _02356_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[919:912] <= _02355_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[911:904] <= _02354_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[903:896] <= _02353_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[895:888] <= _02352_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[887:880] <= _02351_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[879:872] <= _02349_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[871:864] <= _02348_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[863:856] <= _02347_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[855:848] <= _02346_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[847:840] <= _02345_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[839:832] <= _02344_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[831:824] <= _02343_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[823:816] <= _02342_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[815:808] <= _02341_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[807:800] <= _02340_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[799:792] <= _02337_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[791:784] <= _02336_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[783:776] <= _02335_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[775:768] <= _02334_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[767:760] <= _02333_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[759:752] <= _02332_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[751:744] <= _02331_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[743:736] <= _02330_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[735:728] <= _02329_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[727:720] <= _02328_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[719:712] <= _02326_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[711:704] <= _02325_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[703:696] <= _02324_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[695:688] <= _02323_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[687:680] <= _02322_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[679:672] <= _02321_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[671:664] <= _02320_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[663:656] <= _02319_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[655:648] <= _02318_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[647:640] <= _02317_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[639:632] <= _02315_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[631:624] <= _02314_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[623:616] <= _02313_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[615:608] <= _02312_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[607:600] <= _02311_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[599:592] <= _02310_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[591:584] <= _02309_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[583:576] <= _02308_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[575:568] <= _02307_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[567:560] <= _02306_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[559:552] <= _02304_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[551:544] <= _02303_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[543:536] <= _02302_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[535:528] <= _02301_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[527:520] <= _02300_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[519:512] <= _02299_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[511:504] <= _02298_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[503:496] <= _02297_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[495:488] <= _02296_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[487:480] <= _02295_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[479:472] <= _02293_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[471:464] <= _02292_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[463:456] <= _02291_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[455:448] <= _02290_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[447:440] <= _02289_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[439:432] <= _02288_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[431:424] <= _02287_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[423:416] <= _02286_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[415:408] <= _02285_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[407:400] <= _02284_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[399:392] <= _02282_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[391:384] <= _02281_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[383:376] <= _02280_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[375:368] <= _02279_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[367:360] <= _02278_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[359:352] <= _02277_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[351:344] <= _02276_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[343:336] <= _02275_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[335:328] <= _02274_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[327:320] <= _02273_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[319:312] <= _02271_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[311:304] <= _02270_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[303:296] <= _02269_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[295:288] <= _02268_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[287:280] <= _02267_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[279:272] <= _02266_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[271:264] <= _02265_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[263:256] <= _02264_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[255:248] <= _02263_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[247:240] <= _02262_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[239:232] <= _02260_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[231:224] <= _02259_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[223:216] <= _02258_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[215:208] <= _02257_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[207:200] <= _02256_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[199:192] <= _02255_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[191:184] <= _02254_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[183:176] <= _02253_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[175:168] <= _02252_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[167:160] <= _02251_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[159:152] <= _02249_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[151:144] <= _02248_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[143:136] <= _02247_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[135:128] <= _02246_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[127:120] <= _02245_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[119:112] <= _02244_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[111:104] <= _02243_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[103:96] <= _02242_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[95:88] <= _02361_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[87:80] <= _02350_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[79:72] <= _02338_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[71:64] <= _02327_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[63:56] <= _02316_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[55:48] <= _02305_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[47:40] <= _02294_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[39:32] <= _02283_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[31:24] <= _02272_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[23:16] <= _02261_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[15:8] <= _02250_;
  always @(posedge nvdla_core_clk)
      wt4_actv_data[7:0] <= _02339_;
  always @(posedge nvdla_core_clk)
      wt4_actv_nan <= _02367_;
  always @(posedge nvdla_core_clk)
      wt4_actv_nz <= _02368_;
  reg [0:0] \wt4_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt4_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt4_actv_pvld_reg[0]  <= wt4_actv_pvld_w;
  assign wt4_actv_pvld[0] = \wt4_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[1023:1016] <= _01979_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[1015:1008] <= _01978_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[1007:1000] <= _01977_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[999:992] <= _02104_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[991:984] <= _02103_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[983:976] <= _02102_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[975:968] <= _02101_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[967:960] <= _02100_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[959:952] <= _02098_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[951:944] <= _02097_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[943:936] <= _02096_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[935:928] <= _02095_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[927:920] <= _02094_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[919:912] <= _02093_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[911:904] <= _02092_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[903:896] <= _02091_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[895:888] <= _02090_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[887:880] <= _02089_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[879:872] <= _02087_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[871:864] <= _02086_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[863:856] <= _02085_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[855:848] <= _02084_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[847:840] <= _02083_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[839:832] <= _02082_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[831:824] <= _02081_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[823:816] <= _02080_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[815:808] <= _02079_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[807:800] <= _02078_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[799:792] <= _02075_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[791:784] <= _02074_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[783:776] <= _02073_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[775:768] <= _02072_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[767:760] <= _02071_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[759:752] <= _02070_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[751:744] <= _02069_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[743:736] <= _02068_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[735:728] <= _02067_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[727:720] <= _02066_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[719:712] <= _02064_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[711:704] <= _02063_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[703:696] <= _02062_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[695:688] <= _02061_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[687:680] <= _02060_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[679:672] <= _02059_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[671:664] <= _02058_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[663:656] <= _02057_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[655:648] <= _02056_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[647:640] <= _02055_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[639:632] <= _02053_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[631:624] <= _02052_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[623:616] <= _02051_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[615:608] <= _02050_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[607:600] <= _02049_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[599:592] <= _02048_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[591:584] <= _02047_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[583:576] <= _02046_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[575:568] <= _02045_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[567:560] <= _02044_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[559:552] <= _02042_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[551:544] <= _02041_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[543:536] <= _02040_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[535:528] <= _02039_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[527:520] <= _02038_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[519:512] <= _02037_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[511:504] <= _02036_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[503:496] <= _02035_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[495:488] <= _02034_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[487:480] <= _02033_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[479:472] <= _02031_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[471:464] <= _02030_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[463:456] <= _02029_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[455:448] <= _02028_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[447:440] <= _02027_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[439:432] <= _02026_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[431:424] <= _02025_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[423:416] <= _02024_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[415:408] <= _02023_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[407:400] <= _02022_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[399:392] <= _02020_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[391:384] <= _02019_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[383:376] <= _02018_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[375:368] <= _02017_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[367:360] <= _02016_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[359:352] <= _02015_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[351:344] <= _02014_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[343:336] <= _02013_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[335:328] <= _02012_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[327:320] <= _02011_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[319:312] <= _02009_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[311:304] <= _02008_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[303:296] <= _02007_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[295:288] <= _02006_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[287:280] <= _02005_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[279:272] <= _02004_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[271:264] <= _02003_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[263:256] <= _02002_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[255:248] <= _02001_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[247:240] <= _02000_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[239:232] <= _01998_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[231:224] <= _01997_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[223:216] <= _01996_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[215:208] <= _01995_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[207:200] <= _01994_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[199:192] <= _01993_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[191:184] <= _01992_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[183:176] <= _01991_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[175:168] <= _01990_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[167:160] <= _01989_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[159:152] <= _01987_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[151:144] <= _01986_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[143:136] <= _01985_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[135:128] <= _01984_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[127:120] <= _01983_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[119:112] <= _01982_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[111:104] <= _01981_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[103:96] <= _01980_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[95:88] <= _02099_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[87:80] <= _02088_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[79:72] <= _02076_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[71:64] <= _02065_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[63:56] <= _02054_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[55:48] <= _02043_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[47:40] <= _02032_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[39:32] <= _02021_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[31:24] <= _02010_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[23:16] <= _01999_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[15:8] <= _01988_;
  always @(posedge nvdla_core_clk)
      wt3_actv_data[7:0] <= _02077_;
  always @(posedge nvdla_core_clk)
      wt3_actv_nan <= _02105_;
  always @(posedge nvdla_core_clk)
      wt3_actv_nz <= _02106_;
  reg [0:0] \wt3_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt3_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt3_actv_pvld_reg[0]  <= wt3_actv_pvld_w;
  assign wt3_actv_pvld[0] = \wt3_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[1023:1016] <= _01717_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[1015:1008] <= _01716_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[1007:1000] <= _01715_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[999:992] <= _01842_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[991:984] <= _01841_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[983:976] <= _01840_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[975:968] <= _01839_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[967:960] <= _01838_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[959:952] <= _01836_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[951:944] <= _01835_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[943:936] <= _01834_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[935:928] <= _01833_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[927:920] <= _01832_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[919:912] <= _01831_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[911:904] <= _01830_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[903:896] <= _01829_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[895:888] <= _01828_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[887:880] <= _01827_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[879:872] <= _01825_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[871:864] <= _01824_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[863:856] <= _01823_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[855:848] <= _01822_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[847:840] <= _01821_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[839:832] <= _01820_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[831:824] <= _01819_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[823:816] <= _01818_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[815:808] <= _01817_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[807:800] <= _01816_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[799:792] <= _01813_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[791:784] <= _01812_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[783:776] <= _01811_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[775:768] <= _01810_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[767:760] <= _01809_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[759:752] <= _01808_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[751:744] <= _01807_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[743:736] <= _01806_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[735:728] <= _01805_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[727:720] <= _01804_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[719:712] <= _01802_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[711:704] <= _01801_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[703:696] <= _01800_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[695:688] <= _01799_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[687:680] <= _01798_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[679:672] <= _01797_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[671:664] <= _01796_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[663:656] <= _01795_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[655:648] <= _01794_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[647:640] <= _01793_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[639:632] <= _01791_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[631:624] <= _01790_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[623:616] <= _01789_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[615:608] <= _01788_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[607:600] <= _01787_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[599:592] <= _01786_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[591:584] <= _01785_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[583:576] <= _01784_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[575:568] <= _01783_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[567:560] <= _01782_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[559:552] <= _01780_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[551:544] <= _01779_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[543:536] <= _01778_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[535:528] <= _01777_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[527:520] <= _01776_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[519:512] <= _01775_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[511:504] <= _01774_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[503:496] <= _01773_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[495:488] <= _01772_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[487:480] <= _01771_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[479:472] <= _01769_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[471:464] <= _01768_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[463:456] <= _01767_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[455:448] <= _01766_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[447:440] <= _01765_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[439:432] <= _01764_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[431:424] <= _01763_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[423:416] <= _01762_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[415:408] <= _01761_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[407:400] <= _01760_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[399:392] <= _01758_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[391:384] <= _01757_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[383:376] <= _01756_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[375:368] <= _01755_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[367:360] <= _01754_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[359:352] <= _01753_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[351:344] <= _01752_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[343:336] <= _01751_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[335:328] <= _01750_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[327:320] <= _01749_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[319:312] <= _01747_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[311:304] <= _01746_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[303:296] <= _01745_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[295:288] <= _01744_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[287:280] <= _01743_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[279:272] <= _01742_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[271:264] <= _01741_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[263:256] <= _01740_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[255:248] <= _01739_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[247:240] <= _01738_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[239:232] <= _01736_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[231:224] <= _01735_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[223:216] <= _01734_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[215:208] <= _01733_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[207:200] <= _01732_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[199:192] <= _01731_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[191:184] <= _01730_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[183:176] <= _01729_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[175:168] <= _01728_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[167:160] <= _01727_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[159:152] <= _01725_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[151:144] <= _01724_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[143:136] <= _01723_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[135:128] <= _01722_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[127:120] <= _01721_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[119:112] <= _01720_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[111:104] <= _01719_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[103:96] <= _01718_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[95:88] <= _01837_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[87:80] <= _01826_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[79:72] <= _01814_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[71:64] <= _01803_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[63:56] <= _01792_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[55:48] <= _01781_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[47:40] <= _01770_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[39:32] <= _01759_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[31:24] <= _01748_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[23:16] <= _01737_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[15:8] <= _01726_;
  always @(posedge nvdla_core_clk)
      wt2_actv_data[7:0] <= _01815_;
  always @(posedge nvdla_core_clk)
      wt2_actv_nan <= _01843_;
  always @(posedge nvdla_core_clk)
      wt2_actv_nz <= _01844_;
  reg [0:0] \wt2_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt2_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt2_actv_pvld_reg[0]  <= wt2_actv_pvld_w;
  assign wt2_actv_pvld[0] = \wt2_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[1023:1016] <= _01455_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[1015:1008] <= _01454_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[1007:1000] <= _01453_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[999:992] <= _01580_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[991:984] <= _01579_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[983:976] <= _01578_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[975:968] <= _01577_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[967:960] <= _01576_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[959:952] <= _01574_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[951:944] <= _01573_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[943:936] <= _01572_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[935:928] <= _01571_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[927:920] <= _01570_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[919:912] <= _01569_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[911:904] <= _01568_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[903:896] <= _01567_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[895:888] <= _01566_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[887:880] <= _01565_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[879:872] <= _01563_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[871:864] <= _01562_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[863:856] <= _01561_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[855:848] <= _01560_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[847:840] <= _01559_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[839:832] <= _01558_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[831:824] <= _01557_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[823:816] <= _01556_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[815:808] <= _01555_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[807:800] <= _01554_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[799:792] <= _01551_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[791:784] <= _01550_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[783:776] <= _01549_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[775:768] <= _01548_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[767:760] <= _01547_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[759:752] <= _01546_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[751:744] <= _01545_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[743:736] <= _01544_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[735:728] <= _01543_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[727:720] <= _01542_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[719:712] <= _01540_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[711:704] <= _01539_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[703:696] <= _01538_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[695:688] <= _01537_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[687:680] <= _01536_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[679:672] <= _01535_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[671:664] <= _01534_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[663:656] <= _01533_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[655:648] <= _01532_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[647:640] <= _01531_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[639:632] <= _01529_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[631:624] <= _01528_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[623:616] <= _01527_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[615:608] <= _01526_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[607:600] <= _01525_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[599:592] <= _01524_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[591:584] <= _01523_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[583:576] <= _01522_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[575:568] <= _01521_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[567:560] <= _01520_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[559:552] <= _01518_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[551:544] <= _01517_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[543:536] <= _01516_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[535:528] <= _01515_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[527:520] <= _01514_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[519:512] <= _01513_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[511:504] <= _01512_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[503:496] <= _01511_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[495:488] <= _01510_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[487:480] <= _01509_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[479:472] <= _01507_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[471:464] <= _01506_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[463:456] <= _01505_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[455:448] <= _01504_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[447:440] <= _01503_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[439:432] <= _01502_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[431:424] <= _01501_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[423:416] <= _01500_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[415:408] <= _01499_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[407:400] <= _01498_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[399:392] <= _01496_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[391:384] <= _01495_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[383:376] <= _01494_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[375:368] <= _01493_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[367:360] <= _01492_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[359:352] <= _01491_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[351:344] <= _01490_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[343:336] <= _01489_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[335:328] <= _01488_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[327:320] <= _01487_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[319:312] <= _01485_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[311:304] <= _01484_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[303:296] <= _01483_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[295:288] <= _01482_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[287:280] <= _01481_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[279:272] <= _01480_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[271:264] <= _01479_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[263:256] <= _01478_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[255:248] <= _01477_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[247:240] <= _01476_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[239:232] <= _01474_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[231:224] <= _01473_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[223:216] <= _01472_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[215:208] <= _01471_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[207:200] <= _01470_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[199:192] <= _01469_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[191:184] <= _01468_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[183:176] <= _01467_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[175:168] <= _01466_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[167:160] <= _01465_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[159:152] <= _01463_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[151:144] <= _01462_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[143:136] <= _01461_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[135:128] <= _01460_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[127:120] <= _01459_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[119:112] <= _01458_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[111:104] <= _01457_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[103:96] <= _01456_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[95:88] <= _01575_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[87:80] <= _01564_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[79:72] <= _01552_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[71:64] <= _01541_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[63:56] <= _01530_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[55:48] <= _01519_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[47:40] <= _01508_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[39:32] <= _01497_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[31:24] <= _01486_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[23:16] <= _01475_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[15:8] <= _01464_;
  always @(posedge nvdla_core_clk)
      wt1_actv_data[7:0] <= _01553_;
  always @(posedge nvdla_core_clk)
      wt1_actv_nan <= _01581_;
  always @(posedge nvdla_core_clk)
      wt1_actv_nz <= _01582_;
  reg [0:0] \wt1_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt1_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt1_actv_pvld_reg[0]  <= wt1_actv_pvld_w;
  assign wt1_actv_pvld[0] = \wt1_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[1023:1016] <= _01193_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[1015:1008] <= _01192_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[1007:1000] <= _01191_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[999:992] <= _01318_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[991:984] <= _01317_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[983:976] <= _01316_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[975:968] <= _01315_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[967:960] <= _01314_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[959:952] <= _01312_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[951:944] <= _01311_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[943:936] <= _01310_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[935:928] <= _01309_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[927:920] <= _01308_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[919:912] <= _01307_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[911:904] <= _01306_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[903:896] <= _01305_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[895:888] <= _01304_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[887:880] <= _01303_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[879:872] <= _01301_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[871:864] <= _01300_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[863:856] <= _01299_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[855:848] <= _01298_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[847:840] <= _01297_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[839:832] <= _01296_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[831:824] <= _01295_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[823:816] <= _01294_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[815:808] <= _01293_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[807:800] <= _01292_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[799:792] <= _01289_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[791:784] <= _01288_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[783:776] <= _01287_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[775:768] <= _01286_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[767:760] <= _01285_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[759:752] <= _01284_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[751:744] <= _01283_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[743:736] <= _01282_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[735:728] <= _01281_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[727:720] <= _01280_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[719:712] <= _01278_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[711:704] <= _01277_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[703:696] <= _01276_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[695:688] <= _01275_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[687:680] <= _01274_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[679:672] <= _01273_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[671:664] <= _01272_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[663:656] <= _01271_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[655:648] <= _01270_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[647:640] <= _01269_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[639:632] <= _01267_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[631:624] <= _01266_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[623:616] <= _01265_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[615:608] <= _01264_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[607:600] <= _01263_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[599:592] <= _01262_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[591:584] <= _01261_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[583:576] <= _01260_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[575:568] <= _01259_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[567:560] <= _01258_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[559:552] <= _01256_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[551:544] <= _01255_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[543:536] <= _01254_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[535:528] <= _01253_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[527:520] <= _01252_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[519:512] <= _01251_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[511:504] <= _01250_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[503:496] <= _01249_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[495:488] <= _01248_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[487:480] <= _01247_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[479:472] <= _01245_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[471:464] <= _01244_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[463:456] <= _01243_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[455:448] <= _01242_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[447:440] <= _01241_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[439:432] <= _01240_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[431:424] <= _01239_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[423:416] <= _01238_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[415:408] <= _01237_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[407:400] <= _01236_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[399:392] <= _01234_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[391:384] <= _01233_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[383:376] <= _01232_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[375:368] <= _01231_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[367:360] <= _01230_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[359:352] <= _01229_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[351:344] <= _01228_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[343:336] <= _01227_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[335:328] <= _01226_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[327:320] <= _01225_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[319:312] <= _01223_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[311:304] <= _01222_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[303:296] <= _01221_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[295:288] <= _01220_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[287:280] <= _01219_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[279:272] <= _01218_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[271:264] <= _01217_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[263:256] <= _01216_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[255:248] <= _01215_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[247:240] <= _01214_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[239:232] <= _01212_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[231:224] <= _01211_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[223:216] <= _01210_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[215:208] <= _01209_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[207:200] <= _01208_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[199:192] <= _01207_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[191:184] <= _01206_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[183:176] <= _01205_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[175:168] <= _01204_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[167:160] <= _01203_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[159:152] <= _01201_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[151:144] <= _01200_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[143:136] <= _01199_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[135:128] <= _01198_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[127:120] <= _01197_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[119:112] <= _01196_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[111:104] <= _01195_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[103:96] <= _01194_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[95:88] <= _01313_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[87:80] <= _01302_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[79:72] <= _01290_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[71:64] <= _01279_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[63:56] <= _01268_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[55:48] <= _01257_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[47:40] <= _01246_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[39:32] <= _01235_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[31:24] <= _01224_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[23:16] <= _01213_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[15:8] <= _01202_;
  always @(posedge nvdla_core_clk)
      wt0_actv_data[7:0] <= _01291_;
  always @(posedge nvdla_core_clk)
      wt0_actv_nan <= _01319_;
  always @(posedge nvdla_core_clk)
      wt0_actv_nz <= _01320_;
  reg [0:0] \wt0_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \wt0_actv_pvld_reg[0]  <= 1'b0;
    else
      \wt0_actv_pvld_reg[0]  <= wt0_actv_pvld_w;
  assign wt0_actv_pvld[0] = \wt0_actv_pvld_reg[0] ;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[1023:1016] <= _03157_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[1015:1008] <= _03156_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[1007:1000] <= _03155_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[999:992] <= _03282_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[991:984] <= _03281_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[983:976] <= _03280_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[975:968] <= _03279_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[967:960] <= _03278_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[959:952] <= _03276_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[951:944] <= _03275_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[943:936] <= _03274_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[935:928] <= _03273_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[927:920] <= _03272_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[919:912] <= _03271_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[911:904] <= _03270_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[903:896] <= _03269_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[895:888] <= _03268_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[887:880] <= _03267_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[879:872] <= _03265_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[871:864] <= _03264_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[863:856] <= _03263_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[855:848] <= _03262_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[847:840] <= _03261_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[839:832] <= _03260_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[831:824] <= _03259_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[823:816] <= _03258_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[815:808] <= _03257_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[807:800] <= _03256_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[799:792] <= _03253_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[791:784] <= _03252_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[783:776] <= _03251_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[775:768] <= _03250_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[767:760] <= _03249_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[759:752] <= _03248_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[751:744] <= _03247_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[743:736] <= _03246_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[735:728] <= _03245_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[727:720] <= _03244_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[719:712] <= _03242_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[711:704] <= _03241_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[703:696] <= _03240_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[695:688] <= _03239_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[687:680] <= _03238_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[679:672] <= _03237_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[671:664] <= _03236_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[663:656] <= _03235_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[655:648] <= _03234_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[647:640] <= _03233_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[639:632] <= _03231_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[631:624] <= _03230_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[623:616] <= _03229_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[615:608] <= _03228_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[607:600] <= _03227_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[599:592] <= _03226_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[591:584] <= _03225_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[583:576] <= _03224_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[575:568] <= _03223_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[567:560] <= _03222_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[559:552] <= _03220_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[551:544] <= _03219_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[543:536] <= _03218_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[535:528] <= _03217_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[527:520] <= _03216_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[519:512] <= _03215_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[511:504] <= _03214_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[503:496] <= _03213_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[495:488] <= _03212_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[487:480] <= _03211_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[479:472] <= _03209_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[471:464] <= _03208_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[463:456] <= _03207_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[455:448] <= _03206_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[447:440] <= _03205_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[439:432] <= _03204_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[431:424] <= _03203_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[423:416] <= _03202_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[415:408] <= _03201_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[407:400] <= _03200_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[399:392] <= _03198_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[391:384] <= _03197_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[383:376] <= _03196_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[375:368] <= _03195_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[367:360] <= _03194_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[359:352] <= _03193_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[351:344] <= _03192_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[343:336] <= _03191_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[335:328] <= _03190_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[327:320] <= _03189_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[319:312] <= _03187_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[311:304] <= _03186_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[303:296] <= _03185_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[295:288] <= _03184_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[287:280] <= _03183_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[279:272] <= _03182_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[271:264] <= _03181_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[263:256] <= _03180_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[255:248] <= _03179_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[247:240] <= _03178_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[239:232] <= _03176_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[231:224] <= _03175_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[223:216] <= _03174_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[215:208] <= _03173_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[207:200] <= _03172_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[199:192] <= _03171_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[191:184] <= _03170_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[183:176] <= _03169_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[175:168] <= _03168_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[167:160] <= _03167_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[159:152] <= _03165_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[151:144] <= _03164_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[143:136] <= _03163_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[135:128] <= _03162_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[127:120] <= _03161_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[119:112] <= _03160_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[111:104] <= _03159_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[103:96] <= _03158_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[95:88] <= _03277_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[87:80] <= _03266_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[79:72] <= _03254_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[71:64] <= _03243_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[63:56] <= _03232_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[55:48] <= _03221_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[47:40] <= _03210_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[39:32] <= _03199_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[31:24] <= _03188_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[23:16] <= _03177_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[15:8] <= _03166_;
  always @(posedge nvdla_core_clk)
      wt7_sd_data[7:0] <= _03255_;
  always @(posedge nvdla_core_clk)
      wt7_sd_nan <= _03285_;
  always @(posedge nvdla_core_clk)
      wt7_sd_exp <= _03283_;
  always @(posedge nvdla_core_clk)
      wt7_sd_mask <= _03284_;
  always @(posedge nvdla_core_clk)
      wt7_sd_nz <= _03286_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt7_sd_pvld <= 1'b0;
    else
      wt7_sd_pvld <= wt7_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[1023:1016] <= _02895_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[1015:1008] <= _02894_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[1007:1000] <= _02893_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[999:992] <= _03020_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[991:984] <= _03019_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[983:976] <= _03018_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[975:968] <= _03017_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[967:960] <= _03016_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[959:952] <= _03014_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[951:944] <= _03013_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[943:936] <= _03012_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[935:928] <= _03011_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[927:920] <= _03010_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[919:912] <= _03009_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[911:904] <= _03008_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[903:896] <= _03007_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[895:888] <= _03006_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[887:880] <= _03005_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[879:872] <= _03003_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[871:864] <= _03002_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[863:856] <= _03001_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[855:848] <= _03000_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[847:840] <= _02999_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[839:832] <= _02998_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[831:824] <= _02997_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[823:816] <= _02996_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[815:808] <= _02995_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[807:800] <= _02994_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[799:792] <= _02991_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[791:784] <= _02990_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[783:776] <= _02989_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[775:768] <= _02988_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[767:760] <= _02987_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[759:752] <= _02986_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[751:744] <= _02985_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[743:736] <= _02984_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[735:728] <= _02983_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[727:720] <= _02982_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[719:712] <= _02980_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[711:704] <= _02979_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[703:696] <= _02978_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[695:688] <= _02977_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[687:680] <= _02976_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[679:672] <= _02975_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[671:664] <= _02974_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[663:656] <= _02973_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[655:648] <= _02972_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[647:640] <= _02971_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[639:632] <= _02969_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[631:624] <= _02968_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[623:616] <= _02967_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[615:608] <= _02966_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[607:600] <= _02965_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[599:592] <= _02964_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[591:584] <= _02963_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[583:576] <= _02962_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[575:568] <= _02961_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[567:560] <= _02960_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[559:552] <= _02958_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[551:544] <= _02957_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[543:536] <= _02956_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[535:528] <= _02955_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[527:520] <= _02954_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[519:512] <= _02953_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[511:504] <= _02952_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[503:496] <= _02951_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[495:488] <= _02950_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[487:480] <= _02949_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[479:472] <= _02947_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[471:464] <= _02946_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[463:456] <= _02945_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[455:448] <= _02944_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[447:440] <= _02943_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[439:432] <= _02942_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[431:424] <= _02941_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[423:416] <= _02940_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[415:408] <= _02939_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[407:400] <= _02938_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[399:392] <= _02936_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[391:384] <= _02935_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[383:376] <= _02934_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[375:368] <= _02933_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[367:360] <= _02932_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[359:352] <= _02931_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[351:344] <= _02930_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[343:336] <= _02929_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[335:328] <= _02928_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[327:320] <= _02927_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[319:312] <= _02925_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[311:304] <= _02924_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[303:296] <= _02923_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[295:288] <= _02922_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[287:280] <= _02921_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[279:272] <= _02920_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[271:264] <= _02919_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[263:256] <= _02918_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[255:248] <= _02917_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[247:240] <= _02916_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[239:232] <= _02914_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[231:224] <= _02913_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[223:216] <= _02912_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[215:208] <= _02911_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[207:200] <= _02910_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[199:192] <= _02909_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[191:184] <= _02908_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[183:176] <= _02907_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[175:168] <= _02906_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[167:160] <= _02905_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[159:152] <= _02903_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[151:144] <= _02902_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[143:136] <= _02901_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[135:128] <= _02900_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[127:120] <= _02899_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[119:112] <= _02898_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[111:104] <= _02897_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[103:96] <= _02896_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[95:88] <= _03015_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[87:80] <= _03004_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[79:72] <= _02992_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[71:64] <= _02981_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[63:56] <= _02970_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[55:48] <= _02959_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[47:40] <= _02948_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[39:32] <= _02937_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[31:24] <= _02926_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[23:16] <= _02915_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[15:8] <= _02904_;
  always @(posedge nvdla_core_clk)
      wt6_sd_data[7:0] <= _02993_;
  always @(posedge nvdla_core_clk)
      wt6_sd_nan <= _03023_;
  always @(posedge nvdla_core_clk)
      wt6_sd_exp <= _03021_;
  always @(posedge nvdla_core_clk)
      wt6_sd_mask <= _03022_;
  always @(posedge nvdla_core_clk)
      wt6_sd_nz <= _03024_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt6_sd_pvld <= 1'b0;
    else
      wt6_sd_pvld <= wt6_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[1023:1016] <= _02633_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[1015:1008] <= _02632_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[1007:1000] <= _02631_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[999:992] <= _02758_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[991:984] <= _02757_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[983:976] <= _02756_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[975:968] <= _02755_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[967:960] <= _02754_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[959:952] <= _02752_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[951:944] <= _02751_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[943:936] <= _02750_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[935:928] <= _02749_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[927:920] <= _02748_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[919:912] <= _02747_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[911:904] <= _02746_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[903:896] <= _02745_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[895:888] <= _02744_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[887:880] <= _02743_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[879:872] <= _02741_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[871:864] <= _02740_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[863:856] <= _02739_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[855:848] <= _02738_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[847:840] <= _02737_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[839:832] <= _02736_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[831:824] <= _02735_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[823:816] <= _02734_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[815:808] <= _02733_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[807:800] <= _02732_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[799:792] <= _02729_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[791:784] <= _02728_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[783:776] <= _02727_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[775:768] <= _02726_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[767:760] <= _02725_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[759:752] <= _02724_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[751:744] <= _02723_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[743:736] <= _02722_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[735:728] <= _02721_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[727:720] <= _02720_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[719:712] <= _02718_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[711:704] <= _02717_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[703:696] <= _02716_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[695:688] <= _02715_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[687:680] <= _02714_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[679:672] <= _02713_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[671:664] <= _02712_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[663:656] <= _02711_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[655:648] <= _02710_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[647:640] <= _02709_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[639:632] <= _02707_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[631:624] <= _02706_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[623:616] <= _02705_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[615:608] <= _02704_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[607:600] <= _02703_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[599:592] <= _02702_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[591:584] <= _02701_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[583:576] <= _02700_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[575:568] <= _02699_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[567:560] <= _02698_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[559:552] <= _02696_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[551:544] <= _02695_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[543:536] <= _02694_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[535:528] <= _02693_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[527:520] <= _02692_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[519:512] <= _02691_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[511:504] <= _02690_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[503:496] <= _02689_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[495:488] <= _02688_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[487:480] <= _02687_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[479:472] <= _02685_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[471:464] <= _02684_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[463:456] <= _02683_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[455:448] <= _02682_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[447:440] <= _02681_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[439:432] <= _02680_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[431:424] <= _02679_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[423:416] <= _02678_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[415:408] <= _02677_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[407:400] <= _02676_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[399:392] <= _02674_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[391:384] <= _02673_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[383:376] <= _02672_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[375:368] <= _02671_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[367:360] <= _02670_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[359:352] <= _02669_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[351:344] <= _02668_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[343:336] <= _02667_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[335:328] <= _02666_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[327:320] <= _02665_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[319:312] <= _02663_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[311:304] <= _02662_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[303:296] <= _02661_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[295:288] <= _02660_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[287:280] <= _02659_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[279:272] <= _02658_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[271:264] <= _02657_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[263:256] <= _02656_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[255:248] <= _02655_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[247:240] <= _02654_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[239:232] <= _02652_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[231:224] <= _02651_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[223:216] <= _02650_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[215:208] <= _02649_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[207:200] <= _02648_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[199:192] <= _02647_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[191:184] <= _02646_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[183:176] <= _02645_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[175:168] <= _02644_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[167:160] <= _02643_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[159:152] <= _02641_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[151:144] <= _02640_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[143:136] <= _02639_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[135:128] <= _02638_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[127:120] <= _02637_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[119:112] <= _02636_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[111:104] <= _02635_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[103:96] <= _02634_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[95:88] <= _02753_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[87:80] <= _02742_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[79:72] <= _02730_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[71:64] <= _02719_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[63:56] <= _02708_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[55:48] <= _02697_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[47:40] <= _02686_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[39:32] <= _02675_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[31:24] <= _02664_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[23:16] <= _02653_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[15:8] <= _02642_;
  always @(posedge nvdla_core_clk)
      wt5_sd_data[7:0] <= _02731_;
  always @(posedge nvdla_core_clk)
      wt5_sd_nan <= _02761_;
  always @(posedge nvdla_core_clk)
      wt5_sd_exp <= _02759_;
  always @(posedge nvdla_core_clk)
      wt5_sd_mask <= _02760_;
  always @(posedge nvdla_core_clk)
      wt5_sd_nz <= _02762_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt5_sd_pvld <= 1'b0;
    else
      wt5_sd_pvld <= wt5_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[1023:1016] <= _02371_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[1015:1008] <= _02370_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[1007:1000] <= _02369_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[999:992] <= _02496_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[991:984] <= _02495_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[983:976] <= _02494_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[975:968] <= _02493_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[967:960] <= _02492_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[959:952] <= _02490_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[951:944] <= _02489_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[943:936] <= _02488_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[935:928] <= _02487_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[927:920] <= _02486_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[919:912] <= _02485_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[911:904] <= _02484_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[903:896] <= _02483_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[895:888] <= _02482_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[887:880] <= _02481_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[879:872] <= _02479_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[871:864] <= _02478_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[863:856] <= _02477_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[855:848] <= _02476_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[847:840] <= _02475_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[839:832] <= _02474_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[831:824] <= _02473_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[823:816] <= _02472_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[815:808] <= _02471_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[807:800] <= _02470_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[799:792] <= _02467_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[791:784] <= _02466_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[783:776] <= _02465_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[775:768] <= _02464_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[767:760] <= _02463_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[759:752] <= _02462_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[751:744] <= _02461_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[743:736] <= _02460_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[735:728] <= _02459_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[727:720] <= _02458_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[719:712] <= _02456_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[711:704] <= _02455_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[703:696] <= _02454_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[695:688] <= _02453_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[687:680] <= _02452_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[679:672] <= _02451_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[671:664] <= _02450_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[663:656] <= _02449_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[655:648] <= _02448_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[647:640] <= _02447_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[639:632] <= _02445_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[631:624] <= _02444_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[623:616] <= _02443_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[615:608] <= _02442_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[607:600] <= _02441_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[599:592] <= _02440_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[591:584] <= _02439_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[583:576] <= _02438_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[575:568] <= _02437_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[567:560] <= _02436_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[559:552] <= _02434_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[551:544] <= _02433_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[543:536] <= _02432_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[535:528] <= _02431_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[527:520] <= _02430_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[519:512] <= _02429_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[511:504] <= _02428_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[503:496] <= _02427_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[495:488] <= _02426_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[487:480] <= _02425_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[479:472] <= _02423_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[471:464] <= _02422_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[463:456] <= _02421_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[455:448] <= _02420_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[447:440] <= _02419_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[439:432] <= _02418_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[431:424] <= _02417_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[423:416] <= _02416_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[415:408] <= _02415_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[407:400] <= _02414_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[399:392] <= _02412_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[391:384] <= _02411_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[383:376] <= _02410_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[375:368] <= _02409_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[367:360] <= _02408_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[359:352] <= _02407_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[351:344] <= _02406_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[343:336] <= _02405_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[335:328] <= _02404_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[327:320] <= _02403_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[319:312] <= _02401_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[311:304] <= _02400_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[303:296] <= _02399_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[295:288] <= _02398_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[287:280] <= _02397_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[279:272] <= _02396_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[271:264] <= _02395_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[263:256] <= _02394_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[255:248] <= _02393_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[247:240] <= _02392_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[239:232] <= _02390_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[231:224] <= _02389_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[223:216] <= _02388_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[215:208] <= _02387_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[207:200] <= _02386_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[199:192] <= _02385_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[191:184] <= _02384_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[183:176] <= _02383_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[175:168] <= _02382_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[167:160] <= _02381_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[159:152] <= _02379_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[151:144] <= _02378_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[143:136] <= _02377_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[135:128] <= _02376_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[127:120] <= _02375_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[119:112] <= _02374_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[111:104] <= _02373_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[103:96] <= _02372_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[95:88] <= _02491_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[87:80] <= _02480_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[79:72] <= _02468_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[71:64] <= _02457_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[63:56] <= _02446_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[55:48] <= _02435_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[47:40] <= _02424_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[39:32] <= _02413_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[31:24] <= _02402_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[23:16] <= _02391_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[15:8] <= _02380_;
  always @(posedge nvdla_core_clk)
      wt4_sd_data[7:0] <= _02469_;
  always @(posedge nvdla_core_clk)
      wt4_sd_nan <= _02499_;
  always @(posedge nvdla_core_clk)
      wt4_sd_exp <= _02497_;
  always @(posedge nvdla_core_clk)
      wt4_sd_mask <= _02498_;
  always @(posedge nvdla_core_clk)
      wt4_sd_nz <= _02500_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt4_sd_pvld <= 1'b0;
    else
      wt4_sd_pvld <= wt4_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[1023:1016] <= _02109_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[1015:1008] <= _02108_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[1007:1000] <= _02107_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[999:992] <= _02234_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[991:984] <= _02233_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[983:976] <= _02232_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[975:968] <= _02231_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[967:960] <= _02230_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[959:952] <= _02228_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[951:944] <= _02227_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[943:936] <= _02226_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[935:928] <= _02225_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[927:920] <= _02224_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[919:912] <= _02223_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[911:904] <= _02222_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[903:896] <= _02221_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[895:888] <= _02220_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[887:880] <= _02219_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[879:872] <= _02217_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[871:864] <= _02216_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[863:856] <= _02215_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[855:848] <= _02214_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[847:840] <= _02213_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[839:832] <= _02212_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[831:824] <= _02211_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[823:816] <= _02210_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[815:808] <= _02209_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[807:800] <= _02208_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[799:792] <= _02205_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[791:784] <= _02204_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[783:776] <= _02203_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[775:768] <= _02202_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[767:760] <= _02201_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[759:752] <= _02200_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[751:744] <= _02199_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[743:736] <= _02198_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[735:728] <= _02197_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[727:720] <= _02196_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[719:712] <= _02194_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[711:704] <= _02193_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[703:696] <= _02192_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[695:688] <= _02191_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[687:680] <= _02190_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[679:672] <= _02189_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[671:664] <= _02188_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[663:656] <= _02187_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[655:648] <= _02186_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[647:640] <= _02185_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[639:632] <= _02183_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[631:624] <= _02182_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[623:616] <= _02181_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[615:608] <= _02180_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[607:600] <= _02179_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[599:592] <= _02178_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[591:584] <= _02177_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[583:576] <= _02176_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[575:568] <= _02175_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[567:560] <= _02174_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[559:552] <= _02172_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[551:544] <= _02171_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[543:536] <= _02170_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[535:528] <= _02169_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[527:520] <= _02168_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[519:512] <= _02167_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[511:504] <= _02166_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[503:496] <= _02165_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[495:488] <= _02164_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[487:480] <= _02163_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[479:472] <= _02161_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[471:464] <= _02160_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[463:456] <= _02159_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[455:448] <= _02158_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[447:440] <= _02157_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[439:432] <= _02156_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[431:424] <= _02155_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[423:416] <= _02154_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[415:408] <= _02153_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[407:400] <= _02152_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[399:392] <= _02150_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[391:384] <= _02149_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[383:376] <= _02148_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[375:368] <= _02147_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[367:360] <= _02146_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[359:352] <= _02145_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[351:344] <= _02144_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[343:336] <= _02143_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[335:328] <= _02142_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[327:320] <= _02141_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[319:312] <= _02139_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[311:304] <= _02138_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[303:296] <= _02137_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[295:288] <= _02136_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[287:280] <= _02135_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[279:272] <= _02134_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[271:264] <= _02133_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[263:256] <= _02132_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[255:248] <= _02131_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[247:240] <= _02130_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[239:232] <= _02128_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[231:224] <= _02127_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[223:216] <= _02126_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[215:208] <= _02125_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[207:200] <= _02124_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[199:192] <= _02123_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[191:184] <= _02122_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[183:176] <= _02121_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[175:168] <= _02120_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[167:160] <= _02119_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[159:152] <= _02117_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[151:144] <= _02116_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[143:136] <= _02115_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[135:128] <= _02114_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[127:120] <= _02113_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[119:112] <= _02112_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[111:104] <= _02111_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[103:96] <= _02110_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[95:88] <= _02229_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[87:80] <= _02218_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[79:72] <= _02206_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[71:64] <= _02195_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[63:56] <= _02184_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[55:48] <= _02173_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[47:40] <= _02162_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[39:32] <= _02151_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[31:24] <= _02140_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[23:16] <= _02129_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[15:8] <= _02118_;
  always @(posedge nvdla_core_clk)
      wt3_sd_data[7:0] <= _02207_;
  always @(posedge nvdla_core_clk)
      wt3_sd_nan <= _02237_;
  always @(posedge nvdla_core_clk)
      wt3_sd_exp <= _02235_;
  always @(posedge nvdla_core_clk)
      wt3_sd_mask <= _02236_;
  always @(posedge nvdla_core_clk)
      wt3_sd_nz <= _02238_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt3_sd_pvld <= 1'b0;
    else
      wt3_sd_pvld <= wt3_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[1023:1016] <= _01847_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[1015:1008] <= _01846_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[1007:1000] <= _01845_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[999:992] <= _01972_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[991:984] <= _01971_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[983:976] <= _01970_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[975:968] <= _01969_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[967:960] <= _01968_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[959:952] <= _01966_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[951:944] <= _01965_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[943:936] <= _01964_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[935:928] <= _01963_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[927:920] <= _01962_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[919:912] <= _01961_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[911:904] <= _01960_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[903:896] <= _01959_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[895:888] <= _01958_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[887:880] <= _01957_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[879:872] <= _01955_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[871:864] <= _01954_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[863:856] <= _01953_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[855:848] <= _01952_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[847:840] <= _01951_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[839:832] <= _01950_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[831:824] <= _01949_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[823:816] <= _01948_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[815:808] <= _01947_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[807:800] <= _01946_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[799:792] <= _01943_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[791:784] <= _01942_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[783:776] <= _01941_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[775:768] <= _01940_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[767:760] <= _01939_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[759:752] <= _01938_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[751:744] <= _01937_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[743:736] <= _01936_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[735:728] <= _01935_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[727:720] <= _01934_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[719:712] <= _01932_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[711:704] <= _01931_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[703:696] <= _01930_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[695:688] <= _01929_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[687:680] <= _01928_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[679:672] <= _01927_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[671:664] <= _01926_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[663:656] <= _01925_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[655:648] <= _01924_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[647:640] <= _01923_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[639:632] <= _01921_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[631:624] <= _01920_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[623:616] <= _01919_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[615:608] <= _01918_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[607:600] <= _01917_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[599:592] <= _01916_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[591:584] <= _01915_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[583:576] <= _01914_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[575:568] <= _01913_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[567:560] <= _01912_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[559:552] <= _01910_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[551:544] <= _01909_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[543:536] <= _01908_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[535:528] <= _01907_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[527:520] <= _01906_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[519:512] <= _01905_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[511:504] <= _01904_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[503:496] <= _01903_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[495:488] <= _01902_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[487:480] <= _01901_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[479:472] <= _01899_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[471:464] <= _01898_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[463:456] <= _01897_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[455:448] <= _01896_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[447:440] <= _01895_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[439:432] <= _01894_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[431:424] <= _01893_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[423:416] <= _01892_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[415:408] <= _01891_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[407:400] <= _01890_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[399:392] <= _01888_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[391:384] <= _01887_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[383:376] <= _01886_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[375:368] <= _01885_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[367:360] <= _01884_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[359:352] <= _01883_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[351:344] <= _01882_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[343:336] <= _01881_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[335:328] <= _01880_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[327:320] <= _01879_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[319:312] <= _01877_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[311:304] <= _01876_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[303:296] <= _01875_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[295:288] <= _01874_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[287:280] <= _01873_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[279:272] <= _01872_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[271:264] <= _01871_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[263:256] <= _01870_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[255:248] <= _01869_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[247:240] <= _01868_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[239:232] <= _01866_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[231:224] <= _01865_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[223:216] <= _01864_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[215:208] <= _01863_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[207:200] <= _01862_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[199:192] <= _01861_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[191:184] <= _01860_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[183:176] <= _01859_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[175:168] <= _01858_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[167:160] <= _01857_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[159:152] <= _01855_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[151:144] <= _01854_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[143:136] <= _01853_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[135:128] <= _01852_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[127:120] <= _01851_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[119:112] <= _01850_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[111:104] <= _01849_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[103:96] <= _01848_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[95:88] <= _01967_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[87:80] <= _01956_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[79:72] <= _01944_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[71:64] <= _01933_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[63:56] <= _01922_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[55:48] <= _01911_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[47:40] <= _01900_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[39:32] <= _01889_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[31:24] <= _01878_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[23:16] <= _01867_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[15:8] <= _01856_;
  always @(posedge nvdla_core_clk)
      wt2_sd_data[7:0] <= _01945_;
  always @(posedge nvdla_core_clk)
      wt2_sd_nan <= _01975_;
  always @(posedge nvdla_core_clk)
      wt2_sd_exp <= _01973_;
  always @(posedge nvdla_core_clk)
      wt2_sd_mask <= _01974_;
  always @(posedge nvdla_core_clk)
      wt2_sd_nz <= _01976_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt2_sd_pvld <= 1'b0;
    else
      wt2_sd_pvld <= wt2_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[1023:1016] <= _01585_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[1015:1008] <= _01584_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[1007:1000] <= _01583_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[999:992] <= _01710_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[991:984] <= _01709_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[983:976] <= _01708_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[975:968] <= _01707_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[967:960] <= _01706_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[959:952] <= _01704_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[951:944] <= _01703_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[943:936] <= _01702_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[935:928] <= _01701_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[927:920] <= _01700_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[919:912] <= _01699_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[911:904] <= _01698_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[903:896] <= _01697_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[895:888] <= _01696_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[887:880] <= _01695_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[879:872] <= _01693_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[871:864] <= _01692_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[863:856] <= _01691_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[855:848] <= _01690_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[847:840] <= _01689_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[839:832] <= _01688_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[831:824] <= _01687_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[823:816] <= _01686_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[815:808] <= _01685_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[807:800] <= _01684_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[799:792] <= _01681_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[791:784] <= _01680_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[783:776] <= _01679_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[775:768] <= _01678_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[767:760] <= _01677_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[759:752] <= _01676_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[751:744] <= _01675_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[743:736] <= _01674_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[735:728] <= _01673_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[727:720] <= _01672_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[719:712] <= _01670_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[711:704] <= _01669_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[703:696] <= _01668_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[695:688] <= _01667_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[687:680] <= _01666_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[679:672] <= _01665_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[671:664] <= _01664_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[663:656] <= _01663_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[655:648] <= _01662_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[647:640] <= _01661_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[639:632] <= _01659_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[631:624] <= _01658_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[623:616] <= _01657_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[615:608] <= _01656_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[607:600] <= _01655_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[599:592] <= _01654_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[591:584] <= _01653_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[583:576] <= _01652_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[575:568] <= _01651_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[567:560] <= _01650_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[559:552] <= _01648_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[551:544] <= _01647_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[543:536] <= _01646_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[535:528] <= _01645_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[527:520] <= _01644_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[519:512] <= _01643_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[511:504] <= _01642_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[503:496] <= _01641_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[495:488] <= _01640_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[487:480] <= _01639_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[479:472] <= _01637_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[471:464] <= _01636_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[463:456] <= _01635_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[455:448] <= _01634_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[447:440] <= _01633_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[439:432] <= _01632_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[431:424] <= _01631_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[423:416] <= _01630_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[415:408] <= _01629_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[407:400] <= _01628_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[399:392] <= _01626_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[391:384] <= _01625_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[383:376] <= _01624_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[375:368] <= _01623_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[367:360] <= _01622_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[359:352] <= _01621_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[351:344] <= _01620_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[343:336] <= _01619_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[335:328] <= _01618_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[327:320] <= _01617_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[319:312] <= _01615_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[311:304] <= _01614_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[303:296] <= _01613_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[295:288] <= _01612_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[287:280] <= _01611_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[279:272] <= _01610_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[271:264] <= _01609_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[263:256] <= _01608_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[255:248] <= _01607_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[247:240] <= _01606_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[239:232] <= _01604_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[231:224] <= _01603_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[223:216] <= _01602_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[215:208] <= _01601_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[207:200] <= _01600_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[199:192] <= _01599_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[191:184] <= _01598_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[183:176] <= _01597_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[175:168] <= _01596_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[167:160] <= _01595_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[159:152] <= _01593_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[151:144] <= _01592_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[143:136] <= _01591_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[135:128] <= _01590_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[127:120] <= _01589_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[119:112] <= _01588_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[111:104] <= _01587_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[103:96] <= _01586_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[95:88] <= _01705_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[87:80] <= _01694_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[79:72] <= _01682_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[71:64] <= _01671_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[63:56] <= _01660_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[55:48] <= _01649_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[47:40] <= _01638_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[39:32] <= _01627_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[31:24] <= _01616_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[23:16] <= _01605_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[15:8] <= _01594_;
  always @(posedge nvdla_core_clk)
      wt1_sd_data[7:0] <= _01683_;
  always @(posedge nvdla_core_clk)
      wt1_sd_nan <= _01713_;
  always @(posedge nvdla_core_clk)
      wt1_sd_exp <= _01711_;
  always @(posedge nvdla_core_clk)
      wt1_sd_mask <= _01712_;
  always @(posedge nvdla_core_clk)
      wt1_sd_nz <= _01714_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt1_sd_pvld <= 1'b0;
    else
      wt1_sd_pvld <= wt1_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[1023:1016] <= _01323_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[1015:1008] <= _01322_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[1007:1000] <= _01321_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[999:992] <= _01448_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[991:984] <= _01447_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[983:976] <= _01446_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[975:968] <= _01445_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[967:960] <= _01444_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[959:952] <= _01442_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[951:944] <= _01441_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[943:936] <= _01440_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[935:928] <= _01439_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[927:920] <= _01438_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[919:912] <= _01437_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[911:904] <= _01436_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[903:896] <= _01435_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[895:888] <= _01434_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[887:880] <= _01433_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[879:872] <= _01431_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[871:864] <= _01430_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[863:856] <= _01429_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[855:848] <= _01428_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[847:840] <= _01427_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[839:832] <= _01426_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[831:824] <= _01425_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[823:816] <= _01424_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[815:808] <= _01423_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[807:800] <= _01422_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[799:792] <= _01419_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[791:784] <= _01418_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[783:776] <= _01417_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[775:768] <= _01416_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[767:760] <= _01415_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[759:752] <= _01414_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[751:744] <= _01413_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[743:736] <= _01412_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[735:728] <= _01411_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[727:720] <= _01410_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[719:712] <= _01408_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[711:704] <= _01407_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[703:696] <= _01406_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[695:688] <= _01405_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[687:680] <= _01404_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[679:672] <= _01403_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[671:664] <= _01402_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[663:656] <= _01401_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[655:648] <= _01400_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[647:640] <= _01399_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[639:632] <= _01397_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[631:624] <= _01396_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[623:616] <= _01395_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[615:608] <= _01394_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[607:600] <= _01393_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[599:592] <= _01392_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[591:584] <= _01391_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[583:576] <= _01390_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[575:568] <= _01389_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[567:560] <= _01388_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[559:552] <= _01386_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[551:544] <= _01385_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[543:536] <= _01384_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[535:528] <= _01383_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[527:520] <= _01382_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[519:512] <= _01381_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[511:504] <= _01380_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[503:496] <= _01379_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[495:488] <= _01378_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[487:480] <= _01377_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[479:472] <= _01375_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[471:464] <= _01374_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[463:456] <= _01373_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[455:448] <= _01372_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[447:440] <= _01371_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[439:432] <= _01370_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[431:424] <= _01369_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[423:416] <= _01368_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[415:408] <= _01367_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[407:400] <= _01366_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[399:392] <= _01364_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[391:384] <= _01363_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[383:376] <= _01362_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[375:368] <= _01361_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[367:360] <= _01360_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[359:352] <= _01359_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[351:344] <= _01358_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[343:336] <= _01357_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[335:328] <= _01356_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[327:320] <= _01355_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[319:312] <= _01353_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[311:304] <= _01352_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[303:296] <= _01351_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[295:288] <= _01350_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[287:280] <= _01349_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[279:272] <= _01348_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[271:264] <= _01347_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[263:256] <= _01346_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[255:248] <= _01345_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[247:240] <= _01344_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[239:232] <= _01342_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[231:224] <= _01341_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[223:216] <= _01340_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[215:208] <= _01339_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[207:200] <= _01338_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[199:192] <= _01337_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[191:184] <= _01336_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[183:176] <= _01335_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[175:168] <= _01334_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[167:160] <= _01333_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[159:152] <= _01331_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[151:144] <= _01330_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[143:136] <= _01329_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[135:128] <= _01328_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[127:120] <= _01327_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[119:112] <= _01326_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[111:104] <= _01325_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[103:96] <= _01324_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[95:88] <= _01443_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[87:80] <= _01432_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[79:72] <= _01420_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[71:64] <= _01409_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[63:56] <= _01398_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[55:48] <= _01387_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[47:40] <= _01376_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[39:32] <= _01365_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[31:24] <= _01354_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[23:16] <= _01343_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[15:8] <= _01332_;
  always @(posedge nvdla_core_clk)
      wt0_sd_data[7:0] <= _01421_;
  always @(posedge nvdla_core_clk)
      wt0_sd_nan <= _01451_;
  always @(posedge nvdla_core_clk)
      wt0_sd_exp <= _01449_;
  always @(posedge nvdla_core_clk)
      wt0_sd_mask <= _01450_;
  always @(posedge nvdla_core_clk)
      wt0_sd_nz <= _01452_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt0_sd_pvld <= 1'b0;
    else
      wt0_sd_pvld <= wt0_sd_pvld_w;
  always @(posedge nvdla_core_clk)
      wt_pre_data[1023:1016] <= _03289_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[1015:1008] <= _03288_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[1007:1000] <= _03287_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[999:992] <= _03414_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[991:984] <= _03413_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[983:976] <= _03412_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[975:968] <= _03411_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[967:960] <= _03410_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[959:952] <= _03408_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[951:944] <= _03407_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[943:936] <= _03406_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[935:928] <= _03405_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[927:920] <= _03404_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[919:912] <= _03403_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[911:904] <= _03402_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[903:896] <= _03401_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[895:888] <= _03400_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[887:880] <= _03399_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[879:872] <= _03397_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[871:864] <= _03396_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[863:856] <= _03395_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[855:848] <= _03394_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[847:840] <= _03393_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[839:832] <= _03392_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[831:824] <= _03391_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[823:816] <= _03390_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[815:808] <= _03389_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[807:800] <= _03388_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[799:792] <= _03385_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[791:784] <= _03384_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[783:776] <= _03383_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[775:768] <= _03382_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[767:760] <= _03381_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[759:752] <= _03380_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[751:744] <= _03379_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[743:736] <= _03378_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[735:728] <= _03377_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[727:720] <= _03376_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[719:712] <= _03374_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[711:704] <= _03373_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[703:696] <= _03372_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[695:688] <= _03371_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[687:680] <= _03370_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[679:672] <= _03369_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[671:664] <= _03368_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[663:656] <= _03367_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[655:648] <= _03366_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[647:640] <= _03365_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[639:632] <= _03363_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[631:624] <= _03362_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[623:616] <= _03361_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[615:608] <= _03360_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[607:600] <= _03359_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[599:592] <= _03358_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[591:584] <= _03357_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[583:576] <= _03356_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[575:568] <= _03355_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[567:560] <= _03354_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[559:552] <= _03352_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[551:544] <= _03351_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[543:536] <= _03350_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[535:528] <= _03349_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[527:520] <= _03348_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[519:512] <= _03347_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[511:504] <= _03346_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[503:496] <= _03345_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[495:488] <= _03344_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[487:480] <= _03343_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[479:472] <= _03341_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[471:464] <= _03340_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[463:456] <= _03339_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[455:448] <= _03338_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[447:440] <= _03337_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[439:432] <= _03336_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[431:424] <= _03335_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[423:416] <= _03334_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[415:408] <= _03333_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[407:400] <= _03332_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[399:392] <= _03330_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[391:384] <= _03329_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[383:376] <= _03328_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[375:368] <= _03327_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[367:360] <= _03326_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[359:352] <= _03325_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[351:344] <= _03324_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[343:336] <= _03323_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[335:328] <= _03322_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[327:320] <= _03321_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[319:312] <= _03319_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[311:304] <= _03318_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[303:296] <= _03317_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[295:288] <= _03316_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[287:280] <= _03315_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[279:272] <= _03314_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[271:264] <= _03313_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[263:256] <= _03312_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[255:248] <= _03311_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[247:240] <= _03310_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[239:232] <= _03308_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[231:224] <= _03307_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[223:216] <= _03306_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[215:208] <= _03305_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[207:200] <= _03304_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[199:192] <= _03303_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[191:184] <= _03302_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[183:176] <= _03301_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[175:168] <= _03300_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[167:160] <= _03299_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[159:152] <= _03297_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[151:144] <= _03296_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[143:136] <= _03295_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[135:128] <= _03294_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[127:120] <= _03293_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[119:112] <= _03292_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[111:104] <= _03291_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[103:96] <= _03290_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[95:88] <= _03409_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[87:80] <= _03398_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[79:72] <= _03386_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[71:64] <= _03375_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[63:56] <= _03364_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[55:48] <= _03353_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[47:40] <= _03342_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[39:32] <= _03331_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[31:24] <= _03320_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[23:16] <= _03309_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[15:8] <= _03298_;
  always @(posedge nvdla_core_clk)
      wt_pre_data[7:0] <= _03387_;
  always @(posedge nvdla_core_clk)
      wt_pre_nan <= _03417_;
  always @(posedge nvdla_core_clk)
      wt_pre_exp <= _03415_;
  always @(posedge nvdla_core_clk)
      wt_pre_mask <= _03416_;
  always @(posedge nvdla_core_clk)
      wt_pre_nz <= _03418_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wt_pre_sel <= 8'b00000000;
    else
      wt_pre_sel <= in_wt_sel;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_is_int16_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      cfg_is_int16_d1 <= _00001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_is_fp16_d1 <= 98'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      cfg_is_fp16_d1 <= _00000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_is_int8_d1 <= 65'b00000000000000000000000000000000000000000000000000000000000000000;
    else
      cfg_is_int8_d1 <= _00002_;
  assign _00901_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41093" *) dat_pre_data[1023:1016] : dat_actv_data_reg7[1023:1016];
  assign _00900_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41083" *) dat_pre_data[1015:1008] : dat_actv_data_reg7[1015:1008];
  assign _00899_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41073" *) dat_pre_data[1007:1000] : dat_actv_data_reg7[1007:1000];
  assign _01026_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41063" *) dat_pre_data[999:992] : dat_actv_data_reg7[999:992];
  assign _01025_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41053" *) dat_pre_data[991:984] : dat_actv_data_reg7[991:984];
  assign _01024_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41043" *) dat_pre_data[983:976] : dat_actv_data_reg7[983:976];
  assign _01023_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41033" *) dat_pre_data[975:968] : dat_actv_data_reg7[975:968];
  assign _01022_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41023" *) dat_pre_data[967:960] : dat_actv_data_reg7[967:960];
  assign _01020_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41013" *) dat_pre_data[959:952] : dat_actv_data_reg7[959:952];
  assign _01019_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:41003" *) dat_pre_data[951:944] : dat_actv_data_reg7[951:944];
  assign _01018_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40993" *) dat_pre_data[943:936] : dat_actv_data_reg7[943:936];
  assign _01017_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40983" *) dat_pre_data[935:928] : dat_actv_data_reg7[935:928];
  assign _01016_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40973" *) dat_pre_data[927:920] : dat_actv_data_reg7[927:920];
  assign _01015_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40963" *) dat_pre_data[919:912] : dat_actv_data_reg7[919:912];
  assign _01014_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40953" *) dat_pre_data[911:904] : dat_actv_data_reg7[911:904];
  assign _01013_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40943" *) dat_pre_data[903:896] : dat_actv_data_reg7[903:896];
  assign _01012_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40933" *) dat_pre_data[895:888] : dat_actv_data_reg7[895:888];
  assign _01011_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40923" *) dat_pre_data[887:880] : dat_actv_data_reg7[887:880];
  assign _01009_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40913" *) dat_pre_data[879:872] : dat_actv_data_reg7[879:872];
  assign _01008_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40903" *) dat_pre_data[871:864] : dat_actv_data_reg7[871:864];
  assign _01007_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40893" *) dat_pre_data[863:856] : dat_actv_data_reg7[863:856];
  assign _01006_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40883" *) dat_pre_data[855:848] : dat_actv_data_reg7[855:848];
  assign _01005_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40873" *) dat_pre_data[847:840] : dat_actv_data_reg7[847:840];
  assign _01004_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40863" *) dat_pre_data[839:832] : dat_actv_data_reg7[839:832];
  assign _01003_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40853" *) dat_pre_data[831:824] : dat_actv_data_reg7[831:824];
  assign _01002_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40843" *) dat_pre_data[823:816] : dat_actv_data_reg7[823:816];
  assign _01001_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40833" *) dat_pre_data[815:808] : dat_actv_data_reg7[815:808];
  assign _01000_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40823" *) dat_pre_data[807:800] : dat_actv_data_reg7[807:800];
  assign _00997_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40813" *) dat_pre_data[799:792] : dat_actv_data_reg7[799:792];
  assign _00996_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40803" *) dat_pre_data[791:784] : dat_actv_data_reg7[791:784];
  assign _00995_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40793" *) dat_pre_data[783:776] : dat_actv_data_reg7[783:776];
  assign _00994_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40783" *) dat_pre_data[775:768] : dat_actv_data_reg7[775:768];
  assign _00993_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40773" *) dat_pre_data[767:760] : dat_actv_data_reg7[767:760];
  assign _00992_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40763" *) dat_pre_data[759:752] : dat_actv_data_reg7[759:752];
  assign _00991_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40753" *) dat_pre_data[751:744] : dat_actv_data_reg7[751:744];
  assign _00990_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40743" *) dat_pre_data[743:736] : dat_actv_data_reg7[743:736];
  assign _00989_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40733" *) dat_pre_data[735:728] : dat_actv_data_reg7[735:728];
  assign _00988_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40723" *) dat_pre_data[727:720] : dat_actv_data_reg7[727:720];
  assign _00986_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40713" *) dat_pre_data[719:712] : dat_actv_data_reg7[719:712];
  assign _00985_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40703" *) dat_pre_data[711:704] : dat_actv_data_reg7[711:704];
  assign _00984_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40693" *) dat_pre_data[703:696] : dat_actv_data_reg7[703:696];
  assign _00983_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40683" *) dat_pre_data[695:688] : dat_actv_data_reg7[695:688];
  assign _00982_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40673" *) dat_pre_data[687:680] : dat_actv_data_reg7[687:680];
  assign _00981_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40663" *) dat_pre_data[679:672] : dat_actv_data_reg7[679:672];
  assign _00980_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40653" *) dat_pre_data[671:664] : dat_actv_data_reg7[671:664];
  assign _00979_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40643" *) dat_pre_data[663:656] : dat_actv_data_reg7[663:656];
  assign _00978_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40633" *) dat_pre_data[655:648] : dat_actv_data_reg7[655:648];
  assign _00977_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40623" *) dat_pre_data[647:640] : dat_actv_data_reg7[647:640];
  assign _00975_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40613" *) dat_pre_data[639:632] : dat_actv_data_reg7[639:632];
  assign _00974_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40603" *) dat_pre_data[631:624] : dat_actv_data_reg7[631:624];
  assign _00973_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40593" *) dat_pre_data[623:616] : dat_actv_data_reg7[623:616];
  assign _00972_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40583" *) dat_pre_data[615:608] : dat_actv_data_reg7[615:608];
  assign _00971_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40573" *) dat_pre_data[607:600] : dat_actv_data_reg7[607:600];
  assign _00970_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40563" *) dat_pre_data[599:592] : dat_actv_data_reg7[599:592];
  assign _00969_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40553" *) dat_pre_data[591:584] : dat_actv_data_reg7[591:584];
  assign _00968_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40543" *) dat_pre_data[583:576] : dat_actv_data_reg7[583:576];
  assign _00967_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40533" *) dat_pre_data[575:568] : dat_actv_data_reg7[575:568];
  assign _00966_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40523" *) dat_pre_data[567:560] : dat_actv_data_reg7[567:560];
  assign _00964_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40513" *) dat_pre_data[559:552] : dat_actv_data_reg7[559:552];
  assign _00963_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40503" *) dat_pre_data[551:544] : dat_actv_data_reg7[551:544];
  assign _00962_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40493" *) dat_pre_data[543:536] : dat_actv_data_reg7[543:536];
  assign _00961_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40483" *) dat_pre_data[535:528] : dat_actv_data_reg7[535:528];
  assign _00960_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40473" *) dat_pre_data[527:520] : dat_actv_data_reg7[527:520];
  assign _00959_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40463" *) dat_pre_data[519:512] : dat_actv_data_reg7[519:512];
  assign _00958_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40453" *) dat_pre_data[511:504] : dat_actv_data_reg7[511:504];
  assign _00957_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40443" *) dat_pre_data[503:496] : dat_actv_data_reg7[503:496];
  assign _00956_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40433" *) dat_pre_data[495:488] : dat_actv_data_reg7[495:488];
  assign _00955_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40423" *) dat_pre_data[487:480] : dat_actv_data_reg7[487:480];
  assign _00953_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40413" *) dat_pre_data[479:472] : dat_actv_data_reg7[479:472];
  assign _00952_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40403" *) dat_pre_data[471:464] : dat_actv_data_reg7[471:464];
  assign _00951_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40393" *) dat_pre_data[463:456] : dat_actv_data_reg7[463:456];
  assign _00950_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40383" *) dat_pre_data[455:448] : dat_actv_data_reg7[455:448];
  assign _00949_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40373" *) dat_pre_data[447:440] : dat_actv_data_reg7[447:440];
  assign _00948_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40363" *) dat_pre_data[439:432] : dat_actv_data_reg7[439:432];
  assign _00947_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40353" *) dat_pre_data[431:424] : dat_actv_data_reg7[431:424];
  assign _00946_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40343" *) dat_pre_data[423:416] : dat_actv_data_reg7[423:416];
  assign _00945_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40333" *) dat_pre_data[415:408] : dat_actv_data_reg7[415:408];
  assign _00944_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40323" *) dat_pre_data[407:400] : dat_actv_data_reg7[407:400];
  assign _00942_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40313" *) dat_pre_data[399:392] : dat_actv_data_reg7[399:392];
  assign _00941_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40303" *) dat_pre_data[391:384] : dat_actv_data_reg7[391:384];
  assign _00940_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40293" *) dat_pre_data[383:376] : dat_actv_data_reg7[383:376];
  assign _00939_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40283" *) dat_pre_data[375:368] : dat_actv_data_reg7[375:368];
  assign _00938_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40273" *) dat_pre_data[367:360] : dat_actv_data_reg7[367:360];
  assign _00937_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40263" *) dat_pre_data[359:352] : dat_actv_data_reg7[359:352];
  assign _00936_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40253" *) dat_pre_data[351:344] : dat_actv_data_reg7[351:344];
  assign _00935_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40243" *) dat_pre_data[343:336] : dat_actv_data_reg7[343:336];
  assign _00934_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40233" *) dat_pre_data[335:328] : dat_actv_data_reg7[335:328];
  assign _00933_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40223" *) dat_pre_data[327:320] : dat_actv_data_reg7[327:320];
  assign _00931_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40213" *) dat_pre_data[319:312] : dat_actv_data_reg7[319:312];
  assign _00930_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40203" *) dat_pre_data[311:304] : dat_actv_data_reg7[311:304];
  assign _00929_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40193" *) dat_pre_data[303:296] : dat_actv_data_reg7[303:296];
  assign _00928_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40183" *) dat_pre_data[295:288] : dat_actv_data_reg7[295:288];
  assign _00927_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40173" *) dat_pre_data[287:280] : dat_actv_data_reg7[287:280];
  assign _00926_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40163" *) dat_pre_data[279:272] : dat_actv_data_reg7[279:272];
  assign _00925_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40153" *) dat_pre_data[271:264] : dat_actv_data_reg7[271:264];
  assign _00924_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40143" *) dat_pre_data[263:256] : dat_actv_data_reg7[263:256];
  assign _00923_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40133" *) dat_pre_data[255:248] : dat_actv_data_reg7[255:248];
  assign _00922_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40123" *) dat_pre_data[247:240] : dat_actv_data_reg7[247:240];
  assign _00920_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40113" *) dat_pre_data[239:232] : dat_actv_data_reg7[239:232];
  assign _00919_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40103" *) dat_pre_data[231:224] : dat_actv_data_reg7[231:224];
  assign _00918_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40093" *) dat_pre_data[223:216] : dat_actv_data_reg7[223:216];
  assign _00917_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40083" *) dat_pre_data[215:208] : dat_actv_data_reg7[215:208];
  assign _00916_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40073" *) dat_pre_data[207:200] : dat_actv_data_reg7[207:200];
  assign _00915_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40063" *) dat_pre_data[199:192] : dat_actv_data_reg7[199:192];
  assign _00914_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40053" *) dat_pre_data[191:184] : dat_actv_data_reg7[191:184];
  assign _00913_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40043" *) dat_pre_data[183:176] : dat_actv_data_reg7[183:176];
  assign _00912_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40033" *) dat_pre_data[175:168] : dat_actv_data_reg7[175:168];
  assign _00911_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40023" *) dat_pre_data[167:160] : dat_actv_data_reg7[167:160];
  assign _00909_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40013" *) dat_pre_data[159:152] : dat_actv_data_reg7[159:152];
  assign _00908_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:40003" *) dat_pre_data[151:144] : dat_actv_data_reg7[151:144];
  assign _00907_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39993" *) dat_pre_data[143:136] : dat_actv_data_reg7[143:136];
  assign _00906_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39983" *) dat_pre_data[135:128] : dat_actv_data_reg7[135:128];
  assign _00905_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39973" *) dat_pre_data[127:120] : dat_actv_data_reg7[127:120];
  assign _00904_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39963" *) dat_pre_data[119:112] : dat_actv_data_reg7[119:112];
  assign _00903_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39953" *) dat_pre_data[111:104] : dat_actv_data_reg7[111:104];
  assign _00902_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39943" *) dat_pre_data[103:96] : dat_actv_data_reg7[103:96];
  assign _01021_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39933" *) dat_pre_data[95:88] : dat_actv_data_reg7[95:88];
  assign _01010_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39923" *) dat_pre_data[87:80] : dat_actv_data_reg7[87:80];
  assign _00998_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39913" *) dat_pre_data[79:72] : dat_actv_data_reg7[79:72];
  assign _00987_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39903" *) dat_pre_data[71:64] : dat_actv_data_reg7[71:64];
  assign _00976_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39893" *) dat_pre_data[63:56] : dat_actv_data_reg7[63:56];
  assign _00965_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39883" *) dat_pre_data[55:48] : dat_actv_data_reg7[55:48];
  assign _00954_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39873" *) dat_pre_data[47:40] : dat_actv_data_reg7[47:40];
  assign _00943_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39863" *) dat_pre_data[39:32] : dat_actv_data_reg7[39:32];
  assign _00932_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39853" *) dat_pre_data[31:24] : dat_actv_data_reg7[31:24];
  assign _00921_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39843" *) dat_pre_data[23:16] : dat_actv_data_reg7[23:16];
  assign _00910_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39833" *) dat_pre_data[15:8] : dat_actv_data_reg7[15:8];
  assign _00999_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39823" *) dat_pre_data[7:0] : dat_actv_data_reg7[7:0];
  assign _01034_ = _05699_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39813" *) dat_pre_nan : dat_actv_nan_reg7;
  assign _01042_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39803" *) dat_pre_nz : dat_actv_nz_reg7;
  assign _00773_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39786" *) dat_pre_data[1023:1016] : dat_actv_data_reg6[1023:1016];
  assign _00772_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39776" *) dat_pre_data[1015:1008] : dat_actv_data_reg6[1015:1008];
  assign _00771_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39766" *) dat_pre_data[1007:1000] : dat_actv_data_reg6[1007:1000];
  assign _00898_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39756" *) dat_pre_data[999:992] : dat_actv_data_reg6[999:992];
  assign _00897_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39746" *) dat_pre_data[991:984] : dat_actv_data_reg6[991:984];
  assign _00896_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39736" *) dat_pre_data[983:976] : dat_actv_data_reg6[983:976];
  assign _00895_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39726" *) dat_pre_data[975:968] : dat_actv_data_reg6[975:968];
  assign _00894_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39716" *) dat_pre_data[967:960] : dat_actv_data_reg6[967:960];
  assign _00892_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39706" *) dat_pre_data[959:952] : dat_actv_data_reg6[959:952];
  assign _00891_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39696" *) dat_pre_data[951:944] : dat_actv_data_reg6[951:944];
  assign _00890_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39686" *) dat_pre_data[943:936] : dat_actv_data_reg6[943:936];
  assign _00889_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39676" *) dat_pre_data[935:928] : dat_actv_data_reg6[935:928];
  assign _00888_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39666" *) dat_pre_data[927:920] : dat_actv_data_reg6[927:920];
  assign _00887_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39656" *) dat_pre_data[919:912] : dat_actv_data_reg6[919:912];
  assign _00886_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39646" *) dat_pre_data[911:904] : dat_actv_data_reg6[911:904];
  assign _00885_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39636" *) dat_pre_data[903:896] : dat_actv_data_reg6[903:896];
  assign _00884_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39626" *) dat_pre_data[895:888] : dat_actv_data_reg6[895:888];
  assign _00883_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39616" *) dat_pre_data[887:880] : dat_actv_data_reg6[887:880];
  assign _00881_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39606" *) dat_pre_data[879:872] : dat_actv_data_reg6[879:872];
  assign _00880_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39596" *) dat_pre_data[871:864] : dat_actv_data_reg6[871:864];
  assign _00879_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39586" *) dat_pre_data[863:856] : dat_actv_data_reg6[863:856];
  assign _00878_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39576" *) dat_pre_data[855:848] : dat_actv_data_reg6[855:848];
  assign _00877_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39566" *) dat_pre_data[847:840] : dat_actv_data_reg6[847:840];
  assign _00876_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39556" *) dat_pre_data[839:832] : dat_actv_data_reg6[839:832];
  assign _00875_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39546" *) dat_pre_data[831:824] : dat_actv_data_reg6[831:824];
  assign _00874_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39536" *) dat_pre_data[823:816] : dat_actv_data_reg6[823:816];
  assign _00873_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39526" *) dat_pre_data[815:808] : dat_actv_data_reg6[815:808];
  assign _00872_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39516" *) dat_pre_data[807:800] : dat_actv_data_reg6[807:800];
  assign _00869_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39506" *) dat_pre_data[799:792] : dat_actv_data_reg6[799:792];
  assign _00868_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39496" *) dat_pre_data[791:784] : dat_actv_data_reg6[791:784];
  assign _00867_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39486" *) dat_pre_data[783:776] : dat_actv_data_reg6[783:776];
  assign _00866_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39476" *) dat_pre_data[775:768] : dat_actv_data_reg6[775:768];
  assign _00865_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39466" *) dat_pre_data[767:760] : dat_actv_data_reg6[767:760];
  assign _00864_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39456" *) dat_pre_data[759:752] : dat_actv_data_reg6[759:752];
  assign _00863_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39446" *) dat_pre_data[751:744] : dat_actv_data_reg6[751:744];
  assign _00862_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39436" *) dat_pre_data[743:736] : dat_actv_data_reg6[743:736];
  assign _00861_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39426" *) dat_pre_data[735:728] : dat_actv_data_reg6[735:728];
  assign _00860_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39416" *) dat_pre_data[727:720] : dat_actv_data_reg6[727:720];
  assign _00858_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39406" *) dat_pre_data[719:712] : dat_actv_data_reg6[719:712];
  assign _00857_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39396" *) dat_pre_data[711:704] : dat_actv_data_reg6[711:704];
  assign _00856_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39386" *) dat_pre_data[703:696] : dat_actv_data_reg6[703:696];
  assign _00855_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39376" *) dat_pre_data[695:688] : dat_actv_data_reg6[695:688];
  assign _00854_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39366" *) dat_pre_data[687:680] : dat_actv_data_reg6[687:680];
  assign _00853_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39356" *) dat_pre_data[679:672] : dat_actv_data_reg6[679:672];
  assign _00852_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39346" *) dat_pre_data[671:664] : dat_actv_data_reg6[671:664];
  assign _00851_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39336" *) dat_pre_data[663:656] : dat_actv_data_reg6[663:656];
  assign _00850_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39326" *) dat_pre_data[655:648] : dat_actv_data_reg6[655:648];
  assign _00849_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39316" *) dat_pre_data[647:640] : dat_actv_data_reg6[647:640];
  assign _00847_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39306" *) dat_pre_data[639:632] : dat_actv_data_reg6[639:632];
  assign _00846_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39296" *) dat_pre_data[631:624] : dat_actv_data_reg6[631:624];
  assign _00845_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39286" *) dat_pre_data[623:616] : dat_actv_data_reg6[623:616];
  assign _00844_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39276" *) dat_pre_data[615:608] : dat_actv_data_reg6[615:608];
  assign _00843_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39266" *) dat_pre_data[607:600] : dat_actv_data_reg6[607:600];
  assign _00842_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39256" *) dat_pre_data[599:592] : dat_actv_data_reg6[599:592];
  assign _00841_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39246" *) dat_pre_data[591:584] : dat_actv_data_reg6[591:584];
  assign _00840_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39236" *) dat_pre_data[583:576] : dat_actv_data_reg6[583:576];
  assign _00839_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39226" *) dat_pre_data[575:568] : dat_actv_data_reg6[575:568];
  assign _00838_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39216" *) dat_pre_data[567:560] : dat_actv_data_reg6[567:560];
  assign _00836_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39206" *) dat_pre_data[559:552] : dat_actv_data_reg6[559:552];
  assign _00835_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39196" *) dat_pre_data[551:544] : dat_actv_data_reg6[551:544];
  assign _00834_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39186" *) dat_pre_data[543:536] : dat_actv_data_reg6[543:536];
  assign _00833_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39176" *) dat_pre_data[535:528] : dat_actv_data_reg6[535:528];
  assign _00832_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39166" *) dat_pre_data[527:520] : dat_actv_data_reg6[527:520];
  assign _00831_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39156" *) dat_pre_data[519:512] : dat_actv_data_reg6[519:512];
  assign _00830_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39146" *) dat_pre_data[511:504] : dat_actv_data_reg6[511:504];
  assign _00829_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39136" *) dat_pre_data[503:496] : dat_actv_data_reg6[503:496];
  assign _00828_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39126" *) dat_pre_data[495:488] : dat_actv_data_reg6[495:488];
  assign _00827_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39116" *) dat_pre_data[487:480] : dat_actv_data_reg6[487:480];
  assign _00825_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39106" *) dat_pre_data[479:472] : dat_actv_data_reg6[479:472];
  assign _00824_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39096" *) dat_pre_data[471:464] : dat_actv_data_reg6[471:464];
  assign _00823_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39086" *) dat_pre_data[463:456] : dat_actv_data_reg6[463:456];
  assign _00822_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39076" *) dat_pre_data[455:448] : dat_actv_data_reg6[455:448];
  assign _00821_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39066" *) dat_pre_data[447:440] : dat_actv_data_reg6[447:440];
  assign _00820_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39056" *) dat_pre_data[439:432] : dat_actv_data_reg6[439:432];
  assign _00819_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39046" *) dat_pre_data[431:424] : dat_actv_data_reg6[431:424];
  assign _00818_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39036" *) dat_pre_data[423:416] : dat_actv_data_reg6[423:416];
  assign _00817_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39026" *) dat_pre_data[415:408] : dat_actv_data_reg6[415:408];
  assign _00816_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39016" *) dat_pre_data[407:400] : dat_actv_data_reg6[407:400];
  assign _00814_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:39006" *) dat_pre_data[399:392] : dat_actv_data_reg6[399:392];
  assign _00813_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38996" *) dat_pre_data[391:384] : dat_actv_data_reg6[391:384];
  assign _00812_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38986" *) dat_pre_data[383:376] : dat_actv_data_reg6[383:376];
  assign _00811_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38976" *) dat_pre_data[375:368] : dat_actv_data_reg6[375:368];
  assign _00810_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38966" *) dat_pre_data[367:360] : dat_actv_data_reg6[367:360];
  assign _00809_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38956" *) dat_pre_data[359:352] : dat_actv_data_reg6[359:352];
  assign _00808_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38946" *) dat_pre_data[351:344] : dat_actv_data_reg6[351:344];
  assign _00807_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38936" *) dat_pre_data[343:336] : dat_actv_data_reg6[343:336];
  assign _00806_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38926" *) dat_pre_data[335:328] : dat_actv_data_reg6[335:328];
  assign _00805_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38916" *) dat_pre_data[327:320] : dat_actv_data_reg6[327:320];
  assign _00803_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38906" *) dat_pre_data[319:312] : dat_actv_data_reg6[319:312];
  assign _00802_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38896" *) dat_pre_data[311:304] : dat_actv_data_reg6[311:304];
  assign _00801_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38886" *) dat_pre_data[303:296] : dat_actv_data_reg6[303:296];
  assign _00800_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38876" *) dat_pre_data[295:288] : dat_actv_data_reg6[295:288];
  assign _00799_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38866" *) dat_pre_data[287:280] : dat_actv_data_reg6[287:280];
  assign _00798_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38856" *) dat_pre_data[279:272] : dat_actv_data_reg6[279:272];
  assign _00797_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38846" *) dat_pre_data[271:264] : dat_actv_data_reg6[271:264];
  assign _00796_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38836" *) dat_pre_data[263:256] : dat_actv_data_reg6[263:256];
  assign _00795_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38826" *) dat_pre_data[255:248] : dat_actv_data_reg6[255:248];
  assign _00794_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38816" *) dat_pre_data[247:240] : dat_actv_data_reg6[247:240];
  assign _00792_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38806" *) dat_pre_data[239:232] : dat_actv_data_reg6[239:232];
  assign _00791_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38796" *) dat_pre_data[231:224] : dat_actv_data_reg6[231:224];
  assign _00790_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38786" *) dat_pre_data[223:216] : dat_actv_data_reg6[223:216];
  assign _00789_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38776" *) dat_pre_data[215:208] : dat_actv_data_reg6[215:208];
  assign _00788_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38766" *) dat_pre_data[207:200] : dat_actv_data_reg6[207:200];
  assign _00787_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38756" *) dat_pre_data[199:192] : dat_actv_data_reg6[199:192];
  assign _00786_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38746" *) dat_pre_data[191:184] : dat_actv_data_reg6[191:184];
  assign _00785_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38736" *) dat_pre_data[183:176] : dat_actv_data_reg6[183:176];
  assign _00784_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38726" *) dat_pre_data[175:168] : dat_actv_data_reg6[175:168];
  assign _00783_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38716" *) dat_pre_data[167:160] : dat_actv_data_reg6[167:160];
  assign _00781_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38706" *) dat_pre_data[159:152] : dat_actv_data_reg6[159:152];
  assign _00780_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38696" *) dat_pre_data[151:144] : dat_actv_data_reg6[151:144];
  assign _00779_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38686" *) dat_pre_data[143:136] : dat_actv_data_reg6[143:136];
  assign _00778_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38676" *) dat_pre_data[135:128] : dat_actv_data_reg6[135:128];
  assign _00777_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38666" *) dat_pre_data[127:120] : dat_actv_data_reg6[127:120];
  assign _00776_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38656" *) dat_pre_data[119:112] : dat_actv_data_reg6[119:112];
  assign _00775_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38646" *) dat_pre_data[111:104] : dat_actv_data_reg6[111:104];
  assign _00774_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38636" *) dat_pre_data[103:96] : dat_actv_data_reg6[103:96];
  assign _00893_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38626" *) dat_pre_data[95:88] : dat_actv_data_reg6[95:88];
  assign _00882_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38616" *) dat_pre_data[87:80] : dat_actv_data_reg6[87:80];
  assign _00870_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38606" *) dat_pre_data[79:72] : dat_actv_data_reg6[79:72];
  assign _00859_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38596" *) dat_pre_data[71:64] : dat_actv_data_reg6[71:64];
  assign _00848_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38586" *) dat_pre_data[63:56] : dat_actv_data_reg6[63:56];
  assign _00837_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38576" *) dat_pre_data[55:48] : dat_actv_data_reg6[55:48];
  assign _00826_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38566" *) dat_pre_data[47:40] : dat_actv_data_reg6[47:40];
  assign _00815_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38556" *) dat_pre_data[39:32] : dat_actv_data_reg6[39:32];
  assign _00804_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38546" *) dat_pre_data[31:24] : dat_actv_data_reg6[31:24];
  assign _00793_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38536" *) dat_pre_data[23:16] : dat_actv_data_reg6[23:16];
  assign _00782_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38526" *) dat_pre_data[15:8] : dat_actv_data_reg6[15:8];
  assign _00871_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38516" *) dat_pre_data[7:0] : dat_actv_data_reg6[7:0];
  assign _01033_ = _05697_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38506" *) dat_pre_nan : dat_actv_nan_reg6;
  assign _01041_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38496" *) dat_pre_nz : dat_actv_nz_reg6;
  assign _00645_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38479" *) dat_pre_data[1023:1016] : dat_actv_data_reg5[1023:1016];
  assign _00644_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38469" *) dat_pre_data[1015:1008] : dat_actv_data_reg5[1015:1008];
  assign _00643_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38459" *) dat_pre_data[1007:1000] : dat_actv_data_reg5[1007:1000];
  assign _00770_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38449" *) dat_pre_data[999:992] : dat_actv_data_reg5[999:992];
  assign _00769_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38439" *) dat_pre_data[991:984] : dat_actv_data_reg5[991:984];
  assign _00768_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38429" *) dat_pre_data[983:976] : dat_actv_data_reg5[983:976];
  assign _00767_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38419" *) dat_pre_data[975:968] : dat_actv_data_reg5[975:968];
  assign _00766_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38409" *) dat_pre_data[967:960] : dat_actv_data_reg5[967:960];
  assign _00764_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38399" *) dat_pre_data[959:952] : dat_actv_data_reg5[959:952];
  assign _00763_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38389" *) dat_pre_data[951:944] : dat_actv_data_reg5[951:944];
  assign _00762_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38379" *) dat_pre_data[943:936] : dat_actv_data_reg5[943:936];
  assign _00761_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38369" *) dat_pre_data[935:928] : dat_actv_data_reg5[935:928];
  assign _00760_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38359" *) dat_pre_data[927:920] : dat_actv_data_reg5[927:920];
  assign _00759_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38349" *) dat_pre_data[919:912] : dat_actv_data_reg5[919:912];
  assign _00758_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38339" *) dat_pre_data[911:904] : dat_actv_data_reg5[911:904];
  assign _00757_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38329" *) dat_pre_data[903:896] : dat_actv_data_reg5[903:896];
  assign _00756_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38319" *) dat_pre_data[895:888] : dat_actv_data_reg5[895:888];
  assign _00755_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38309" *) dat_pre_data[887:880] : dat_actv_data_reg5[887:880];
  assign _00753_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38299" *) dat_pre_data[879:872] : dat_actv_data_reg5[879:872];
  assign _00752_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38289" *) dat_pre_data[871:864] : dat_actv_data_reg5[871:864];
  assign _00751_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38279" *) dat_pre_data[863:856] : dat_actv_data_reg5[863:856];
  assign _00750_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38269" *) dat_pre_data[855:848] : dat_actv_data_reg5[855:848];
  assign _00749_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38259" *) dat_pre_data[847:840] : dat_actv_data_reg5[847:840];
  assign _00748_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38249" *) dat_pre_data[839:832] : dat_actv_data_reg5[839:832];
  assign _00747_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38239" *) dat_pre_data[831:824] : dat_actv_data_reg5[831:824];
  assign _00746_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38229" *) dat_pre_data[823:816] : dat_actv_data_reg5[823:816];
  assign _00745_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38219" *) dat_pre_data[815:808] : dat_actv_data_reg5[815:808];
  assign _00744_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38209" *) dat_pre_data[807:800] : dat_actv_data_reg5[807:800];
  assign _00741_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38199" *) dat_pre_data[799:792] : dat_actv_data_reg5[799:792];
  assign _00740_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38189" *) dat_pre_data[791:784] : dat_actv_data_reg5[791:784];
  assign _00739_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38179" *) dat_pre_data[783:776] : dat_actv_data_reg5[783:776];
  assign _00738_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38169" *) dat_pre_data[775:768] : dat_actv_data_reg5[775:768];
  assign _00737_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38159" *) dat_pre_data[767:760] : dat_actv_data_reg5[767:760];
  assign _00736_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38149" *) dat_pre_data[759:752] : dat_actv_data_reg5[759:752];
  assign _00735_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38139" *) dat_pre_data[751:744] : dat_actv_data_reg5[751:744];
  assign _00734_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38129" *) dat_pre_data[743:736] : dat_actv_data_reg5[743:736];
  assign _00733_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38119" *) dat_pre_data[735:728] : dat_actv_data_reg5[735:728];
  assign _00732_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38109" *) dat_pre_data[727:720] : dat_actv_data_reg5[727:720];
  assign _00730_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38099" *) dat_pre_data[719:712] : dat_actv_data_reg5[719:712];
  assign _00729_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38089" *) dat_pre_data[711:704] : dat_actv_data_reg5[711:704];
  assign _00728_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38079" *) dat_pre_data[703:696] : dat_actv_data_reg5[703:696];
  assign _00727_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38069" *) dat_pre_data[695:688] : dat_actv_data_reg5[695:688];
  assign _00726_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38059" *) dat_pre_data[687:680] : dat_actv_data_reg5[687:680];
  assign _00725_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38049" *) dat_pre_data[679:672] : dat_actv_data_reg5[679:672];
  assign _00724_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38039" *) dat_pre_data[671:664] : dat_actv_data_reg5[671:664];
  assign _00723_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38029" *) dat_pre_data[663:656] : dat_actv_data_reg5[663:656];
  assign _00722_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38019" *) dat_pre_data[655:648] : dat_actv_data_reg5[655:648];
  assign _00721_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:38009" *) dat_pre_data[647:640] : dat_actv_data_reg5[647:640];
  assign _00719_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37999" *) dat_pre_data[639:632] : dat_actv_data_reg5[639:632];
  assign _00718_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37989" *) dat_pre_data[631:624] : dat_actv_data_reg5[631:624];
  assign _00717_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37979" *) dat_pre_data[623:616] : dat_actv_data_reg5[623:616];
  assign _00716_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37969" *) dat_pre_data[615:608] : dat_actv_data_reg5[615:608];
  assign _00715_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37959" *) dat_pre_data[607:600] : dat_actv_data_reg5[607:600];
  assign _00714_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37949" *) dat_pre_data[599:592] : dat_actv_data_reg5[599:592];
  assign _00713_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37939" *) dat_pre_data[591:584] : dat_actv_data_reg5[591:584];
  assign _00712_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37929" *) dat_pre_data[583:576] : dat_actv_data_reg5[583:576];
  assign _00711_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37919" *) dat_pre_data[575:568] : dat_actv_data_reg5[575:568];
  assign _00710_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37909" *) dat_pre_data[567:560] : dat_actv_data_reg5[567:560];
  assign _00708_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37899" *) dat_pre_data[559:552] : dat_actv_data_reg5[559:552];
  assign _00707_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37889" *) dat_pre_data[551:544] : dat_actv_data_reg5[551:544];
  assign _00706_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37879" *) dat_pre_data[543:536] : dat_actv_data_reg5[543:536];
  assign _00705_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37869" *) dat_pre_data[535:528] : dat_actv_data_reg5[535:528];
  assign _00704_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37859" *) dat_pre_data[527:520] : dat_actv_data_reg5[527:520];
  assign _00703_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37849" *) dat_pre_data[519:512] : dat_actv_data_reg5[519:512];
  assign _00702_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37839" *) dat_pre_data[511:504] : dat_actv_data_reg5[511:504];
  assign _00701_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37829" *) dat_pre_data[503:496] : dat_actv_data_reg5[503:496];
  assign _00700_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37819" *) dat_pre_data[495:488] : dat_actv_data_reg5[495:488];
  assign _00699_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37809" *) dat_pre_data[487:480] : dat_actv_data_reg5[487:480];
  assign _00697_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37799" *) dat_pre_data[479:472] : dat_actv_data_reg5[479:472];
  assign _00696_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37789" *) dat_pre_data[471:464] : dat_actv_data_reg5[471:464];
  assign _00695_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37779" *) dat_pre_data[463:456] : dat_actv_data_reg5[463:456];
  assign _00694_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37769" *) dat_pre_data[455:448] : dat_actv_data_reg5[455:448];
  assign _00693_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37759" *) dat_pre_data[447:440] : dat_actv_data_reg5[447:440];
  assign _00692_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37749" *) dat_pre_data[439:432] : dat_actv_data_reg5[439:432];
  assign _00691_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37739" *) dat_pre_data[431:424] : dat_actv_data_reg5[431:424];
  assign _00690_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37729" *) dat_pre_data[423:416] : dat_actv_data_reg5[423:416];
  assign _00689_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37719" *) dat_pre_data[415:408] : dat_actv_data_reg5[415:408];
  assign _00688_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37709" *) dat_pre_data[407:400] : dat_actv_data_reg5[407:400];
  assign _00686_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37699" *) dat_pre_data[399:392] : dat_actv_data_reg5[399:392];
  assign _00685_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37689" *) dat_pre_data[391:384] : dat_actv_data_reg5[391:384];
  assign _00684_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37679" *) dat_pre_data[383:376] : dat_actv_data_reg5[383:376];
  assign _00683_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37669" *) dat_pre_data[375:368] : dat_actv_data_reg5[375:368];
  assign _00682_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37659" *) dat_pre_data[367:360] : dat_actv_data_reg5[367:360];
  assign _00681_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37649" *) dat_pre_data[359:352] : dat_actv_data_reg5[359:352];
  assign _00680_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37639" *) dat_pre_data[351:344] : dat_actv_data_reg5[351:344];
  assign _00679_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37629" *) dat_pre_data[343:336] : dat_actv_data_reg5[343:336];
  assign _00678_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37619" *) dat_pre_data[335:328] : dat_actv_data_reg5[335:328];
  assign _00677_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37609" *) dat_pre_data[327:320] : dat_actv_data_reg5[327:320];
  assign _00675_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37599" *) dat_pre_data[319:312] : dat_actv_data_reg5[319:312];
  assign _00674_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37589" *) dat_pre_data[311:304] : dat_actv_data_reg5[311:304];
  assign _00673_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37579" *) dat_pre_data[303:296] : dat_actv_data_reg5[303:296];
  assign _00672_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37569" *) dat_pre_data[295:288] : dat_actv_data_reg5[295:288];
  assign _00671_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37559" *) dat_pre_data[287:280] : dat_actv_data_reg5[287:280];
  assign _00670_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37549" *) dat_pre_data[279:272] : dat_actv_data_reg5[279:272];
  assign _00669_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37539" *) dat_pre_data[271:264] : dat_actv_data_reg5[271:264];
  assign _00668_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37529" *) dat_pre_data[263:256] : dat_actv_data_reg5[263:256];
  assign _00667_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37519" *) dat_pre_data[255:248] : dat_actv_data_reg5[255:248];
  assign _00666_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37509" *) dat_pre_data[247:240] : dat_actv_data_reg5[247:240];
  assign _00664_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37499" *) dat_pre_data[239:232] : dat_actv_data_reg5[239:232];
  assign _00663_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37489" *) dat_pre_data[231:224] : dat_actv_data_reg5[231:224];
  assign _00662_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37479" *) dat_pre_data[223:216] : dat_actv_data_reg5[223:216];
  assign _00661_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37469" *) dat_pre_data[215:208] : dat_actv_data_reg5[215:208];
  assign _00660_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37459" *) dat_pre_data[207:200] : dat_actv_data_reg5[207:200];
  assign _00659_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37449" *) dat_pre_data[199:192] : dat_actv_data_reg5[199:192];
  assign _00658_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37439" *) dat_pre_data[191:184] : dat_actv_data_reg5[191:184];
  assign _00657_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37429" *) dat_pre_data[183:176] : dat_actv_data_reg5[183:176];
  assign _00656_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37419" *) dat_pre_data[175:168] : dat_actv_data_reg5[175:168];
  assign _00655_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37409" *) dat_pre_data[167:160] : dat_actv_data_reg5[167:160];
  assign _00653_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37399" *) dat_pre_data[159:152] : dat_actv_data_reg5[159:152];
  assign _00652_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37389" *) dat_pre_data[151:144] : dat_actv_data_reg5[151:144];
  assign _00651_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37379" *) dat_pre_data[143:136] : dat_actv_data_reg5[143:136];
  assign _00650_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37369" *) dat_pre_data[135:128] : dat_actv_data_reg5[135:128];
  assign _00649_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37359" *) dat_pre_data[127:120] : dat_actv_data_reg5[127:120];
  assign _00648_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37349" *) dat_pre_data[119:112] : dat_actv_data_reg5[119:112];
  assign _00647_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37339" *) dat_pre_data[111:104] : dat_actv_data_reg5[111:104];
  assign _00646_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37329" *) dat_pre_data[103:96] : dat_actv_data_reg5[103:96];
  assign _00765_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37319" *) dat_pre_data[95:88] : dat_actv_data_reg5[95:88];
  assign _00754_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37309" *) dat_pre_data[87:80] : dat_actv_data_reg5[87:80];
  assign _00742_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37299" *) dat_pre_data[79:72] : dat_actv_data_reg5[79:72];
  assign _00731_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37289" *) dat_pre_data[71:64] : dat_actv_data_reg5[71:64];
  assign _00720_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37279" *) dat_pre_data[63:56] : dat_actv_data_reg5[63:56];
  assign _00709_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37269" *) dat_pre_data[55:48] : dat_actv_data_reg5[55:48];
  assign _00698_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37259" *) dat_pre_data[47:40] : dat_actv_data_reg5[47:40];
  assign _00687_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37249" *) dat_pre_data[39:32] : dat_actv_data_reg5[39:32];
  assign _00676_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37239" *) dat_pre_data[31:24] : dat_actv_data_reg5[31:24];
  assign _00665_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37229" *) dat_pre_data[23:16] : dat_actv_data_reg5[23:16];
  assign _00654_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37219" *) dat_pre_data[15:8] : dat_actv_data_reg5[15:8];
  assign _00743_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37209" *) dat_pre_data[7:0] : dat_actv_data_reg5[7:0];
  assign _01032_ = _05696_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37199" *) dat_pre_nan : dat_actv_nan_reg5;
  assign _01040_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37189" *) dat_pre_nz : dat_actv_nz_reg5;
  assign _00517_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37172" *) dat_pre_data[1023:1016] : dat_actv_data_reg4[1023:1016];
  assign _00516_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37162" *) dat_pre_data[1015:1008] : dat_actv_data_reg4[1015:1008];
  assign _00515_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37152" *) dat_pre_data[1007:1000] : dat_actv_data_reg4[1007:1000];
  assign _00642_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37142" *) dat_pre_data[999:992] : dat_actv_data_reg4[999:992];
  assign _00641_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37132" *) dat_pre_data[991:984] : dat_actv_data_reg4[991:984];
  assign _00640_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37122" *) dat_pre_data[983:976] : dat_actv_data_reg4[983:976];
  assign _00639_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37112" *) dat_pre_data[975:968] : dat_actv_data_reg4[975:968];
  assign _00638_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37102" *) dat_pre_data[967:960] : dat_actv_data_reg4[967:960];
  assign _00636_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37092" *) dat_pre_data[959:952] : dat_actv_data_reg4[959:952];
  assign _00635_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37082" *) dat_pre_data[951:944] : dat_actv_data_reg4[951:944];
  assign _00634_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37072" *) dat_pre_data[943:936] : dat_actv_data_reg4[943:936];
  assign _00633_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37062" *) dat_pre_data[935:928] : dat_actv_data_reg4[935:928];
  assign _00632_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37052" *) dat_pre_data[927:920] : dat_actv_data_reg4[927:920];
  assign _00631_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37042" *) dat_pre_data[919:912] : dat_actv_data_reg4[919:912];
  assign _00630_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37032" *) dat_pre_data[911:904] : dat_actv_data_reg4[911:904];
  assign _00629_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37022" *) dat_pre_data[903:896] : dat_actv_data_reg4[903:896];
  assign _00628_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37012" *) dat_pre_data[895:888] : dat_actv_data_reg4[895:888];
  assign _00627_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:37002" *) dat_pre_data[887:880] : dat_actv_data_reg4[887:880];
  assign _00625_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36992" *) dat_pre_data[879:872] : dat_actv_data_reg4[879:872];
  assign _00624_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36982" *) dat_pre_data[871:864] : dat_actv_data_reg4[871:864];
  assign _00623_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36972" *) dat_pre_data[863:856] : dat_actv_data_reg4[863:856];
  assign _00622_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36962" *) dat_pre_data[855:848] : dat_actv_data_reg4[855:848];
  assign _00621_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36952" *) dat_pre_data[847:840] : dat_actv_data_reg4[847:840];
  assign _00620_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36942" *) dat_pre_data[839:832] : dat_actv_data_reg4[839:832];
  assign _00619_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36932" *) dat_pre_data[831:824] : dat_actv_data_reg4[831:824];
  assign _00618_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36922" *) dat_pre_data[823:816] : dat_actv_data_reg4[823:816];
  assign _00617_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36912" *) dat_pre_data[815:808] : dat_actv_data_reg4[815:808];
  assign _00616_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36902" *) dat_pre_data[807:800] : dat_actv_data_reg4[807:800];
  assign _00613_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36892" *) dat_pre_data[799:792] : dat_actv_data_reg4[799:792];
  assign _00612_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36882" *) dat_pre_data[791:784] : dat_actv_data_reg4[791:784];
  assign _00611_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36872" *) dat_pre_data[783:776] : dat_actv_data_reg4[783:776];
  assign _00610_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36862" *) dat_pre_data[775:768] : dat_actv_data_reg4[775:768];
  assign _00609_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36852" *) dat_pre_data[767:760] : dat_actv_data_reg4[767:760];
  assign _00608_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36842" *) dat_pre_data[759:752] : dat_actv_data_reg4[759:752];
  assign _00607_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36832" *) dat_pre_data[751:744] : dat_actv_data_reg4[751:744];
  assign _00606_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36822" *) dat_pre_data[743:736] : dat_actv_data_reg4[743:736];
  assign _00605_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36812" *) dat_pre_data[735:728] : dat_actv_data_reg4[735:728];
  assign _00604_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36802" *) dat_pre_data[727:720] : dat_actv_data_reg4[727:720];
  assign _00602_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36792" *) dat_pre_data[719:712] : dat_actv_data_reg4[719:712];
  assign _00601_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36782" *) dat_pre_data[711:704] : dat_actv_data_reg4[711:704];
  assign _00600_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36772" *) dat_pre_data[703:696] : dat_actv_data_reg4[703:696];
  assign _00599_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36762" *) dat_pre_data[695:688] : dat_actv_data_reg4[695:688];
  assign _00598_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36752" *) dat_pre_data[687:680] : dat_actv_data_reg4[687:680];
  assign _00597_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36742" *) dat_pre_data[679:672] : dat_actv_data_reg4[679:672];
  assign _00596_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36732" *) dat_pre_data[671:664] : dat_actv_data_reg4[671:664];
  assign _00595_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36722" *) dat_pre_data[663:656] : dat_actv_data_reg4[663:656];
  assign _00594_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36712" *) dat_pre_data[655:648] : dat_actv_data_reg4[655:648];
  assign _00593_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36702" *) dat_pre_data[647:640] : dat_actv_data_reg4[647:640];
  assign _00591_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36692" *) dat_pre_data[639:632] : dat_actv_data_reg4[639:632];
  assign _00590_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36682" *) dat_pre_data[631:624] : dat_actv_data_reg4[631:624];
  assign _00589_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36672" *) dat_pre_data[623:616] : dat_actv_data_reg4[623:616];
  assign _00588_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36662" *) dat_pre_data[615:608] : dat_actv_data_reg4[615:608];
  assign _00587_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36652" *) dat_pre_data[607:600] : dat_actv_data_reg4[607:600];
  assign _00586_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36642" *) dat_pre_data[599:592] : dat_actv_data_reg4[599:592];
  assign _00585_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36632" *) dat_pre_data[591:584] : dat_actv_data_reg4[591:584];
  assign _00584_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36622" *) dat_pre_data[583:576] : dat_actv_data_reg4[583:576];
  assign _00583_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36612" *) dat_pre_data[575:568] : dat_actv_data_reg4[575:568];
  assign _00582_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36602" *) dat_pre_data[567:560] : dat_actv_data_reg4[567:560];
  assign _00580_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36592" *) dat_pre_data[559:552] : dat_actv_data_reg4[559:552];
  assign _00579_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36582" *) dat_pre_data[551:544] : dat_actv_data_reg4[551:544];
  assign _00578_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36572" *) dat_pre_data[543:536] : dat_actv_data_reg4[543:536];
  assign _00577_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36562" *) dat_pre_data[535:528] : dat_actv_data_reg4[535:528];
  assign _00576_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36552" *) dat_pre_data[527:520] : dat_actv_data_reg4[527:520];
  assign _00575_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36542" *) dat_pre_data[519:512] : dat_actv_data_reg4[519:512];
  assign _00574_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36532" *) dat_pre_data[511:504] : dat_actv_data_reg4[511:504];
  assign _00573_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36522" *) dat_pre_data[503:496] : dat_actv_data_reg4[503:496];
  assign _00572_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36512" *) dat_pre_data[495:488] : dat_actv_data_reg4[495:488];
  assign _00571_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36502" *) dat_pre_data[487:480] : dat_actv_data_reg4[487:480];
  assign _00569_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36492" *) dat_pre_data[479:472] : dat_actv_data_reg4[479:472];
  assign _00568_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36482" *) dat_pre_data[471:464] : dat_actv_data_reg4[471:464];
  assign _00567_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36472" *) dat_pre_data[463:456] : dat_actv_data_reg4[463:456];
  assign _00566_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36462" *) dat_pre_data[455:448] : dat_actv_data_reg4[455:448];
  assign _00565_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36452" *) dat_pre_data[447:440] : dat_actv_data_reg4[447:440];
  assign _00564_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36442" *) dat_pre_data[439:432] : dat_actv_data_reg4[439:432];
  assign _00563_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36432" *) dat_pre_data[431:424] : dat_actv_data_reg4[431:424];
  assign _00562_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36422" *) dat_pre_data[423:416] : dat_actv_data_reg4[423:416];
  assign _00561_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36412" *) dat_pre_data[415:408] : dat_actv_data_reg4[415:408];
  assign _00560_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36402" *) dat_pre_data[407:400] : dat_actv_data_reg4[407:400];
  assign _00558_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36392" *) dat_pre_data[399:392] : dat_actv_data_reg4[399:392];
  assign _00557_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36382" *) dat_pre_data[391:384] : dat_actv_data_reg4[391:384];
  assign _00556_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36372" *) dat_pre_data[383:376] : dat_actv_data_reg4[383:376];
  assign _00555_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36362" *) dat_pre_data[375:368] : dat_actv_data_reg4[375:368];
  assign _00554_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36352" *) dat_pre_data[367:360] : dat_actv_data_reg4[367:360];
  assign _00553_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36342" *) dat_pre_data[359:352] : dat_actv_data_reg4[359:352];
  assign _00552_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36332" *) dat_pre_data[351:344] : dat_actv_data_reg4[351:344];
  assign _00551_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36322" *) dat_pre_data[343:336] : dat_actv_data_reg4[343:336];
  assign _00550_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36312" *) dat_pre_data[335:328] : dat_actv_data_reg4[335:328];
  assign _00549_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36302" *) dat_pre_data[327:320] : dat_actv_data_reg4[327:320];
  assign _00547_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36292" *) dat_pre_data[319:312] : dat_actv_data_reg4[319:312];
  assign _00546_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36282" *) dat_pre_data[311:304] : dat_actv_data_reg4[311:304];
  assign _00545_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36272" *) dat_pre_data[303:296] : dat_actv_data_reg4[303:296];
  assign _00544_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36262" *) dat_pre_data[295:288] : dat_actv_data_reg4[295:288];
  assign _00543_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36252" *) dat_pre_data[287:280] : dat_actv_data_reg4[287:280];
  assign _00542_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36242" *) dat_pre_data[279:272] : dat_actv_data_reg4[279:272];
  assign _00541_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36232" *) dat_pre_data[271:264] : dat_actv_data_reg4[271:264];
  assign _00540_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36222" *) dat_pre_data[263:256] : dat_actv_data_reg4[263:256];
  assign _00539_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36212" *) dat_pre_data[255:248] : dat_actv_data_reg4[255:248];
  assign _00538_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36202" *) dat_pre_data[247:240] : dat_actv_data_reg4[247:240];
  assign _00536_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36192" *) dat_pre_data[239:232] : dat_actv_data_reg4[239:232];
  assign _00535_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36182" *) dat_pre_data[231:224] : dat_actv_data_reg4[231:224];
  assign _00534_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36172" *) dat_pre_data[223:216] : dat_actv_data_reg4[223:216];
  assign _00533_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36162" *) dat_pre_data[215:208] : dat_actv_data_reg4[215:208];
  assign _00532_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36152" *) dat_pre_data[207:200] : dat_actv_data_reg4[207:200];
  assign _00531_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36142" *) dat_pre_data[199:192] : dat_actv_data_reg4[199:192];
  assign _00530_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36132" *) dat_pre_data[191:184] : dat_actv_data_reg4[191:184];
  assign _00529_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36122" *) dat_pre_data[183:176] : dat_actv_data_reg4[183:176];
  assign _00528_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36112" *) dat_pre_data[175:168] : dat_actv_data_reg4[175:168];
  assign _00527_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36102" *) dat_pre_data[167:160] : dat_actv_data_reg4[167:160];
  assign _00525_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36092" *) dat_pre_data[159:152] : dat_actv_data_reg4[159:152];
  assign _00524_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36082" *) dat_pre_data[151:144] : dat_actv_data_reg4[151:144];
  assign _00523_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36072" *) dat_pre_data[143:136] : dat_actv_data_reg4[143:136];
  assign _00522_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36062" *) dat_pre_data[135:128] : dat_actv_data_reg4[135:128];
  assign _00521_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36052" *) dat_pre_data[127:120] : dat_actv_data_reg4[127:120];
  assign _00520_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36042" *) dat_pre_data[119:112] : dat_actv_data_reg4[119:112];
  assign _00519_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36032" *) dat_pre_data[111:104] : dat_actv_data_reg4[111:104];
  assign _00518_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36022" *) dat_pre_data[103:96] : dat_actv_data_reg4[103:96];
  assign _00637_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36012" *) dat_pre_data[95:88] : dat_actv_data_reg4[95:88];
  assign _00626_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:36002" *) dat_pre_data[87:80] : dat_actv_data_reg4[87:80];
  assign _00614_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35992" *) dat_pre_data[79:72] : dat_actv_data_reg4[79:72];
  assign _00603_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35982" *) dat_pre_data[71:64] : dat_actv_data_reg4[71:64];
  assign _00592_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35972" *) dat_pre_data[63:56] : dat_actv_data_reg4[63:56];
  assign _00581_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35962" *) dat_pre_data[55:48] : dat_actv_data_reg4[55:48];
  assign _00570_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35952" *) dat_pre_data[47:40] : dat_actv_data_reg4[47:40];
  assign _00559_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35942" *) dat_pre_data[39:32] : dat_actv_data_reg4[39:32];
  assign _00548_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35932" *) dat_pre_data[31:24] : dat_actv_data_reg4[31:24];
  assign _00537_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35922" *) dat_pre_data[23:16] : dat_actv_data_reg4[23:16];
  assign _00526_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35912" *) dat_pre_data[15:8] : dat_actv_data_reg4[15:8];
  assign _00615_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35902" *) dat_pre_data[7:0] : dat_actv_data_reg4[7:0];
  assign _01031_ = _05695_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35892" *) dat_pre_nan : dat_actv_nan_reg4;
  assign _01039_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35882" *) dat_pre_nz : dat_actv_nz_reg4;
  assign _00389_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35865" *) dat_pre_data[1023:1016] : dat_actv_data_reg3[1023:1016];
  assign _00388_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35855" *) dat_pre_data[1015:1008] : dat_actv_data_reg3[1015:1008];
  assign _00387_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35845" *) dat_pre_data[1007:1000] : dat_actv_data_reg3[1007:1000];
  assign _00514_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35835" *) dat_pre_data[999:992] : dat_actv_data_reg3[999:992];
  assign _00513_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35825" *) dat_pre_data[991:984] : dat_actv_data_reg3[991:984];
  assign _00512_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35815" *) dat_pre_data[983:976] : dat_actv_data_reg3[983:976];
  assign _00511_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35805" *) dat_pre_data[975:968] : dat_actv_data_reg3[975:968];
  assign _00510_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35795" *) dat_pre_data[967:960] : dat_actv_data_reg3[967:960];
  assign _00508_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35785" *) dat_pre_data[959:952] : dat_actv_data_reg3[959:952];
  assign _00507_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35775" *) dat_pre_data[951:944] : dat_actv_data_reg3[951:944];
  assign _00506_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35765" *) dat_pre_data[943:936] : dat_actv_data_reg3[943:936];
  assign _00505_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35755" *) dat_pre_data[935:928] : dat_actv_data_reg3[935:928];
  assign _00504_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35745" *) dat_pre_data[927:920] : dat_actv_data_reg3[927:920];
  assign _00503_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35735" *) dat_pre_data[919:912] : dat_actv_data_reg3[919:912];
  assign _00502_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35725" *) dat_pre_data[911:904] : dat_actv_data_reg3[911:904];
  assign _00501_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35715" *) dat_pre_data[903:896] : dat_actv_data_reg3[903:896];
  assign _00500_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35705" *) dat_pre_data[895:888] : dat_actv_data_reg3[895:888];
  assign _00499_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35695" *) dat_pre_data[887:880] : dat_actv_data_reg3[887:880];
  assign _00497_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35685" *) dat_pre_data[879:872] : dat_actv_data_reg3[879:872];
  assign _00496_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35675" *) dat_pre_data[871:864] : dat_actv_data_reg3[871:864];
  assign _00495_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35665" *) dat_pre_data[863:856] : dat_actv_data_reg3[863:856];
  assign _00494_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35655" *) dat_pre_data[855:848] : dat_actv_data_reg3[855:848];
  assign _00493_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35645" *) dat_pre_data[847:840] : dat_actv_data_reg3[847:840];
  assign _00492_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35635" *) dat_pre_data[839:832] : dat_actv_data_reg3[839:832];
  assign _00491_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35625" *) dat_pre_data[831:824] : dat_actv_data_reg3[831:824];
  assign _00490_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35615" *) dat_pre_data[823:816] : dat_actv_data_reg3[823:816];
  assign _00489_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35605" *) dat_pre_data[815:808] : dat_actv_data_reg3[815:808];
  assign _00488_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35595" *) dat_pre_data[807:800] : dat_actv_data_reg3[807:800];
  assign _00485_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35585" *) dat_pre_data[799:792] : dat_actv_data_reg3[799:792];
  assign _00484_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35575" *) dat_pre_data[791:784] : dat_actv_data_reg3[791:784];
  assign _00483_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35565" *) dat_pre_data[783:776] : dat_actv_data_reg3[783:776];
  assign _00482_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35555" *) dat_pre_data[775:768] : dat_actv_data_reg3[775:768];
  assign _00481_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35545" *) dat_pre_data[767:760] : dat_actv_data_reg3[767:760];
  assign _00480_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35535" *) dat_pre_data[759:752] : dat_actv_data_reg3[759:752];
  assign _00479_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35525" *) dat_pre_data[751:744] : dat_actv_data_reg3[751:744];
  assign _00478_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35515" *) dat_pre_data[743:736] : dat_actv_data_reg3[743:736];
  assign _00477_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35505" *) dat_pre_data[735:728] : dat_actv_data_reg3[735:728];
  assign _00476_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35495" *) dat_pre_data[727:720] : dat_actv_data_reg3[727:720];
  assign _00474_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35485" *) dat_pre_data[719:712] : dat_actv_data_reg3[719:712];
  assign _00473_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35475" *) dat_pre_data[711:704] : dat_actv_data_reg3[711:704];
  assign _00472_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35465" *) dat_pre_data[703:696] : dat_actv_data_reg3[703:696];
  assign _00471_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35455" *) dat_pre_data[695:688] : dat_actv_data_reg3[695:688];
  assign _00470_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35445" *) dat_pre_data[687:680] : dat_actv_data_reg3[687:680];
  assign _00469_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35435" *) dat_pre_data[679:672] : dat_actv_data_reg3[679:672];
  assign _00468_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35425" *) dat_pre_data[671:664] : dat_actv_data_reg3[671:664];
  assign _00467_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35415" *) dat_pre_data[663:656] : dat_actv_data_reg3[663:656];
  assign _00466_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35405" *) dat_pre_data[655:648] : dat_actv_data_reg3[655:648];
  assign _00465_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35395" *) dat_pre_data[647:640] : dat_actv_data_reg3[647:640];
  assign _00463_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35385" *) dat_pre_data[639:632] : dat_actv_data_reg3[639:632];
  assign _00462_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35375" *) dat_pre_data[631:624] : dat_actv_data_reg3[631:624];
  assign _00461_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35365" *) dat_pre_data[623:616] : dat_actv_data_reg3[623:616];
  assign _00460_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35355" *) dat_pre_data[615:608] : dat_actv_data_reg3[615:608];
  assign _00459_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35345" *) dat_pre_data[607:600] : dat_actv_data_reg3[607:600];
  assign _00458_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35335" *) dat_pre_data[599:592] : dat_actv_data_reg3[599:592];
  assign _00457_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35325" *) dat_pre_data[591:584] : dat_actv_data_reg3[591:584];
  assign _00456_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35315" *) dat_pre_data[583:576] : dat_actv_data_reg3[583:576];
  assign _00455_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35305" *) dat_pre_data[575:568] : dat_actv_data_reg3[575:568];
  assign _00454_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35295" *) dat_pre_data[567:560] : dat_actv_data_reg3[567:560];
  assign _00452_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35285" *) dat_pre_data[559:552] : dat_actv_data_reg3[559:552];
  assign _00451_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35275" *) dat_pre_data[551:544] : dat_actv_data_reg3[551:544];
  assign _00450_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35265" *) dat_pre_data[543:536] : dat_actv_data_reg3[543:536];
  assign _00449_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35255" *) dat_pre_data[535:528] : dat_actv_data_reg3[535:528];
  assign _00448_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35245" *) dat_pre_data[527:520] : dat_actv_data_reg3[527:520];
  assign _00447_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35235" *) dat_pre_data[519:512] : dat_actv_data_reg3[519:512];
  assign _00446_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35225" *) dat_pre_data[511:504] : dat_actv_data_reg3[511:504];
  assign _00445_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35215" *) dat_pre_data[503:496] : dat_actv_data_reg3[503:496];
  assign _00444_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35205" *) dat_pre_data[495:488] : dat_actv_data_reg3[495:488];
  assign _00443_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35195" *) dat_pre_data[487:480] : dat_actv_data_reg3[487:480];
  assign _00441_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35185" *) dat_pre_data[479:472] : dat_actv_data_reg3[479:472];
  assign _00440_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35175" *) dat_pre_data[471:464] : dat_actv_data_reg3[471:464];
  assign _00439_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35165" *) dat_pre_data[463:456] : dat_actv_data_reg3[463:456];
  assign _00438_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35155" *) dat_pre_data[455:448] : dat_actv_data_reg3[455:448];
  assign _00437_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35145" *) dat_pre_data[447:440] : dat_actv_data_reg3[447:440];
  assign _00436_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35135" *) dat_pre_data[439:432] : dat_actv_data_reg3[439:432];
  assign _00435_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35125" *) dat_pre_data[431:424] : dat_actv_data_reg3[431:424];
  assign _00434_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35115" *) dat_pre_data[423:416] : dat_actv_data_reg3[423:416];
  assign _00433_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35105" *) dat_pre_data[415:408] : dat_actv_data_reg3[415:408];
  assign _00432_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35095" *) dat_pre_data[407:400] : dat_actv_data_reg3[407:400];
  assign _00430_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35085" *) dat_pre_data[399:392] : dat_actv_data_reg3[399:392];
  assign _00429_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35075" *) dat_pre_data[391:384] : dat_actv_data_reg3[391:384];
  assign _00428_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35065" *) dat_pre_data[383:376] : dat_actv_data_reg3[383:376];
  assign _00427_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35055" *) dat_pre_data[375:368] : dat_actv_data_reg3[375:368];
  assign _00426_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35045" *) dat_pre_data[367:360] : dat_actv_data_reg3[367:360];
  assign _00425_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35035" *) dat_pre_data[359:352] : dat_actv_data_reg3[359:352];
  assign _00424_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35025" *) dat_pre_data[351:344] : dat_actv_data_reg3[351:344];
  assign _00423_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35015" *) dat_pre_data[343:336] : dat_actv_data_reg3[343:336];
  assign _00422_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:35005" *) dat_pre_data[335:328] : dat_actv_data_reg3[335:328];
  assign _00421_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34995" *) dat_pre_data[327:320] : dat_actv_data_reg3[327:320];
  assign _00419_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34985" *) dat_pre_data[319:312] : dat_actv_data_reg3[319:312];
  assign _00418_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34975" *) dat_pre_data[311:304] : dat_actv_data_reg3[311:304];
  assign _00417_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34965" *) dat_pre_data[303:296] : dat_actv_data_reg3[303:296];
  assign _00416_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34955" *) dat_pre_data[295:288] : dat_actv_data_reg3[295:288];
  assign _00415_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34945" *) dat_pre_data[287:280] : dat_actv_data_reg3[287:280];
  assign _00414_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34935" *) dat_pre_data[279:272] : dat_actv_data_reg3[279:272];
  assign _00413_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34925" *) dat_pre_data[271:264] : dat_actv_data_reg3[271:264];
  assign _00412_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34915" *) dat_pre_data[263:256] : dat_actv_data_reg3[263:256];
  assign _00411_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34905" *) dat_pre_data[255:248] : dat_actv_data_reg3[255:248];
  assign _00410_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34895" *) dat_pre_data[247:240] : dat_actv_data_reg3[247:240];
  assign _00408_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34885" *) dat_pre_data[239:232] : dat_actv_data_reg3[239:232];
  assign _00407_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34875" *) dat_pre_data[231:224] : dat_actv_data_reg3[231:224];
  assign _00406_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34865" *) dat_pre_data[223:216] : dat_actv_data_reg3[223:216];
  assign _00405_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34855" *) dat_pre_data[215:208] : dat_actv_data_reg3[215:208];
  assign _00404_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34845" *) dat_pre_data[207:200] : dat_actv_data_reg3[207:200];
  assign _00403_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34835" *) dat_pre_data[199:192] : dat_actv_data_reg3[199:192];
  assign _00402_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34825" *) dat_pre_data[191:184] : dat_actv_data_reg3[191:184];
  assign _00401_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34815" *) dat_pre_data[183:176] : dat_actv_data_reg3[183:176];
  assign _00400_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34805" *) dat_pre_data[175:168] : dat_actv_data_reg3[175:168];
  assign _00399_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34795" *) dat_pre_data[167:160] : dat_actv_data_reg3[167:160];
  assign _00397_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34785" *) dat_pre_data[159:152] : dat_actv_data_reg3[159:152];
  assign _00396_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34775" *) dat_pre_data[151:144] : dat_actv_data_reg3[151:144];
  assign _00395_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34765" *) dat_pre_data[143:136] : dat_actv_data_reg3[143:136];
  assign _00394_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34755" *) dat_pre_data[135:128] : dat_actv_data_reg3[135:128];
  assign _00393_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34745" *) dat_pre_data[127:120] : dat_actv_data_reg3[127:120];
  assign _00392_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34735" *) dat_pre_data[119:112] : dat_actv_data_reg3[119:112];
  assign _00391_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34725" *) dat_pre_data[111:104] : dat_actv_data_reg3[111:104];
  assign _00390_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34715" *) dat_pre_data[103:96] : dat_actv_data_reg3[103:96];
  assign _00509_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34705" *) dat_pre_data[95:88] : dat_actv_data_reg3[95:88];
  assign _00498_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34695" *) dat_pre_data[87:80] : dat_actv_data_reg3[87:80];
  assign _00486_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34685" *) dat_pre_data[79:72] : dat_actv_data_reg3[79:72];
  assign _00475_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34675" *) dat_pre_data[71:64] : dat_actv_data_reg3[71:64];
  assign _00464_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34665" *) dat_pre_data[63:56] : dat_actv_data_reg3[63:56];
  assign _00453_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34655" *) dat_pre_data[55:48] : dat_actv_data_reg3[55:48];
  assign _00442_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34645" *) dat_pre_data[47:40] : dat_actv_data_reg3[47:40];
  assign _00431_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34635" *) dat_pre_data[39:32] : dat_actv_data_reg3[39:32];
  assign _00420_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34625" *) dat_pre_data[31:24] : dat_actv_data_reg3[31:24];
  assign _00409_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34615" *) dat_pre_data[23:16] : dat_actv_data_reg3[23:16];
  assign _00398_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34605" *) dat_pre_data[15:8] : dat_actv_data_reg3[15:8];
  assign _00487_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34595" *) dat_pre_data[7:0] : dat_actv_data_reg3[7:0];
  assign _01030_ = _05694_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34585" *) dat_pre_nan : dat_actv_nan_reg3;
  assign _01038_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34575" *) dat_pre_nz : dat_actv_nz_reg3;
  assign _00261_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34558" *) dat_pre_data[1023:1016] : dat_actv_data_reg2[1023:1016];
  assign _00260_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34548" *) dat_pre_data[1015:1008] : dat_actv_data_reg2[1015:1008];
  assign _00259_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34538" *) dat_pre_data[1007:1000] : dat_actv_data_reg2[1007:1000];
  assign _00386_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34528" *) dat_pre_data[999:992] : dat_actv_data_reg2[999:992];
  assign _00385_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34518" *) dat_pre_data[991:984] : dat_actv_data_reg2[991:984];
  assign _00384_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34508" *) dat_pre_data[983:976] : dat_actv_data_reg2[983:976];
  assign _00383_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34498" *) dat_pre_data[975:968] : dat_actv_data_reg2[975:968];
  assign _00382_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34488" *) dat_pre_data[967:960] : dat_actv_data_reg2[967:960];
  assign _00380_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34478" *) dat_pre_data[959:952] : dat_actv_data_reg2[959:952];
  assign _00379_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34468" *) dat_pre_data[951:944] : dat_actv_data_reg2[951:944];
  assign _00378_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34458" *) dat_pre_data[943:936] : dat_actv_data_reg2[943:936];
  assign _00377_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34448" *) dat_pre_data[935:928] : dat_actv_data_reg2[935:928];
  assign _00376_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34438" *) dat_pre_data[927:920] : dat_actv_data_reg2[927:920];
  assign _00375_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34428" *) dat_pre_data[919:912] : dat_actv_data_reg2[919:912];
  assign _00374_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34418" *) dat_pre_data[911:904] : dat_actv_data_reg2[911:904];
  assign _00373_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34408" *) dat_pre_data[903:896] : dat_actv_data_reg2[903:896];
  assign _00372_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34398" *) dat_pre_data[895:888] : dat_actv_data_reg2[895:888];
  assign _00371_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34388" *) dat_pre_data[887:880] : dat_actv_data_reg2[887:880];
  assign _00369_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34378" *) dat_pre_data[879:872] : dat_actv_data_reg2[879:872];
  assign _00368_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34368" *) dat_pre_data[871:864] : dat_actv_data_reg2[871:864];
  assign _00367_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34358" *) dat_pre_data[863:856] : dat_actv_data_reg2[863:856];
  assign _00366_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34348" *) dat_pre_data[855:848] : dat_actv_data_reg2[855:848];
  assign _00365_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34338" *) dat_pre_data[847:840] : dat_actv_data_reg2[847:840];
  assign _00364_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34328" *) dat_pre_data[839:832] : dat_actv_data_reg2[839:832];
  assign _00363_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34318" *) dat_pre_data[831:824] : dat_actv_data_reg2[831:824];
  assign _00362_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34308" *) dat_pre_data[823:816] : dat_actv_data_reg2[823:816];
  assign _00361_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34298" *) dat_pre_data[815:808] : dat_actv_data_reg2[815:808];
  assign _00360_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34288" *) dat_pre_data[807:800] : dat_actv_data_reg2[807:800];
  assign _00357_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34278" *) dat_pre_data[799:792] : dat_actv_data_reg2[799:792];
  assign _00356_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34268" *) dat_pre_data[791:784] : dat_actv_data_reg2[791:784];
  assign _00355_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34258" *) dat_pre_data[783:776] : dat_actv_data_reg2[783:776];
  assign _00354_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34248" *) dat_pre_data[775:768] : dat_actv_data_reg2[775:768];
  assign _00353_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34238" *) dat_pre_data[767:760] : dat_actv_data_reg2[767:760];
  assign _00352_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34228" *) dat_pre_data[759:752] : dat_actv_data_reg2[759:752];
  assign _00351_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34218" *) dat_pre_data[751:744] : dat_actv_data_reg2[751:744];
  assign _00350_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34208" *) dat_pre_data[743:736] : dat_actv_data_reg2[743:736];
  assign _00349_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34198" *) dat_pre_data[735:728] : dat_actv_data_reg2[735:728];
  assign _00348_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34188" *) dat_pre_data[727:720] : dat_actv_data_reg2[727:720];
  assign _00346_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34178" *) dat_pre_data[719:712] : dat_actv_data_reg2[719:712];
  assign _00345_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34168" *) dat_pre_data[711:704] : dat_actv_data_reg2[711:704];
  assign _00344_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34158" *) dat_pre_data[703:696] : dat_actv_data_reg2[703:696];
  assign _00343_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34148" *) dat_pre_data[695:688] : dat_actv_data_reg2[695:688];
  assign _00342_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34138" *) dat_pre_data[687:680] : dat_actv_data_reg2[687:680];
  assign _00341_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34128" *) dat_pre_data[679:672] : dat_actv_data_reg2[679:672];
  assign _00340_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34118" *) dat_pre_data[671:664] : dat_actv_data_reg2[671:664];
  assign _00339_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34108" *) dat_pre_data[663:656] : dat_actv_data_reg2[663:656];
  assign _00338_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34098" *) dat_pre_data[655:648] : dat_actv_data_reg2[655:648];
  assign _00337_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34088" *) dat_pre_data[647:640] : dat_actv_data_reg2[647:640];
  assign _00335_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34078" *) dat_pre_data[639:632] : dat_actv_data_reg2[639:632];
  assign _00334_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34068" *) dat_pre_data[631:624] : dat_actv_data_reg2[631:624];
  assign _00333_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34058" *) dat_pre_data[623:616] : dat_actv_data_reg2[623:616];
  assign _00332_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34048" *) dat_pre_data[615:608] : dat_actv_data_reg2[615:608];
  assign _00331_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34038" *) dat_pre_data[607:600] : dat_actv_data_reg2[607:600];
  assign _00330_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34028" *) dat_pre_data[599:592] : dat_actv_data_reg2[599:592];
  assign _00329_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34018" *) dat_pre_data[591:584] : dat_actv_data_reg2[591:584];
  assign _00328_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:34008" *) dat_pre_data[583:576] : dat_actv_data_reg2[583:576];
  assign _00327_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33998" *) dat_pre_data[575:568] : dat_actv_data_reg2[575:568];
  assign _00326_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33988" *) dat_pre_data[567:560] : dat_actv_data_reg2[567:560];
  assign _00324_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33978" *) dat_pre_data[559:552] : dat_actv_data_reg2[559:552];
  assign _00323_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33968" *) dat_pre_data[551:544] : dat_actv_data_reg2[551:544];
  assign _00322_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33958" *) dat_pre_data[543:536] : dat_actv_data_reg2[543:536];
  assign _00321_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33948" *) dat_pre_data[535:528] : dat_actv_data_reg2[535:528];
  assign _00320_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33938" *) dat_pre_data[527:520] : dat_actv_data_reg2[527:520];
  assign _00319_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33928" *) dat_pre_data[519:512] : dat_actv_data_reg2[519:512];
  assign _00318_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33918" *) dat_pre_data[511:504] : dat_actv_data_reg2[511:504];
  assign _00317_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33908" *) dat_pre_data[503:496] : dat_actv_data_reg2[503:496];
  assign _00316_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33898" *) dat_pre_data[495:488] : dat_actv_data_reg2[495:488];
  assign _00315_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33888" *) dat_pre_data[487:480] : dat_actv_data_reg2[487:480];
  assign _00313_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33878" *) dat_pre_data[479:472] : dat_actv_data_reg2[479:472];
  assign _00312_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33868" *) dat_pre_data[471:464] : dat_actv_data_reg2[471:464];
  assign _00311_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33858" *) dat_pre_data[463:456] : dat_actv_data_reg2[463:456];
  assign _00310_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33848" *) dat_pre_data[455:448] : dat_actv_data_reg2[455:448];
  assign _00309_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33838" *) dat_pre_data[447:440] : dat_actv_data_reg2[447:440];
  assign _00308_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33828" *) dat_pre_data[439:432] : dat_actv_data_reg2[439:432];
  assign _00307_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33818" *) dat_pre_data[431:424] : dat_actv_data_reg2[431:424];
  assign _00306_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33808" *) dat_pre_data[423:416] : dat_actv_data_reg2[423:416];
  assign _00305_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33798" *) dat_pre_data[415:408] : dat_actv_data_reg2[415:408];
  assign _00304_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33788" *) dat_pre_data[407:400] : dat_actv_data_reg2[407:400];
  assign _00302_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33778" *) dat_pre_data[399:392] : dat_actv_data_reg2[399:392];
  assign _00301_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33768" *) dat_pre_data[391:384] : dat_actv_data_reg2[391:384];
  assign _00300_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33758" *) dat_pre_data[383:376] : dat_actv_data_reg2[383:376];
  assign _00299_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33748" *) dat_pre_data[375:368] : dat_actv_data_reg2[375:368];
  assign _00298_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33738" *) dat_pre_data[367:360] : dat_actv_data_reg2[367:360];
  assign _00297_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33728" *) dat_pre_data[359:352] : dat_actv_data_reg2[359:352];
  assign _00296_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33718" *) dat_pre_data[351:344] : dat_actv_data_reg2[351:344];
  assign _00295_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33708" *) dat_pre_data[343:336] : dat_actv_data_reg2[343:336];
  assign _00294_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33698" *) dat_pre_data[335:328] : dat_actv_data_reg2[335:328];
  assign _00293_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33688" *) dat_pre_data[327:320] : dat_actv_data_reg2[327:320];
  assign _00291_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33678" *) dat_pre_data[319:312] : dat_actv_data_reg2[319:312];
  assign _00290_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33668" *) dat_pre_data[311:304] : dat_actv_data_reg2[311:304];
  assign _00289_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33658" *) dat_pre_data[303:296] : dat_actv_data_reg2[303:296];
  assign _00288_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33648" *) dat_pre_data[295:288] : dat_actv_data_reg2[295:288];
  assign _00287_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33638" *) dat_pre_data[287:280] : dat_actv_data_reg2[287:280];
  assign _00286_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33628" *) dat_pre_data[279:272] : dat_actv_data_reg2[279:272];
  assign _00285_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33618" *) dat_pre_data[271:264] : dat_actv_data_reg2[271:264];
  assign _00284_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33608" *) dat_pre_data[263:256] : dat_actv_data_reg2[263:256];
  assign _00283_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33598" *) dat_pre_data[255:248] : dat_actv_data_reg2[255:248];
  assign _00282_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33588" *) dat_pre_data[247:240] : dat_actv_data_reg2[247:240];
  assign _00280_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33578" *) dat_pre_data[239:232] : dat_actv_data_reg2[239:232];
  assign _00279_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33568" *) dat_pre_data[231:224] : dat_actv_data_reg2[231:224];
  assign _00278_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33558" *) dat_pre_data[223:216] : dat_actv_data_reg2[223:216];
  assign _00277_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33548" *) dat_pre_data[215:208] : dat_actv_data_reg2[215:208];
  assign _00276_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33538" *) dat_pre_data[207:200] : dat_actv_data_reg2[207:200];
  assign _00275_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33528" *) dat_pre_data[199:192] : dat_actv_data_reg2[199:192];
  assign _00274_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33518" *) dat_pre_data[191:184] : dat_actv_data_reg2[191:184];
  assign _00273_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33508" *) dat_pre_data[183:176] : dat_actv_data_reg2[183:176];
  assign _00272_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33498" *) dat_pre_data[175:168] : dat_actv_data_reg2[175:168];
  assign _00271_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33488" *) dat_pre_data[167:160] : dat_actv_data_reg2[167:160];
  assign _00269_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33478" *) dat_pre_data[159:152] : dat_actv_data_reg2[159:152];
  assign _00268_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33468" *) dat_pre_data[151:144] : dat_actv_data_reg2[151:144];
  assign _00267_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33458" *) dat_pre_data[143:136] : dat_actv_data_reg2[143:136];
  assign _00266_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33448" *) dat_pre_data[135:128] : dat_actv_data_reg2[135:128];
  assign _00265_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33438" *) dat_pre_data[127:120] : dat_actv_data_reg2[127:120];
  assign _00264_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33428" *) dat_pre_data[119:112] : dat_actv_data_reg2[119:112];
  assign _00263_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33418" *) dat_pre_data[111:104] : dat_actv_data_reg2[111:104];
  assign _00262_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33408" *) dat_pre_data[103:96] : dat_actv_data_reg2[103:96];
  assign _00381_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33398" *) dat_pre_data[95:88] : dat_actv_data_reg2[95:88];
  assign _00370_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33388" *) dat_pre_data[87:80] : dat_actv_data_reg2[87:80];
  assign _00358_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33378" *) dat_pre_data[79:72] : dat_actv_data_reg2[79:72];
  assign _00347_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33368" *) dat_pre_data[71:64] : dat_actv_data_reg2[71:64];
  assign _00336_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33358" *) dat_pre_data[63:56] : dat_actv_data_reg2[63:56];
  assign _00325_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33348" *) dat_pre_data[55:48] : dat_actv_data_reg2[55:48];
  assign _00314_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33338" *) dat_pre_data[47:40] : dat_actv_data_reg2[47:40];
  assign _00303_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33328" *) dat_pre_data[39:32] : dat_actv_data_reg2[39:32];
  assign _00292_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33318" *) dat_pre_data[31:24] : dat_actv_data_reg2[31:24];
  assign _00281_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33308" *) dat_pre_data[23:16] : dat_actv_data_reg2[23:16];
  assign _00270_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33298" *) dat_pre_data[15:8] : dat_actv_data_reg2[15:8];
  assign _00359_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33288" *) dat_pre_data[7:0] : dat_actv_data_reg2[7:0];
  assign _01029_ = _05693_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33278" *) dat_pre_nan : dat_actv_nan_reg2;
  assign _01037_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33268" *) dat_pre_nz : dat_actv_nz_reg2;
  assign _00133_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33251" *) dat_pre_data[1023:1016] : dat_actv_data_reg1[1023:1016];
  assign _00132_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33241" *) dat_pre_data[1015:1008] : dat_actv_data_reg1[1015:1008];
  assign _00131_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33231" *) dat_pre_data[1007:1000] : dat_actv_data_reg1[1007:1000];
  assign _00258_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33221" *) dat_pre_data[999:992] : dat_actv_data_reg1[999:992];
  assign _00257_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33211" *) dat_pre_data[991:984] : dat_actv_data_reg1[991:984];
  assign _00256_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33201" *) dat_pre_data[983:976] : dat_actv_data_reg1[983:976];
  assign _00255_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33191" *) dat_pre_data[975:968] : dat_actv_data_reg1[975:968];
  assign _00254_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33181" *) dat_pre_data[967:960] : dat_actv_data_reg1[967:960];
  assign _00252_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33171" *) dat_pre_data[959:952] : dat_actv_data_reg1[959:952];
  assign _00251_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33161" *) dat_pre_data[951:944] : dat_actv_data_reg1[951:944];
  assign _00250_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33151" *) dat_pre_data[943:936] : dat_actv_data_reg1[943:936];
  assign _00249_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33141" *) dat_pre_data[935:928] : dat_actv_data_reg1[935:928];
  assign _00248_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33131" *) dat_pre_data[927:920] : dat_actv_data_reg1[927:920];
  assign _00247_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33121" *) dat_pre_data[919:912] : dat_actv_data_reg1[919:912];
  assign _00246_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33111" *) dat_pre_data[911:904] : dat_actv_data_reg1[911:904];
  assign _00245_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33101" *) dat_pre_data[903:896] : dat_actv_data_reg1[903:896];
  assign _00244_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33091" *) dat_pre_data[895:888] : dat_actv_data_reg1[895:888];
  assign _00243_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33081" *) dat_pre_data[887:880] : dat_actv_data_reg1[887:880];
  assign _00241_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33071" *) dat_pre_data[879:872] : dat_actv_data_reg1[879:872];
  assign _00240_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33061" *) dat_pre_data[871:864] : dat_actv_data_reg1[871:864];
  assign _00239_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33051" *) dat_pre_data[863:856] : dat_actv_data_reg1[863:856];
  assign _00238_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33041" *) dat_pre_data[855:848] : dat_actv_data_reg1[855:848];
  assign _00237_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33031" *) dat_pre_data[847:840] : dat_actv_data_reg1[847:840];
  assign _00236_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33021" *) dat_pre_data[839:832] : dat_actv_data_reg1[839:832];
  assign _00235_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33011" *) dat_pre_data[831:824] : dat_actv_data_reg1[831:824];
  assign _00234_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:33001" *) dat_pre_data[823:816] : dat_actv_data_reg1[823:816];
  assign _00233_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32991" *) dat_pre_data[815:808] : dat_actv_data_reg1[815:808];
  assign _00232_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32981" *) dat_pre_data[807:800] : dat_actv_data_reg1[807:800];
  assign _00229_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32971" *) dat_pre_data[799:792] : dat_actv_data_reg1[799:792];
  assign _00228_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32961" *) dat_pre_data[791:784] : dat_actv_data_reg1[791:784];
  assign _00227_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32951" *) dat_pre_data[783:776] : dat_actv_data_reg1[783:776];
  assign _00226_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32941" *) dat_pre_data[775:768] : dat_actv_data_reg1[775:768];
  assign _00225_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32931" *) dat_pre_data[767:760] : dat_actv_data_reg1[767:760];
  assign _00224_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32921" *) dat_pre_data[759:752] : dat_actv_data_reg1[759:752];
  assign _00223_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32911" *) dat_pre_data[751:744] : dat_actv_data_reg1[751:744];
  assign _00222_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32901" *) dat_pre_data[743:736] : dat_actv_data_reg1[743:736];
  assign _00221_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32891" *) dat_pre_data[735:728] : dat_actv_data_reg1[735:728];
  assign _00220_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32881" *) dat_pre_data[727:720] : dat_actv_data_reg1[727:720];
  assign _00218_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32871" *) dat_pre_data[719:712] : dat_actv_data_reg1[719:712];
  assign _00217_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32861" *) dat_pre_data[711:704] : dat_actv_data_reg1[711:704];
  assign _00216_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32851" *) dat_pre_data[703:696] : dat_actv_data_reg1[703:696];
  assign _00215_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32841" *) dat_pre_data[695:688] : dat_actv_data_reg1[695:688];
  assign _00214_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32831" *) dat_pre_data[687:680] : dat_actv_data_reg1[687:680];
  assign _00213_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32821" *) dat_pre_data[679:672] : dat_actv_data_reg1[679:672];
  assign _00212_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32811" *) dat_pre_data[671:664] : dat_actv_data_reg1[671:664];
  assign _00211_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32801" *) dat_pre_data[663:656] : dat_actv_data_reg1[663:656];
  assign _00210_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32791" *) dat_pre_data[655:648] : dat_actv_data_reg1[655:648];
  assign _00209_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32781" *) dat_pre_data[647:640] : dat_actv_data_reg1[647:640];
  assign _00207_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32771" *) dat_pre_data[639:632] : dat_actv_data_reg1[639:632];
  assign _00206_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32761" *) dat_pre_data[631:624] : dat_actv_data_reg1[631:624];
  assign _00205_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32751" *) dat_pre_data[623:616] : dat_actv_data_reg1[623:616];
  assign _00204_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32741" *) dat_pre_data[615:608] : dat_actv_data_reg1[615:608];
  assign _00203_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32731" *) dat_pre_data[607:600] : dat_actv_data_reg1[607:600];
  assign _00202_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32721" *) dat_pre_data[599:592] : dat_actv_data_reg1[599:592];
  assign _00201_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32711" *) dat_pre_data[591:584] : dat_actv_data_reg1[591:584];
  assign _00200_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32701" *) dat_pre_data[583:576] : dat_actv_data_reg1[583:576];
  assign _00199_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32691" *) dat_pre_data[575:568] : dat_actv_data_reg1[575:568];
  assign _00198_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32681" *) dat_pre_data[567:560] : dat_actv_data_reg1[567:560];
  assign _00196_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32671" *) dat_pre_data[559:552] : dat_actv_data_reg1[559:552];
  assign _00195_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32661" *) dat_pre_data[551:544] : dat_actv_data_reg1[551:544];
  assign _00194_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32651" *) dat_pre_data[543:536] : dat_actv_data_reg1[543:536];
  assign _00193_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32641" *) dat_pre_data[535:528] : dat_actv_data_reg1[535:528];
  assign _00192_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32631" *) dat_pre_data[527:520] : dat_actv_data_reg1[527:520];
  assign _00191_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32621" *) dat_pre_data[519:512] : dat_actv_data_reg1[519:512];
  assign _00190_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32611" *) dat_pre_data[511:504] : dat_actv_data_reg1[511:504];
  assign _00189_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32601" *) dat_pre_data[503:496] : dat_actv_data_reg1[503:496];
  assign _00188_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32591" *) dat_pre_data[495:488] : dat_actv_data_reg1[495:488];
  assign _00187_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32581" *) dat_pre_data[487:480] : dat_actv_data_reg1[487:480];
  assign _00185_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32571" *) dat_pre_data[479:472] : dat_actv_data_reg1[479:472];
  assign _00184_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32561" *) dat_pre_data[471:464] : dat_actv_data_reg1[471:464];
  assign _00183_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32551" *) dat_pre_data[463:456] : dat_actv_data_reg1[463:456];
  assign _00182_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32541" *) dat_pre_data[455:448] : dat_actv_data_reg1[455:448];
  assign _00181_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32531" *) dat_pre_data[447:440] : dat_actv_data_reg1[447:440];
  assign _00180_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32521" *) dat_pre_data[439:432] : dat_actv_data_reg1[439:432];
  assign _00179_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32511" *) dat_pre_data[431:424] : dat_actv_data_reg1[431:424];
  assign _00178_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32501" *) dat_pre_data[423:416] : dat_actv_data_reg1[423:416];
  assign _00177_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32491" *) dat_pre_data[415:408] : dat_actv_data_reg1[415:408];
  assign _00176_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32481" *) dat_pre_data[407:400] : dat_actv_data_reg1[407:400];
  assign _00174_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32471" *) dat_pre_data[399:392] : dat_actv_data_reg1[399:392];
  assign _00173_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32461" *) dat_pre_data[391:384] : dat_actv_data_reg1[391:384];
  assign _00172_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32451" *) dat_pre_data[383:376] : dat_actv_data_reg1[383:376];
  assign _00171_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32441" *) dat_pre_data[375:368] : dat_actv_data_reg1[375:368];
  assign _00170_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32431" *) dat_pre_data[367:360] : dat_actv_data_reg1[367:360];
  assign _00169_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32421" *) dat_pre_data[359:352] : dat_actv_data_reg1[359:352];
  assign _00168_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32411" *) dat_pre_data[351:344] : dat_actv_data_reg1[351:344];
  assign _00167_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32401" *) dat_pre_data[343:336] : dat_actv_data_reg1[343:336];
  assign _00166_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32391" *) dat_pre_data[335:328] : dat_actv_data_reg1[335:328];
  assign _00165_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32381" *) dat_pre_data[327:320] : dat_actv_data_reg1[327:320];
  assign _00163_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32371" *) dat_pre_data[319:312] : dat_actv_data_reg1[319:312];
  assign _00162_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32361" *) dat_pre_data[311:304] : dat_actv_data_reg1[311:304];
  assign _00161_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32351" *) dat_pre_data[303:296] : dat_actv_data_reg1[303:296];
  assign _00160_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32341" *) dat_pre_data[295:288] : dat_actv_data_reg1[295:288];
  assign _00159_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32331" *) dat_pre_data[287:280] : dat_actv_data_reg1[287:280];
  assign _00158_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32321" *) dat_pre_data[279:272] : dat_actv_data_reg1[279:272];
  assign _00157_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32311" *) dat_pre_data[271:264] : dat_actv_data_reg1[271:264];
  assign _00156_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32301" *) dat_pre_data[263:256] : dat_actv_data_reg1[263:256];
  assign _00155_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32291" *) dat_pre_data[255:248] : dat_actv_data_reg1[255:248];
  assign _00154_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32281" *) dat_pre_data[247:240] : dat_actv_data_reg1[247:240];
  assign _00152_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32271" *) dat_pre_data[239:232] : dat_actv_data_reg1[239:232];
  assign _00151_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32261" *) dat_pre_data[231:224] : dat_actv_data_reg1[231:224];
  assign _00150_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32251" *) dat_pre_data[223:216] : dat_actv_data_reg1[223:216];
  assign _00149_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32241" *) dat_pre_data[215:208] : dat_actv_data_reg1[215:208];
  assign _00148_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32231" *) dat_pre_data[207:200] : dat_actv_data_reg1[207:200];
  assign _00147_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32221" *) dat_pre_data[199:192] : dat_actv_data_reg1[199:192];
  assign _00146_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32211" *) dat_pre_data[191:184] : dat_actv_data_reg1[191:184];
  assign _00145_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32201" *) dat_pre_data[183:176] : dat_actv_data_reg1[183:176];
  assign _00144_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32191" *) dat_pre_data[175:168] : dat_actv_data_reg1[175:168];
  assign _00143_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32181" *) dat_pre_data[167:160] : dat_actv_data_reg1[167:160];
  assign _00141_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32171" *) dat_pre_data[159:152] : dat_actv_data_reg1[159:152];
  assign _00140_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32161" *) dat_pre_data[151:144] : dat_actv_data_reg1[151:144];
  assign _00139_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32151" *) dat_pre_data[143:136] : dat_actv_data_reg1[143:136];
  assign _00138_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32141" *) dat_pre_data[135:128] : dat_actv_data_reg1[135:128];
  assign _00137_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32131" *) dat_pre_data[127:120] : dat_actv_data_reg1[127:120];
  assign _00136_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32121" *) dat_pre_data[119:112] : dat_actv_data_reg1[119:112];
  assign _00135_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32111" *) dat_pre_data[111:104] : dat_actv_data_reg1[111:104];
  assign _00134_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32101" *) dat_pre_data[103:96] : dat_actv_data_reg1[103:96];
  assign _00253_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32091" *) dat_pre_data[95:88] : dat_actv_data_reg1[95:88];
  assign _00242_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32081" *) dat_pre_data[87:80] : dat_actv_data_reg1[87:80];
  assign _00230_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32071" *) dat_pre_data[79:72] : dat_actv_data_reg1[79:72];
  assign _00219_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32061" *) dat_pre_data[71:64] : dat_actv_data_reg1[71:64];
  assign _00208_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32051" *) dat_pre_data[63:56] : dat_actv_data_reg1[63:56];
  assign _00197_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32041" *) dat_pre_data[55:48] : dat_actv_data_reg1[55:48];
  assign _00186_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32031" *) dat_pre_data[47:40] : dat_actv_data_reg1[47:40];
  assign _00175_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32021" *) dat_pre_data[39:32] : dat_actv_data_reg1[39:32];
  assign _00164_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32011" *) dat_pre_data[31:24] : dat_actv_data_reg1[31:24];
  assign _00153_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:32001" *) dat_pre_data[23:16] : dat_actv_data_reg1[23:16];
  assign _00142_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31991" *) dat_pre_data[15:8] : dat_actv_data_reg1[15:8];
  assign _00231_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31981" *) dat_pre_data[7:0] : dat_actv_data_reg1[7:0];
  assign _01028_ = _05692_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31971" *) dat_pre_nan : dat_actv_nan_reg1;
  assign _01036_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31961" *) dat_pre_nz : dat_actv_nz_reg1;
  assign _00005_ = _05691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31944" *) dat_pre_data[1023:1016] : dat_actv_data_reg0[1023:1016];
  assign _00004_ = _05690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31934" *) dat_pre_data[1015:1008] : dat_actv_data_reg0[1015:1008];
  assign _00003_ = _05689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31924" *) dat_pre_data[1007:1000] : dat_actv_data_reg0[1007:1000];
  assign _00130_ = _05688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31914" *) dat_pre_data[999:992] : dat_actv_data_reg0[999:992];
  assign _00129_ = _05687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31904" *) dat_pre_data[991:984] : dat_actv_data_reg0[991:984];
  assign _00128_ = _05686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31894" *) dat_pre_data[983:976] : dat_actv_data_reg0[983:976];
  assign _00127_ = _05685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31884" *) dat_pre_data[975:968] : dat_actv_data_reg0[975:968];
  assign _00126_ = _05684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31874" *) dat_pre_data[967:960] : dat_actv_data_reg0[967:960];
  assign _00124_ = _05683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31864" *) dat_pre_data[959:952] : dat_actv_data_reg0[959:952];
  assign _00123_ = _05682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31854" *) dat_pre_data[951:944] : dat_actv_data_reg0[951:944];
  assign _00122_ = _05681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31844" *) dat_pre_data[943:936] : dat_actv_data_reg0[943:936];
  assign _00121_ = _05680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31834" *) dat_pre_data[935:928] : dat_actv_data_reg0[935:928];
  assign _00120_ = _05679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31824" *) dat_pre_data[927:920] : dat_actv_data_reg0[927:920];
  assign _00119_ = _05678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31814" *) dat_pre_data[919:912] : dat_actv_data_reg0[919:912];
  assign _00118_ = _05677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31804" *) dat_pre_data[911:904] : dat_actv_data_reg0[911:904];
  assign _00117_ = _05676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31794" *) dat_pre_data[903:896] : dat_actv_data_reg0[903:896];
  assign _00116_ = _05675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31784" *) dat_pre_data[895:888] : dat_actv_data_reg0[895:888];
  assign _00115_ = _05674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31774" *) dat_pre_data[887:880] : dat_actv_data_reg0[887:880];
  assign _00113_ = _05673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31764" *) dat_pre_data[879:872] : dat_actv_data_reg0[879:872];
  assign _00112_ = _05672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31754" *) dat_pre_data[871:864] : dat_actv_data_reg0[871:864];
  assign _00111_ = _05671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31744" *) dat_pre_data[863:856] : dat_actv_data_reg0[863:856];
  assign _00110_ = _05670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31734" *) dat_pre_data[855:848] : dat_actv_data_reg0[855:848];
  assign _00109_ = _05669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31724" *) dat_pre_data[847:840] : dat_actv_data_reg0[847:840];
  assign _00108_ = _05668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31714" *) dat_pre_data[839:832] : dat_actv_data_reg0[839:832];
  assign _00107_ = _05667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31704" *) dat_pre_data[831:824] : dat_actv_data_reg0[831:824];
  assign _00106_ = _05666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31694" *) dat_pre_data[823:816] : dat_actv_data_reg0[823:816];
  assign _00105_ = _05665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31684" *) dat_pre_data[815:808] : dat_actv_data_reg0[815:808];
  assign _00104_ = _05664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31674" *) dat_pre_data[807:800] : dat_actv_data_reg0[807:800];
  assign _00101_ = _05663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31664" *) dat_pre_data[799:792] : dat_actv_data_reg0[799:792];
  assign _00100_ = _05662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31654" *) dat_pre_data[791:784] : dat_actv_data_reg0[791:784];
  assign _00099_ = _05661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31644" *) dat_pre_data[783:776] : dat_actv_data_reg0[783:776];
  assign _00098_ = _05660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31634" *) dat_pre_data[775:768] : dat_actv_data_reg0[775:768];
  assign _00097_ = _05659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31624" *) dat_pre_data[767:760] : dat_actv_data_reg0[767:760];
  assign _00096_ = _05658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31614" *) dat_pre_data[759:752] : dat_actv_data_reg0[759:752];
  assign _00095_ = _05657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31604" *) dat_pre_data[751:744] : dat_actv_data_reg0[751:744];
  assign _00094_ = _05656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31594" *) dat_pre_data[743:736] : dat_actv_data_reg0[743:736];
  assign _00093_ = _05655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31584" *) dat_pre_data[735:728] : dat_actv_data_reg0[735:728];
  assign _00092_ = _05654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31574" *) dat_pre_data[727:720] : dat_actv_data_reg0[727:720];
  assign _00090_ = _05653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31564" *) dat_pre_data[719:712] : dat_actv_data_reg0[719:712];
  assign _00089_ = _05652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31554" *) dat_pre_data[711:704] : dat_actv_data_reg0[711:704];
  assign _00088_ = _05651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31544" *) dat_pre_data[703:696] : dat_actv_data_reg0[703:696];
  assign _00087_ = _05650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31534" *) dat_pre_data[695:688] : dat_actv_data_reg0[695:688];
  assign _00086_ = _05649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31524" *) dat_pre_data[687:680] : dat_actv_data_reg0[687:680];
  assign _00085_ = _05648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31514" *) dat_pre_data[679:672] : dat_actv_data_reg0[679:672];
  assign _00084_ = _05647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31504" *) dat_pre_data[671:664] : dat_actv_data_reg0[671:664];
  assign _00083_ = _05646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31494" *) dat_pre_data[663:656] : dat_actv_data_reg0[663:656];
  assign _00082_ = _05645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31484" *) dat_pre_data[655:648] : dat_actv_data_reg0[655:648];
  assign _00081_ = _05644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31474" *) dat_pre_data[647:640] : dat_actv_data_reg0[647:640];
  assign _00079_ = _05643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31464" *) dat_pre_data[639:632] : dat_actv_data_reg0[639:632];
  assign _00078_ = _05642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31454" *) dat_pre_data[631:624] : dat_actv_data_reg0[631:624];
  assign _00077_ = _05641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31444" *) dat_pre_data[623:616] : dat_actv_data_reg0[623:616];
  assign _00076_ = _05640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31434" *) dat_pre_data[615:608] : dat_actv_data_reg0[615:608];
  assign _00075_ = _05639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31424" *) dat_pre_data[607:600] : dat_actv_data_reg0[607:600];
  assign _00074_ = _05638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31414" *) dat_pre_data[599:592] : dat_actv_data_reg0[599:592];
  assign _00073_ = _05637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31404" *) dat_pre_data[591:584] : dat_actv_data_reg0[591:584];
  assign _00072_ = _05636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31394" *) dat_pre_data[583:576] : dat_actv_data_reg0[583:576];
  assign _00071_ = _05635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31384" *) dat_pre_data[575:568] : dat_actv_data_reg0[575:568];
  assign _00070_ = _05634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31374" *) dat_pre_data[567:560] : dat_actv_data_reg0[567:560];
  assign _00068_ = _05633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31364" *) dat_pre_data[559:552] : dat_actv_data_reg0[559:552];
  assign _00067_ = _05632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31354" *) dat_pre_data[551:544] : dat_actv_data_reg0[551:544];
  assign _00066_ = _05631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31344" *) dat_pre_data[543:536] : dat_actv_data_reg0[543:536];
  assign _00065_ = _05630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31334" *) dat_pre_data[535:528] : dat_actv_data_reg0[535:528];
  assign _00064_ = _05629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31324" *) dat_pre_data[527:520] : dat_actv_data_reg0[527:520];
  assign _00063_ = _05628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31314" *) dat_pre_data[519:512] : dat_actv_data_reg0[519:512];
  assign _00062_ = _05627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31304" *) dat_pre_data[511:504] : dat_actv_data_reg0[511:504];
  assign _00061_ = _05626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31294" *) dat_pre_data[503:496] : dat_actv_data_reg0[503:496];
  assign _00060_ = _05625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31284" *) dat_pre_data[495:488] : dat_actv_data_reg0[495:488];
  assign _00059_ = _05624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31274" *) dat_pre_data[487:480] : dat_actv_data_reg0[487:480];
  assign _00057_ = _05623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31264" *) dat_pre_data[479:472] : dat_actv_data_reg0[479:472];
  assign _00056_ = _05622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31254" *) dat_pre_data[471:464] : dat_actv_data_reg0[471:464];
  assign _00055_ = _05621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31244" *) dat_pre_data[463:456] : dat_actv_data_reg0[463:456];
  assign _00054_ = _05620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31234" *) dat_pre_data[455:448] : dat_actv_data_reg0[455:448];
  assign _00053_ = _05619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31224" *) dat_pre_data[447:440] : dat_actv_data_reg0[447:440];
  assign _00052_ = _05618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31214" *) dat_pre_data[439:432] : dat_actv_data_reg0[439:432];
  assign _00051_ = _05617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31204" *) dat_pre_data[431:424] : dat_actv_data_reg0[431:424];
  assign _00050_ = _05616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31194" *) dat_pre_data[423:416] : dat_actv_data_reg0[423:416];
  assign _00049_ = _05615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31184" *) dat_pre_data[415:408] : dat_actv_data_reg0[415:408];
  assign _00048_ = _05614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31174" *) dat_pre_data[407:400] : dat_actv_data_reg0[407:400];
  assign _00046_ = _05613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31164" *) dat_pre_data[399:392] : dat_actv_data_reg0[399:392];
  assign _00045_ = _05612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31154" *) dat_pre_data[391:384] : dat_actv_data_reg0[391:384];
  assign _00044_ = _05611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31144" *) dat_pre_data[383:376] : dat_actv_data_reg0[383:376];
  assign _00043_ = _05610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31134" *) dat_pre_data[375:368] : dat_actv_data_reg0[375:368];
  assign _00042_ = _05609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31124" *) dat_pre_data[367:360] : dat_actv_data_reg0[367:360];
  assign _00041_ = _05608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31114" *) dat_pre_data[359:352] : dat_actv_data_reg0[359:352];
  assign _00040_ = _05607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31104" *) dat_pre_data[351:344] : dat_actv_data_reg0[351:344];
  assign _00039_ = _05606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31094" *) dat_pre_data[343:336] : dat_actv_data_reg0[343:336];
  assign _00038_ = _05605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31084" *) dat_pre_data[335:328] : dat_actv_data_reg0[335:328];
  assign _00037_ = _05604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31074" *) dat_pre_data[327:320] : dat_actv_data_reg0[327:320];
  assign _00035_ = _05603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31064" *) dat_pre_data[319:312] : dat_actv_data_reg0[319:312];
  assign _00034_ = _05602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31054" *) dat_pre_data[311:304] : dat_actv_data_reg0[311:304];
  assign _00033_ = _05601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31044" *) dat_pre_data[303:296] : dat_actv_data_reg0[303:296];
  assign _00032_ = _05600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31034" *) dat_pre_data[295:288] : dat_actv_data_reg0[295:288];
  assign _00031_ = _05599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31024" *) dat_pre_data[287:280] : dat_actv_data_reg0[287:280];
  assign _00030_ = _05598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31014" *) dat_pre_data[279:272] : dat_actv_data_reg0[279:272];
  assign _00029_ = _05597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:31004" *) dat_pre_data[271:264] : dat_actv_data_reg0[271:264];
  assign _00028_ = _05596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30994" *) dat_pre_data[263:256] : dat_actv_data_reg0[263:256];
  assign _00027_ = _05595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30984" *) dat_pre_data[255:248] : dat_actv_data_reg0[255:248];
  assign _00026_ = _05594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30974" *) dat_pre_data[247:240] : dat_actv_data_reg0[247:240];
  assign _00024_ = _05593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30964" *) dat_pre_data[239:232] : dat_actv_data_reg0[239:232];
  assign _00023_ = _05592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30954" *) dat_pre_data[231:224] : dat_actv_data_reg0[231:224];
  assign _00022_ = _05591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30944" *) dat_pre_data[223:216] : dat_actv_data_reg0[223:216];
  assign _00021_ = _05590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30934" *) dat_pre_data[215:208] : dat_actv_data_reg0[215:208];
  assign _00020_ = _05589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30924" *) dat_pre_data[207:200] : dat_actv_data_reg0[207:200];
  assign _00019_ = _05588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30914" *) dat_pre_data[199:192] : dat_actv_data_reg0[199:192];
  assign _00018_ = _05587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30904" *) dat_pre_data[191:184] : dat_actv_data_reg0[191:184];
  assign _00017_ = _05586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30894" *) dat_pre_data[183:176] : dat_actv_data_reg0[183:176];
  assign _00016_ = _05585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30884" *) dat_pre_data[175:168] : dat_actv_data_reg0[175:168];
  assign _00015_ = _05584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30874" *) dat_pre_data[167:160] : dat_actv_data_reg0[167:160];
  assign _00013_ = _05583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30864" *) dat_pre_data[159:152] : dat_actv_data_reg0[159:152];
  assign _00012_ = _05582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30854" *) dat_pre_data[151:144] : dat_actv_data_reg0[151:144];
  assign _00011_ = _05581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30844" *) dat_pre_data[143:136] : dat_actv_data_reg0[143:136];
  assign _00010_ = _05580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30834" *) dat_pre_data[135:128] : dat_actv_data_reg0[135:128];
  assign _00009_ = _05579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30824" *) dat_pre_data[127:120] : dat_actv_data_reg0[127:120];
  assign _00008_ = _05578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30814" *) dat_pre_data[119:112] : dat_actv_data_reg0[119:112];
  assign _00007_ = _05577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30804" *) dat_pre_data[111:104] : dat_actv_data_reg0[111:104];
  assign _00006_ = _05576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30794" *) dat_pre_data[103:96] : dat_actv_data_reg0[103:96];
  assign _00125_ = _05575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30784" *) dat_pre_data[95:88] : dat_actv_data_reg0[95:88];
  assign _00114_ = _05574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30774" *) dat_pre_data[87:80] : dat_actv_data_reg0[87:80];
  assign _00102_ = _05573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30764" *) dat_pre_data[79:72] : dat_actv_data_reg0[79:72];
  assign _00091_ = _05572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30754" *) dat_pre_data[71:64] : dat_actv_data_reg0[71:64];
  assign _00080_ = _05571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30744" *) dat_pre_data[63:56] : dat_actv_data_reg0[63:56];
  assign _00069_ = _05570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30734" *) dat_pre_data[55:48] : dat_actv_data_reg0[55:48];
  assign _00058_ = _05569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30724" *) dat_pre_data[47:40] : dat_actv_data_reg0[47:40];
  assign _00047_ = _05568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30714" *) dat_pre_data[39:32] : dat_actv_data_reg0[39:32];
  assign _00036_ = _05567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30704" *) dat_pre_data[31:24] : dat_actv_data_reg0[31:24];
  assign _00025_ = _05566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30694" *) dat_pre_data[23:16] : dat_actv_data_reg0[23:16];
  assign _00014_ = _05565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30684" *) dat_pre_data[15:8] : dat_actv_data_reg0[15:8];
  assign _00103_ = _05564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30674" *) dat_pre_data[7:0] : dat_actv_data_reg0[7:0];
  assign _01027_ = _05563_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30664" *) dat_pre_nan : dat_actv_nan_reg0;
  assign _01035_ = dat_pre_pvld[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30654" *) dat_pre_nz : dat_actv_nz_reg0;
  assign _01178_ = _05562_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30530" *) dat_pre_exp_w : dat_pre_exp_reg7;
  assign _01186_ = _05562_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30520" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask7;
  assign _01177_ = _05561_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30510" *) dat_pre_exp_w : dat_pre_exp_reg6;
  assign _01185_ = _05561_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30500" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask6;
  assign _01176_ = _05560_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30490" *) dat_pre_exp_w : dat_pre_exp_reg5;
  assign _01184_ = _05560_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30480" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask5;
  assign _01175_ = _05559_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30470" *) dat_pre_exp_w : dat_pre_exp_reg4;
  assign _01183_ = _05559_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30460" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask4;
  assign _01174_ = _05558_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30450" *) dat_pre_exp_w : dat_pre_exp_reg3;
  assign _01182_ = _05558_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30440" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask3;
  assign _01173_ = _05557_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30430" *) dat_pre_exp_w : dat_pre_exp_reg2;
  assign _01181_ = _05557_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30420" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask2;
  assign _01172_ = _05556_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30410" *) dat_pre_exp_w : dat_pre_exp_reg1;
  assign _01180_ = _05556_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30400" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask1;
  assign _01171_ = _05555_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30390" *) dat_pre_exp_w : dat_pre_exp_reg0;
  assign _01179_ = _05555_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30380" *) { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] } : dat_pre_mask0;
  assign _01045_ = _05554_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30356" *) dat_pre_data_w[1023:1016] : dat_pre_data[1023:1016];
  assign _01044_ = _05553_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30346" *) dat_pre_data_w[1015:1008] : dat_pre_data[1015:1008];
  assign _01043_ = _05552_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30336" *) dat_pre_data_w[1007:1000] : dat_pre_data[1007:1000];
  assign _01170_ = _05551_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30326" *) dat_pre_data_w[999:992] : dat_pre_data[999:992];
  assign _01169_ = _05550_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30316" *) dat_pre_data_w[991:984] : dat_pre_data[991:984];
  assign _01168_ = _05549_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30306" *) dat_pre_data_w[983:976] : dat_pre_data[983:976];
  assign _01167_ = _05548_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30296" *) dat_pre_data_w[975:968] : dat_pre_data[975:968];
  assign _01166_ = _05547_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30286" *) dat_pre_data_w[967:960] : dat_pre_data[967:960];
  assign _01164_ = _05546_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30276" *) dat_pre_data_w[959:952] : dat_pre_data[959:952];
  assign _01163_ = _05545_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30266" *) dat_pre_data_w[951:944] : dat_pre_data[951:944];
  assign _01162_ = _05544_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30256" *) dat_pre_data_w[943:936] : dat_pre_data[943:936];
  assign _01161_ = _05543_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30246" *) dat_pre_data_w[935:928] : dat_pre_data[935:928];
  assign _01160_ = _05542_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30236" *) dat_pre_data_w[927:920] : dat_pre_data[927:920];
  assign _01159_ = _05541_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30226" *) dat_pre_data_w[919:912] : dat_pre_data[919:912];
  assign _01158_ = _05540_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30216" *) dat_pre_data_w[911:904] : dat_pre_data[911:904];
  assign _01157_ = _05539_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30206" *) dat_pre_data_w[903:896] : dat_pre_data[903:896];
  assign _01156_ = _05538_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30196" *) dat_pre_data_w[895:888] : dat_pre_data[895:888];
  assign _01155_ = _05537_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30186" *) dat_pre_data_w[887:880] : dat_pre_data[887:880];
  assign _01153_ = _05536_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30176" *) dat_pre_data_w[879:872] : dat_pre_data[879:872];
  assign _01152_ = _05535_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30166" *) dat_pre_data_w[871:864] : dat_pre_data[871:864];
  assign _01151_ = _05534_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30156" *) dat_pre_data_w[863:856] : dat_pre_data[863:856];
  assign _01150_ = _05533_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30146" *) dat_pre_data_w[855:848] : dat_pre_data[855:848];
  assign _01149_ = _05532_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30136" *) dat_pre_data_w[847:840] : dat_pre_data[847:840];
  assign _01148_ = _05531_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30126" *) dat_pre_data_w[839:832] : dat_pre_data[839:832];
  assign _01147_ = _05530_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30116" *) dat_pre_data_w[831:824] : dat_pre_data[831:824];
  assign _01146_ = _05529_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30106" *) dat_pre_data_w[823:816] : dat_pre_data[823:816];
  assign _01145_ = _05528_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30096" *) dat_pre_data_w[815:808] : dat_pre_data[815:808];
  assign _01144_ = _05527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30086" *) dat_pre_data_w[807:800] : dat_pre_data[807:800];
  assign _01141_ = _05526_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30076" *) dat_pre_data_w[799:792] : dat_pre_data[799:792];
  assign _01140_ = _05525_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30066" *) dat_pre_data_w[791:784] : dat_pre_data[791:784];
  assign _01139_ = _05524_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30056" *) dat_pre_data_w[783:776] : dat_pre_data[783:776];
  assign _01138_ = _05523_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30046" *) dat_pre_data_w[775:768] : dat_pre_data[775:768];
  assign _01137_ = _05522_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30036" *) dat_pre_data_w[767:760] : dat_pre_data[767:760];
  assign _01136_ = _05521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30026" *) dat_pre_data_w[759:752] : dat_pre_data[759:752];
  assign _01135_ = _05520_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30016" *) dat_pre_data_w[751:744] : dat_pre_data[751:744];
  assign _01134_ = _05519_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:30006" *) dat_pre_data_w[743:736] : dat_pre_data[743:736];
  assign _01133_ = _05518_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29996" *) dat_pre_data_w[735:728] : dat_pre_data[735:728];
  assign _01132_ = _05517_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29986" *) dat_pre_data_w[727:720] : dat_pre_data[727:720];
  assign _01130_ = _05516_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29976" *) dat_pre_data_w[719:712] : dat_pre_data[719:712];
  assign _01129_ = _05515_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29966" *) dat_pre_data_w[711:704] : dat_pre_data[711:704];
  assign _01128_ = _05514_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29956" *) dat_pre_data_w[703:696] : dat_pre_data[703:696];
  assign _01127_ = _05513_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29946" *) dat_pre_data_w[695:688] : dat_pre_data[695:688];
  assign _01126_ = _05512_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29936" *) dat_pre_data_w[687:680] : dat_pre_data[687:680];
  assign _01125_ = _05511_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29926" *) dat_pre_data_w[679:672] : dat_pre_data[679:672];
  assign _01124_ = _05510_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29916" *) dat_pre_data_w[671:664] : dat_pre_data[671:664];
  assign _01123_ = _05509_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29906" *) dat_pre_data_w[663:656] : dat_pre_data[663:656];
  assign _01122_ = _05508_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29896" *) dat_pre_data_w[655:648] : dat_pre_data[655:648];
  assign _01121_ = _05507_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29886" *) dat_pre_data_w[647:640] : dat_pre_data[647:640];
  assign _01119_ = _05506_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29876" *) dat_pre_data_w[639:632] : dat_pre_data[639:632];
  assign _01118_ = _05505_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29866" *) dat_pre_data_w[631:624] : dat_pre_data[631:624];
  assign _01117_ = _05504_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29856" *) dat_pre_data_w[623:616] : dat_pre_data[623:616];
  assign _01116_ = _05503_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29846" *) dat_pre_data_w[615:608] : dat_pre_data[615:608];
  assign _01115_ = _05502_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29836" *) dat_pre_data_w[607:600] : dat_pre_data[607:600];
  assign _01114_ = _05501_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29826" *) dat_pre_data_w[599:592] : dat_pre_data[599:592];
  assign _01113_ = _05500_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29816" *) dat_pre_data_w[591:584] : dat_pre_data[591:584];
  assign _01112_ = _05499_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29806" *) dat_pre_data_w[583:576] : dat_pre_data[583:576];
  assign _01111_ = _05498_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29796" *) dat_pre_data_w[575:568] : dat_pre_data[575:568];
  assign _01110_ = _05497_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29786" *) dat_pre_data_w[567:560] : dat_pre_data[567:560];
  assign _01108_ = _05496_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29776" *) dat_pre_data_w[559:552] : dat_pre_data[559:552];
  assign _01107_ = _05495_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29766" *) dat_pre_data_w[551:544] : dat_pre_data[551:544];
  assign _01106_ = _05494_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29756" *) dat_pre_data_w[543:536] : dat_pre_data[543:536];
  assign _01105_ = _05493_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29746" *) dat_pre_data_w[535:528] : dat_pre_data[535:528];
  assign _01104_ = _05492_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29736" *) dat_pre_data_w[527:520] : dat_pre_data[527:520];
  assign _01103_ = _05491_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29726" *) dat_pre_data_w[519:512] : dat_pre_data[519:512];
  assign _01102_ = _05490_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29716" *) dat_pre_data_w[511:504] : dat_pre_data[511:504];
  assign _01101_ = _05489_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29706" *) dat_pre_data_w[503:496] : dat_pre_data[503:496];
  assign _01100_ = _05488_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29696" *) dat_pre_data_w[495:488] : dat_pre_data[495:488];
  assign _01099_ = _05487_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29686" *) dat_pre_data_w[487:480] : dat_pre_data[487:480];
  assign _01097_ = _05486_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29676" *) dat_pre_data_w[479:472] : dat_pre_data[479:472];
  assign _01096_ = _05485_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29666" *) dat_pre_data_w[471:464] : dat_pre_data[471:464];
  assign _01095_ = _05484_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29656" *) dat_pre_data_w[463:456] : dat_pre_data[463:456];
  assign _01094_ = _05483_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29646" *) dat_pre_data_w[455:448] : dat_pre_data[455:448];
  assign _01093_ = _05482_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29636" *) dat_pre_data_w[447:440] : dat_pre_data[447:440];
  assign _01092_ = _05481_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29626" *) dat_pre_data_w[439:432] : dat_pre_data[439:432];
  assign _01091_ = _05480_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29616" *) dat_pre_data_w[431:424] : dat_pre_data[431:424];
  assign _01090_ = _05479_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29606" *) dat_pre_data_w[423:416] : dat_pre_data[423:416];
  assign _01089_ = _05478_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29596" *) dat_pre_data_w[415:408] : dat_pre_data[415:408];
  assign _01088_ = _05477_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29586" *) dat_pre_data_w[407:400] : dat_pre_data[407:400];
  assign _01086_ = _05476_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29576" *) dat_pre_data_w[399:392] : dat_pre_data[399:392];
  assign _01085_ = _05475_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29566" *) dat_pre_data_w[391:384] : dat_pre_data[391:384];
  assign _01084_ = _05474_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29556" *) dat_pre_data_w[383:376] : dat_pre_data[383:376];
  assign _01083_ = _05473_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29546" *) dat_pre_data_w[375:368] : dat_pre_data[375:368];
  assign _01082_ = _05472_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29536" *) dat_pre_data_w[367:360] : dat_pre_data[367:360];
  assign _01081_ = _05471_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29526" *) dat_pre_data_w[359:352] : dat_pre_data[359:352];
  assign _01080_ = _05470_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29516" *) dat_pre_data_w[351:344] : dat_pre_data[351:344];
  assign _01079_ = _05469_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29506" *) dat_pre_data_w[343:336] : dat_pre_data[343:336];
  assign _01078_ = _05468_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29496" *) dat_pre_data_w[335:328] : dat_pre_data[335:328];
  assign _01077_ = _05467_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29486" *) dat_pre_data_w[327:320] : dat_pre_data[327:320];
  assign _01075_ = _05466_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29476" *) dat_pre_data_w[319:312] : dat_pre_data[319:312];
  assign _01074_ = _05465_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29466" *) dat_pre_data_w[311:304] : dat_pre_data[311:304];
  assign _01073_ = _05464_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29456" *) dat_pre_data_w[303:296] : dat_pre_data[303:296];
  assign _01072_ = _05463_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29446" *) dat_pre_data_w[295:288] : dat_pre_data[295:288];
  assign _01071_ = _05462_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29436" *) dat_pre_data_w[287:280] : dat_pre_data[287:280];
  assign _01070_ = _05461_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29426" *) dat_pre_data_w[279:272] : dat_pre_data[279:272];
  assign _01069_ = _05460_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29416" *) dat_pre_data_w[271:264] : dat_pre_data[271:264];
  assign _01068_ = _05459_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29406" *) dat_pre_data_w[263:256] : dat_pre_data[263:256];
  assign _01067_ = _05458_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29396" *) dat_pre_data_w[255:248] : dat_pre_data[255:248];
  assign _01066_ = _05457_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29386" *) dat_pre_data_w[247:240] : dat_pre_data[247:240];
  assign _01064_ = _05456_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29376" *) dat_pre_data_w[239:232] : dat_pre_data[239:232];
  assign _01063_ = _05455_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29366" *) dat_pre_data_w[231:224] : dat_pre_data[231:224];
  assign _01062_ = _05454_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29356" *) dat_pre_data_w[223:216] : dat_pre_data[223:216];
  assign _01061_ = _05453_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29346" *) dat_pre_data_w[215:208] : dat_pre_data[215:208];
  assign _01060_ = _05452_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29336" *) dat_pre_data_w[207:200] : dat_pre_data[207:200];
  assign _01059_ = _05451_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29326" *) dat_pre_data_w[199:192] : dat_pre_data[199:192];
  assign _01058_ = _05450_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29316" *) dat_pre_data_w[191:184] : dat_pre_data[191:184];
  assign _01057_ = _05449_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29306" *) dat_pre_data_w[183:176] : dat_pre_data[183:176];
  assign _01056_ = _05448_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29296" *) dat_pre_data_w[175:168] : dat_pre_data[175:168];
  assign _01055_ = _05447_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29286" *) dat_pre_data_w[167:160] : dat_pre_data[167:160];
  assign _01053_ = _05446_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29276" *) dat_pre_data_w[159:152] : dat_pre_data[159:152];
  assign _01052_ = _05445_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29266" *) dat_pre_data_w[151:144] : dat_pre_data[151:144];
  assign _01051_ = _05444_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29256" *) dat_pre_data_w[143:136] : dat_pre_data[143:136];
  assign _01050_ = _05443_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29246" *) dat_pre_data_w[135:128] : dat_pre_data[135:128];
  assign _01049_ = _05442_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29236" *) dat_pre_data_w[127:120] : dat_pre_data[127:120];
  assign _01048_ = _05441_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29226" *) dat_pre_data_w[119:112] : dat_pre_data[119:112];
  assign _01047_ = _05440_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29216" *) dat_pre_data_w[111:104] : dat_pre_data[111:104];
  assign _01046_ = _05439_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29206" *) dat_pre_data_w[103:96] : dat_pre_data[103:96];
  assign _01165_ = _05438_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29196" *) dat_pre_data_w[95:88] : dat_pre_data[95:88];
  assign _01154_ = _05437_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29186" *) dat_pre_data_w[87:80] : dat_pre_data[87:80];
  assign _01142_ = _05436_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29176" *) dat_pre_data_w[79:72] : dat_pre_data[79:72];
  assign _01131_ = _05435_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29166" *) dat_pre_data_w[71:64] : dat_pre_data[71:64];
  assign _01120_ = _05434_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29156" *) dat_pre_data_w[63:56] : dat_pre_data[63:56];
  assign _01109_ = _05433_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29146" *) dat_pre_data_w[55:48] : dat_pre_data[55:48];
  assign _01098_ = _05432_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29136" *) dat_pre_data_w[47:40] : dat_pre_data[47:40];
  assign _01087_ = _05431_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29126" *) dat_pre_data_w[39:32] : dat_pre_data[39:32];
  assign _01076_ = _05430_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29116" *) dat_pre_data_w[31:24] : dat_pre_data[31:24];
  assign _01065_ = _05429_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29106" *) dat_pre_data_w[23:16] : dat_pre_data[23:16];
  assign _01054_ = _05428_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29096" *) dat_pre_data_w[15:8] : dat_pre_data[15:8];
  assign _01143_ = _05427_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29086" *) dat_pre_data_w[7:0] : dat_pre_data[7:0];
  assign _01187_ = _05426_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29076" *) in_dat_nan : dat_pre_nan;
  assign _01188_ = in_dat_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29066" *) dat_pre_nz_w : dat_pre_nz;
  assign _03027_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26586" *) _05169_ : wt7_actv_data[1023:1016];
  assign _03026_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26576" *) _05167_ : wt7_actv_data[1015:1008];
  assign _03025_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26566" *) _05166_ : wt7_actv_data[1007:1000];
  assign _03152_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26556" *) _05165_ : wt7_actv_data[999:992];
  assign _03151_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26546" *) _05164_ : wt7_actv_data[991:984];
  assign _03150_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26536" *) _05163_ : wt7_actv_data[983:976];
  assign _03149_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26526" *) _05162_ : wt7_actv_data[975:968];
  assign _03148_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26516" *) _05161_ : wt7_actv_data[967:960];
  assign _03146_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26506" *) _05158_ : wt7_actv_data[959:952];
  assign _03145_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26496" *) _05155_ : wt7_actv_data[951:944];
  assign _03144_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26486" *) _05152_ : wt7_actv_data[943:936];
  assign _03143_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26476" *) _05149_ : wt7_actv_data[935:928];
  assign _03142_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26466" *) _05146_ : wt7_actv_data[927:920];
  assign _03141_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26456" *) _05143_ : wt7_actv_data[919:912];
  assign _03140_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26446" *) _05140_ : wt7_actv_data[911:904];
  assign _03139_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26436" *) _05137_ : wt7_actv_data[903:896];
  assign _03138_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26426" *) _05134_ : wt7_actv_data[895:888];
  assign _03137_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26416" *) _05131_ : wt7_actv_data[887:880];
  assign _03135_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26406" *) _05128_ : wt7_actv_data[879:872];
  assign _03134_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26396" *) _05125_ : wt7_actv_data[871:864];
  assign _03133_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26386" *) _05122_ : wt7_actv_data[863:856];
  assign _03132_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26376" *) _05119_ : wt7_actv_data[855:848];
  assign _03131_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26366" *) _05116_ : wt7_actv_data[847:840];
  assign _03130_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26356" *) _05113_ : wt7_actv_data[839:832];
  assign _03129_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26346" *) _05110_ : wt7_actv_data[831:824];
  assign _03128_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26336" *) _05107_ : wt7_actv_data[823:816];
  assign _03127_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26326" *) _05104_ : wt7_actv_data[815:808];
  assign _03126_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26316" *) _05101_ : wt7_actv_data[807:800];
  assign _03123_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26306" *) _05098_ : wt7_actv_data[799:792];
  assign _03122_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26296" *) _05095_ : wt7_actv_data[791:784];
  assign _03121_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26286" *) _05092_ : wt7_actv_data[783:776];
  assign _03120_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26276" *) _05089_ : wt7_actv_data[775:768];
  assign _03119_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26266" *) _05086_ : wt7_actv_data[767:760];
  assign _03118_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26256" *) _05083_ : wt7_actv_data[759:752];
  assign _03117_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26246" *) _05080_ : wt7_actv_data[751:744];
  assign _03116_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26236" *) _05077_ : wt7_actv_data[743:736];
  assign _03115_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26226" *) _05074_ : wt7_actv_data[735:728];
  assign _03114_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26216" *) _05071_ : wt7_actv_data[727:720];
  assign _03112_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26206" *) _05068_ : wt7_actv_data[719:712];
  assign _03111_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26196" *) _05065_ : wt7_actv_data[711:704];
  assign _03110_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26186" *) _05062_ : wt7_actv_data[703:696];
  assign _03109_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26176" *) _05059_ : wt7_actv_data[695:688];
  assign _03108_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26166" *) _05056_ : wt7_actv_data[687:680];
  assign _03107_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26156" *) _05053_ : wt7_actv_data[679:672];
  assign _03106_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26146" *) _05050_ : wt7_actv_data[671:664];
  assign _03105_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26136" *) _05047_ : wt7_actv_data[663:656];
  assign _03104_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26126" *) _05044_ : wt7_actv_data[655:648];
  assign _03103_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26116" *) _05041_ : wt7_actv_data[647:640];
  assign _03101_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26106" *) _05038_ : wt7_actv_data[639:632];
  assign _03100_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26096" *) _05035_ : wt7_actv_data[631:624];
  assign _03099_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26086" *) _05032_ : wt7_actv_data[623:616];
  assign _03098_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26076" *) _05029_ : wt7_actv_data[615:608];
  assign _03097_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26066" *) _05026_ : wt7_actv_data[607:600];
  assign _03096_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26056" *) _05023_ : wt7_actv_data[599:592];
  assign _03095_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26046" *) _05020_ : wt7_actv_data[591:584];
  assign _03094_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26036" *) _05017_ : wt7_actv_data[583:576];
  assign _03093_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26026" *) _05014_ : wt7_actv_data[575:568];
  assign _03092_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26016" *) _05011_ : wt7_actv_data[567:560];
  assign _03090_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:26006" *) _05008_ : wt7_actv_data[559:552];
  assign _03089_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25996" *) _05005_ : wt7_actv_data[551:544];
  assign _03088_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25986" *) _05002_ : wt7_actv_data[543:536];
  assign _03087_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25976" *) _04999_ : wt7_actv_data[535:528];
  assign _03086_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25966" *) _04996_ : wt7_actv_data[527:520];
  assign _03085_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25956" *) _04993_ : wt7_actv_data[519:512];
  assign _03084_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25946" *) _04990_ : wt7_actv_data[511:504];
  assign _03083_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25936" *) _04987_ : wt7_actv_data[503:496];
  assign _03082_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25926" *) _04984_ : wt7_actv_data[495:488];
  assign _03081_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25916" *) _04981_ : wt7_actv_data[487:480];
  assign _03079_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25906" *) _04978_ : wt7_actv_data[479:472];
  assign _03078_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25896" *) _04975_ : wt7_actv_data[471:464];
  assign _03077_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25886" *) _04972_ : wt7_actv_data[463:456];
  assign _03076_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25876" *) _04969_ : wt7_actv_data[455:448];
  assign _03075_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25866" *) _04968_ : wt7_actv_data[447:440];
  assign _03074_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25856" *) _04967_ : wt7_actv_data[439:432];
  assign _03073_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25846" *) _04966_ : wt7_actv_data[431:424];
  assign _03072_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25836" *) _04965_ : wt7_actv_data[423:416];
  assign _03071_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25826" *) _04964_ : wt7_actv_data[415:408];
  assign _03070_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25816" *) _04963_ : wt7_actv_data[407:400];
  assign _03068_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25806" *) _04962_ : wt7_actv_data[399:392];
  assign _03067_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25796" *) _04961_ : wt7_actv_data[391:384];
  assign _03066_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25786" *) _04960_ : wt7_actv_data[383:376];
  assign _03065_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25776" *) _04959_ : wt7_actv_data[375:368];
  assign _03064_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25766" *) _04958_ : wt7_actv_data[367:360];
  assign _03063_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25756" *) _04957_ : wt7_actv_data[359:352];
  assign _03062_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25746" *) _04956_ : wt7_actv_data[351:344];
  assign _03061_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25736" *) _04955_ : wt7_actv_data[343:336];
  assign _03060_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25726" *) _04954_ : wt7_actv_data[335:328];
  assign _03059_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25716" *) _04953_ : wt7_actv_data[327:320];
  assign _03057_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25706" *) _04952_ : wt7_actv_data[319:312];
  assign _03056_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25696" *) _04951_ : wt7_actv_data[311:304];
  assign _03055_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25686" *) _04950_ : wt7_actv_data[303:296];
  assign _03054_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25676" *) _04949_ : wt7_actv_data[295:288];
  assign _03053_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25666" *) _04948_ : wt7_actv_data[287:280];
  assign _03052_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25656" *) _04947_ : wt7_actv_data[279:272];
  assign _03051_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25646" *) _04946_ : wt7_actv_data[271:264];
  assign _03050_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25636" *) _04945_ : wt7_actv_data[263:256];
  assign _03049_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25626" *) _04944_ : wt7_actv_data[255:248];
  assign _03048_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25616" *) _04943_ : wt7_actv_data[247:240];
  assign _03046_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25606" *) _04942_ : wt7_actv_data[239:232];
  assign _03045_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25596" *) _04941_ : wt7_actv_data[231:224];
  assign _03044_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25586" *) _04940_ : wt7_actv_data[223:216];
  assign _03043_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25576" *) _04939_ : wt7_actv_data[215:208];
  assign _03042_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25566" *) _04938_ : wt7_actv_data[207:200];
  assign _03041_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25556" *) _04937_ : wt7_actv_data[199:192];
  assign _03040_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25546" *) _04936_ : wt7_actv_data[191:184];
  assign _03039_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25536" *) _04935_ : wt7_actv_data[183:176];
  assign _03038_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25526" *) _04934_ : wt7_actv_data[175:168];
  assign _03037_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25516" *) _04933_ : wt7_actv_data[167:160];
  assign _03035_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25506" *) _04932_ : wt7_actv_data[159:152];
  assign _03034_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25496" *) _04931_ : wt7_actv_data[151:144];
  assign _03033_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25486" *) _04930_ : wt7_actv_data[143:136];
  assign _03032_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25476" *) _04929_ : wt7_actv_data[135:128];
  assign _03031_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25466" *) _04928_ : wt7_actv_data[127:120];
  assign _03030_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25456" *) _04927_ : wt7_actv_data[119:112];
  assign _03029_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25446" *) _04926_ : wt7_actv_data[111:104];
  assign _03028_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25436" *) _04925_ : wt7_actv_data[103:96];
  assign _03147_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25426" *) _04924_ : wt7_actv_data[95:88];
  assign _03136_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25416" *) _04923_ : wt7_actv_data[87:80];
  assign _03124_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25406" *) _04922_ : wt7_actv_data[79:72];
  assign _03113_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25396" *) _04921_ : wt7_actv_data[71:64];
  assign _03102_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25386" *) _04920_ : wt7_actv_data[63:56];
  assign _03091_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25376" *) _04919_ : wt7_actv_data[55:48];
  assign _03080_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25366" *) _04918_ : wt7_actv_data[47:40];
  assign _03069_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25356" *) _04917_ : wt7_actv_data[39:32];
  assign _03058_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25346" *) _04916_ : wt7_actv_data[31:24];
  assign _03047_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25336" *) _04915_ : wt7_actv_data[23:16];
  assign _03036_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25326" *) _04914_ : wt7_actv_data[15:8];
  assign _03125_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25316" *) _04913_ : wt7_actv_data[7:0];
  assign _03153_ = _04912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25306" *) wt7_sd_nan : wt7_actv_nan;
  assign _03154_ = _04911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25296" *) wt7_sd_nz : wt7_actv_nz;
  assign _02765_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25262" *) _04910_ : wt6_actv_data[1023:1016];
  assign _02764_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25252" *) _04909_ : wt6_actv_data[1015:1008];
  assign _02763_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25242" *) _04908_ : wt6_actv_data[1007:1000];
  assign _02890_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25232" *) _04907_ : wt6_actv_data[999:992];
  assign _02889_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25222" *) _04906_ : wt6_actv_data[991:984];
  assign _02888_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25212" *) _04905_ : wt6_actv_data[983:976];
  assign _02887_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25202" *) _04904_ : wt6_actv_data[975:968];
  assign _02886_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25192" *) _04903_ : wt6_actv_data[967:960];
  assign _02884_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25182" *) _04902_ : wt6_actv_data[959:952];
  assign _02883_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25172" *) _04901_ : wt6_actv_data[951:944];
  assign _02882_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25162" *) _04900_ : wt6_actv_data[943:936];
  assign _02881_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25152" *) _04899_ : wt6_actv_data[935:928];
  assign _02880_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25142" *) _04898_ : wt6_actv_data[927:920];
  assign _02879_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25132" *) _04897_ : wt6_actv_data[919:912];
  assign _02878_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25122" *) _04896_ : wt6_actv_data[911:904];
  assign _02877_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25112" *) _04895_ : wt6_actv_data[903:896];
  assign _02876_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25102" *) _04894_ : wt6_actv_data[895:888];
  assign _02875_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25092" *) _04893_ : wt6_actv_data[887:880];
  assign _02873_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25082" *) _04892_ : wt6_actv_data[879:872];
  assign _02872_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25072" *) _04891_ : wt6_actv_data[871:864];
  assign _02871_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25062" *) _04890_ : wt6_actv_data[863:856];
  assign _02870_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25052" *) _04889_ : wt6_actv_data[855:848];
  assign _02869_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25042" *) _04888_ : wt6_actv_data[847:840];
  assign _02868_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25032" *) _04887_ : wt6_actv_data[839:832];
  assign _02867_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25022" *) _04886_ : wt6_actv_data[831:824];
  assign _02866_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25012" *) _04885_ : wt6_actv_data[823:816];
  assign _02865_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25002" *) _04884_ : wt6_actv_data[815:808];
  assign _02864_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24992" *) _04883_ : wt6_actv_data[807:800];
  assign _02861_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24982" *) _04882_ : wt6_actv_data[799:792];
  assign _02860_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24972" *) _04881_ : wt6_actv_data[791:784];
  assign _02859_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24962" *) _04880_ : wt6_actv_data[783:776];
  assign _02858_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24952" *) _04879_ : wt6_actv_data[775:768];
  assign _02857_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24942" *) _04878_ : wt6_actv_data[767:760];
  assign _02856_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24932" *) _04877_ : wt6_actv_data[759:752];
  assign _02855_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24922" *) _04876_ : wt6_actv_data[751:744];
  assign _02854_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24912" *) _04875_ : wt6_actv_data[743:736];
  assign _02853_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24902" *) _04874_ : wt6_actv_data[735:728];
  assign _02852_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24892" *) _04873_ : wt6_actv_data[727:720];
  assign _02850_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24882" *) _04872_ : wt6_actv_data[719:712];
  assign _02849_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24872" *) _04871_ : wt6_actv_data[711:704];
  assign _02848_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24862" *) _04870_ : wt6_actv_data[703:696];
  assign _02847_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24852" *) _04869_ : wt6_actv_data[695:688];
  assign _02846_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24842" *) _04868_ : wt6_actv_data[687:680];
  assign _02845_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24832" *) _04867_ : wt6_actv_data[679:672];
  assign _02844_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24822" *) _04866_ : wt6_actv_data[671:664];
  assign _02843_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24812" *) _04865_ : wt6_actv_data[663:656];
  assign _02842_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24802" *) _04864_ : wt6_actv_data[655:648];
  assign _02841_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24792" *) _04863_ : wt6_actv_data[647:640];
  assign _02839_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24782" *) _04862_ : wt6_actv_data[639:632];
  assign _02838_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24772" *) _04861_ : wt6_actv_data[631:624];
  assign _02837_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24762" *) _04860_ : wt6_actv_data[623:616];
  assign _02836_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24752" *) _04859_ : wt6_actv_data[615:608];
  assign _02835_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24742" *) _04858_ : wt6_actv_data[607:600];
  assign _02834_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24732" *) _04857_ : wt6_actv_data[599:592];
  assign _02833_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24722" *) _04856_ : wt6_actv_data[591:584];
  assign _02832_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24712" *) _04855_ : wt6_actv_data[583:576];
  assign _02831_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24702" *) _04854_ : wt6_actv_data[575:568];
  assign _02830_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24692" *) _04853_ : wt6_actv_data[567:560];
  assign _02828_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24682" *) _04852_ : wt6_actv_data[559:552];
  assign _02827_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24672" *) _04851_ : wt6_actv_data[551:544];
  assign _02826_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24662" *) _04850_ : wt6_actv_data[543:536];
  assign _02825_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24652" *) _04849_ : wt6_actv_data[535:528];
  assign _02824_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24642" *) _04848_ : wt6_actv_data[527:520];
  assign _02823_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24632" *) _04847_ : wt6_actv_data[519:512];
  assign _02822_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24622" *) _04846_ : wt6_actv_data[511:504];
  assign _02821_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24612" *) _04845_ : wt6_actv_data[503:496];
  assign _02820_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24602" *) _04844_ : wt6_actv_data[495:488];
  assign _02819_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24592" *) _04843_ : wt6_actv_data[487:480];
  assign _02817_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24582" *) _04842_ : wt6_actv_data[479:472];
  assign _02816_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24572" *) _04841_ : wt6_actv_data[471:464];
  assign _02815_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24562" *) _04840_ : wt6_actv_data[463:456];
  assign _02814_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24552" *) _04839_ : wt6_actv_data[455:448];
  assign _02813_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24542" *) _04838_ : wt6_actv_data[447:440];
  assign _02812_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24532" *) _04837_ : wt6_actv_data[439:432];
  assign _02811_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24522" *) _04836_ : wt6_actv_data[431:424];
  assign _02810_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24512" *) _04835_ : wt6_actv_data[423:416];
  assign _02809_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24502" *) _04834_ : wt6_actv_data[415:408];
  assign _02808_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24492" *) _04833_ : wt6_actv_data[407:400];
  assign _02806_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24482" *) _04832_ : wt6_actv_data[399:392];
  assign _02805_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24472" *) _04831_ : wt6_actv_data[391:384];
  assign _02804_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24462" *) _04830_ : wt6_actv_data[383:376];
  assign _02803_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24452" *) _04829_ : wt6_actv_data[375:368];
  assign _02802_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24442" *) _04828_ : wt6_actv_data[367:360];
  assign _02801_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24432" *) _04827_ : wt6_actv_data[359:352];
  assign _02800_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24422" *) _04826_ : wt6_actv_data[351:344];
  assign _02799_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24412" *) _04825_ : wt6_actv_data[343:336];
  assign _02798_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24402" *) _04824_ : wt6_actv_data[335:328];
  assign _02797_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24392" *) _04823_ : wt6_actv_data[327:320];
  assign _02795_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24382" *) _04822_ : wt6_actv_data[319:312];
  assign _02794_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24372" *) _04821_ : wt6_actv_data[311:304];
  assign _02793_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24362" *) _04820_ : wt6_actv_data[303:296];
  assign _02792_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24352" *) _04819_ : wt6_actv_data[295:288];
  assign _02791_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24342" *) _04818_ : wt6_actv_data[287:280];
  assign _02790_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24332" *) _04817_ : wt6_actv_data[279:272];
  assign _02789_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24322" *) _04816_ : wt6_actv_data[271:264];
  assign _02788_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24312" *) _04815_ : wt6_actv_data[263:256];
  assign _02787_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24302" *) _04814_ : wt6_actv_data[255:248];
  assign _02786_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24292" *) _04813_ : wt6_actv_data[247:240];
  assign _02784_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24282" *) _04812_ : wt6_actv_data[239:232];
  assign _02783_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24272" *) _04811_ : wt6_actv_data[231:224];
  assign _02782_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24262" *) _04810_ : wt6_actv_data[223:216];
  assign _02781_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24252" *) _04809_ : wt6_actv_data[215:208];
  assign _02780_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24242" *) _04808_ : wt6_actv_data[207:200];
  assign _02779_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24232" *) _04807_ : wt6_actv_data[199:192];
  assign _02778_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24222" *) _04806_ : wt6_actv_data[191:184];
  assign _02777_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24212" *) _04805_ : wt6_actv_data[183:176];
  assign _02776_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24202" *) _04804_ : wt6_actv_data[175:168];
  assign _02775_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24192" *) _04803_ : wt6_actv_data[167:160];
  assign _02773_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24182" *) _04802_ : wt6_actv_data[159:152];
  assign _02772_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24172" *) _04801_ : wt6_actv_data[151:144];
  assign _02771_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24162" *) _04800_ : wt6_actv_data[143:136];
  assign _02770_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24152" *) _04799_ : wt6_actv_data[135:128];
  assign _02769_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24142" *) _04798_ : wt6_actv_data[127:120];
  assign _02768_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24132" *) _04797_ : wt6_actv_data[119:112];
  assign _02767_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24122" *) _04796_ : wt6_actv_data[111:104];
  assign _02766_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24112" *) _04795_ : wt6_actv_data[103:96];
  assign _02885_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24102" *) _04794_ : wt6_actv_data[95:88];
  assign _02874_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24092" *) _04793_ : wt6_actv_data[87:80];
  assign _02862_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24082" *) _04792_ : wt6_actv_data[79:72];
  assign _02851_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24072" *) _04791_ : wt6_actv_data[71:64];
  assign _02840_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24062" *) _04790_ : wt6_actv_data[63:56];
  assign _02829_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24052" *) _04789_ : wt6_actv_data[55:48];
  assign _02818_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24042" *) _04788_ : wt6_actv_data[47:40];
  assign _02807_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24032" *) _04787_ : wt6_actv_data[39:32];
  assign _02796_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24022" *) _04786_ : wt6_actv_data[31:24];
  assign _02785_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24012" *) _04785_ : wt6_actv_data[23:16];
  assign _02774_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:24002" *) _04784_ : wt6_actv_data[15:8];
  assign _02863_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23992" *) _04783_ : wt6_actv_data[7:0];
  assign _02891_ = _04782_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23982" *) wt6_sd_nan : wt6_actv_nan;
  assign _02892_ = _04781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23972" *) wt6_sd_nz : wt6_actv_nz;
  assign _02503_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23938" *) _04780_ : wt5_actv_data[1023:1016];
  assign _02502_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23928" *) _04779_ : wt5_actv_data[1015:1008];
  assign _02501_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23918" *) _04778_ : wt5_actv_data[1007:1000];
  assign _02628_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23908" *) _04777_ : wt5_actv_data[999:992];
  assign _02627_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23898" *) _04776_ : wt5_actv_data[991:984];
  assign _02626_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23888" *) _04775_ : wt5_actv_data[983:976];
  assign _02625_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23878" *) _04774_ : wt5_actv_data[975:968];
  assign _02624_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23868" *) _04773_ : wt5_actv_data[967:960];
  assign _02622_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23858" *) _04772_ : wt5_actv_data[959:952];
  assign _02621_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23848" *) _04771_ : wt5_actv_data[951:944];
  assign _02620_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23838" *) _04770_ : wt5_actv_data[943:936];
  assign _02619_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23828" *) _04769_ : wt5_actv_data[935:928];
  assign _02618_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23818" *) _04768_ : wt5_actv_data[927:920];
  assign _02617_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23808" *) _04767_ : wt5_actv_data[919:912];
  assign _02616_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23798" *) _04766_ : wt5_actv_data[911:904];
  assign _02615_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23788" *) _04765_ : wt5_actv_data[903:896];
  assign _02614_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23778" *) _04764_ : wt5_actv_data[895:888];
  assign _02613_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23768" *) _04763_ : wt5_actv_data[887:880];
  assign _02611_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23758" *) _04762_ : wt5_actv_data[879:872];
  assign _02610_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23748" *) _04761_ : wt5_actv_data[871:864];
  assign _02609_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23738" *) _04760_ : wt5_actv_data[863:856];
  assign _02608_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23728" *) _04759_ : wt5_actv_data[855:848];
  assign _02607_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23718" *) _04758_ : wt5_actv_data[847:840];
  assign _02606_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23708" *) _04757_ : wt5_actv_data[839:832];
  assign _02605_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23698" *) _04756_ : wt5_actv_data[831:824];
  assign _02604_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23688" *) _04755_ : wt5_actv_data[823:816];
  assign _02603_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23678" *) _04754_ : wt5_actv_data[815:808];
  assign _02602_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23668" *) _04753_ : wt5_actv_data[807:800];
  assign _02599_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23658" *) _04752_ : wt5_actv_data[799:792];
  assign _02598_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23648" *) _04751_ : wt5_actv_data[791:784];
  assign _02597_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23638" *) _04750_ : wt5_actv_data[783:776];
  assign _02596_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23628" *) _04749_ : wt5_actv_data[775:768];
  assign _02595_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23618" *) _04748_ : wt5_actv_data[767:760];
  assign _02594_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23608" *) _04747_ : wt5_actv_data[759:752];
  assign _02593_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23598" *) _04746_ : wt5_actv_data[751:744];
  assign _02592_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23588" *) _04745_ : wt5_actv_data[743:736];
  assign _02591_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23578" *) _04744_ : wt5_actv_data[735:728];
  assign _02590_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23568" *) _04743_ : wt5_actv_data[727:720];
  assign _02588_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23558" *) _04742_ : wt5_actv_data[719:712];
  assign _02587_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23548" *) _04741_ : wt5_actv_data[711:704];
  assign _02586_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23538" *) _04740_ : wt5_actv_data[703:696];
  assign _02585_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23528" *) _04739_ : wt5_actv_data[695:688];
  assign _02584_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23518" *) _04738_ : wt5_actv_data[687:680];
  assign _02583_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23508" *) _04737_ : wt5_actv_data[679:672];
  assign _02582_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23498" *) _04736_ : wt5_actv_data[671:664];
  assign _02581_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23488" *) _04735_ : wt5_actv_data[663:656];
  assign _02580_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23478" *) _04734_ : wt5_actv_data[655:648];
  assign _02579_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23468" *) _04733_ : wt5_actv_data[647:640];
  assign _02577_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23458" *) _04732_ : wt5_actv_data[639:632];
  assign _02576_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23448" *) _04731_ : wt5_actv_data[631:624];
  assign _02575_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23438" *) _04730_ : wt5_actv_data[623:616];
  assign _02574_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23428" *) _04729_ : wt5_actv_data[615:608];
  assign _02573_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23418" *) _04728_ : wt5_actv_data[607:600];
  assign _02572_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23408" *) _04727_ : wt5_actv_data[599:592];
  assign _02571_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23398" *) _04726_ : wt5_actv_data[591:584];
  assign _02570_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23388" *) _04725_ : wt5_actv_data[583:576];
  assign _02569_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23378" *) _04724_ : wt5_actv_data[575:568];
  assign _02568_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23368" *) _04723_ : wt5_actv_data[567:560];
  assign _02566_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23358" *) _04722_ : wt5_actv_data[559:552];
  assign _02565_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23348" *) _04721_ : wt5_actv_data[551:544];
  assign _02564_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23338" *) _04720_ : wt5_actv_data[543:536];
  assign _02563_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23328" *) _04719_ : wt5_actv_data[535:528];
  assign _02562_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23318" *) _04718_ : wt5_actv_data[527:520];
  assign _02561_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23308" *) _04717_ : wt5_actv_data[519:512];
  assign _02560_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23298" *) _04716_ : wt5_actv_data[511:504];
  assign _02559_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23288" *) _04715_ : wt5_actv_data[503:496];
  assign _02558_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23278" *) _04714_ : wt5_actv_data[495:488];
  assign _02557_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23268" *) _04713_ : wt5_actv_data[487:480];
  assign _02555_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23258" *) _04712_ : wt5_actv_data[479:472];
  assign _02554_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23248" *) _04711_ : wt5_actv_data[471:464];
  assign _02553_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23238" *) _04710_ : wt5_actv_data[463:456];
  assign _02552_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23228" *) _04709_ : wt5_actv_data[455:448];
  assign _02551_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23218" *) _04708_ : wt5_actv_data[447:440];
  assign _02550_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23208" *) _04707_ : wt5_actv_data[439:432];
  assign _02549_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23198" *) _04706_ : wt5_actv_data[431:424];
  assign _02548_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23188" *) _04705_ : wt5_actv_data[423:416];
  assign _02547_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23178" *) _04704_ : wt5_actv_data[415:408];
  assign _02546_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23168" *) _04703_ : wt5_actv_data[407:400];
  assign _02544_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23158" *) _04702_ : wt5_actv_data[399:392];
  assign _02543_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23148" *) _04701_ : wt5_actv_data[391:384];
  assign _02542_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23138" *) _04700_ : wt5_actv_data[383:376];
  assign _02541_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23128" *) _04699_ : wt5_actv_data[375:368];
  assign _02540_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23118" *) _04698_ : wt5_actv_data[367:360];
  assign _02539_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23108" *) _04697_ : wt5_actv_data[359:352];
  assign _02538_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23098" *) _04696_ : wt5_actv_data[351:344];
  assign _02537_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23088" *) _04695_ : wt5_actv_data[343:336];
  assign _02536_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23078" *) _04694_ : wt5_actv_data[335:328];
  assign _02535_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23068" *) _04693_ : wt5_actv_data[327:320];
  assign _02533_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23058" *) _04692_ : wt5_actv_data[319:312];
  assign _02532_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23048" *) _04691_ : wt5_actv_data[311:304];
  assign _02531_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23038" *) _04690_ : wt5_actv_data[303:296];
  assign _02530_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23028" *) _04689_ : wt5_actv_data[295:288];
  assign _02529_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23018" *) _04688_ : wt5_actv_data[287:280];
  assign _02528_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23008" *) _04687_ : wt5_actv_data[279:272];
  assign _02527_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22998" *) _04686_ : wt5_actv_data[271:264];
  assign _02526_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22988" *) _04685_ : wt5_actv_data[263:256];
  assign _02525_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22978" *) _04684_ : wt5_actv_data[255:248];
  assign _02524_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22968" *) _04683_ : wt5_actv_data[247:240];
  assign _02522_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22958" *) _04682_ : wt5_actv_data[239:232];
  assign _02521_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22948" *) _04681_ : wt5_actv_data[231:224];
  assign _02520_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22938" *) _04680_ : wt5_actv_data[223:216];
  assign _02519_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22928" *) _04679_ : wt5_actv_data[215:208];
  assign _02518_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22918" *) _04678_ : wt5_actv_data[207:200];
  assign _02517_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22908" *) _04677_ : wt5_actv_data[199:192];
  assign _02516_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22898" *) _04676_ : wt5_actv_data[191:184];
  assign _02515_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22888" *) _04675_ : wt5_actv_data[183:176];
  assign _02514_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22878" *) _04674_ : wt5_actv_data[175:168];
  assign _02513_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22868" *) _04673_ : wt5_actv_data[167:160];
  assign _02511_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22858" *) _04672_ : wt5_actv_data[159:152];
  assign _02510_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22848" *) _04671_ : wt5_actv_data[151:144];
  assign _02509_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22838" *) _04670_ : wt5_actv_data[143:136];
  assign _02508_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22828" *) _04669_ : wt5_actv_data[135:128];
  assign _02507_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22818" *) _04668_ : wt5_actv_data[127:120];
  assign _02506_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22808" *) _04667_ : wt5_actv_data[119:112];
  assign _02505_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22798" *) _04666_ : wt5_actv_data[111:104];
  assign _02504_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22788" *) _04665_ : wt5_actv_data[103:96];
  assign _02623_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22778" *) _04664_ : wt5_actv_data[95:88];
  assign _02612_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22768" *) _04663_ : wt5_actv_data[87:80];
  assign _02600_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22758" *) _04662_ : wt5_actv_data[79:72];
  assign _02589_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22748" *) _04661_ : wt5_actv_data[71:64];
  assign _02578_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22738" *) _04660_ : wt5_actv_data[63:56];
  assign _02567_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22728" *) _04659_ : wt5_actv_data[55:48];
  assign _02556_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22718" *) _04658_ : wt5_actv_data[47:40];
  assign _02545_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22708" *) _04657_ : wt5_actv_data[39:32];
  assign _02534_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22698" *) _04656_ : wt5_actv_data[31:24];
  assign _02523_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22688" *) _04655_ : wt5_actv_data[23:16];
  assign _02512_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22678" *) _04654_ : wt5_actv_data[15:8];
  assign _02601_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22668" *) _04653_ : wt5_actv_data[7:0];
  assign _02629_ = _04652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22658" *) wt5_sd_nan : wt5_actv_nan;
  assign _02630_ = _04651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22648" *) wt5_sd_nz : wt5_actv_nz;
  assign _02241_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22614" *) _04650_ : wt4_actv_data[1023:1016];
  assign _02240_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22604" *) _04649_ : wt4_actv_data[1015:1008];
  assign _02239_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22594" *) _04648_ : wt4_actv_data[1007:1000];
  assign _02366_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22584" *) _04647_ : wt4_actv_data[999:992];
  assign _02365_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22574" *) _04646_ : wt4_actv_data[991:984];
  assign _02364_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22564" *) _04645_ : wt4_actv_data[983:976];
  assign _02363_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22554" *) _04644_ : wt4_actv_data[975:968];
  assign _02362_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22544" *) _04643_ : wt4_actv_data[967:960];
  assign _02360_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22534" *) _04642_ : wt4_actv_data[959:952];
  assign _02359_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22524" *) _04641_ : wt4_actv_data[951:944];
  assign _02358_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22514" *) _04640_ : wt4_actv_data[943:936];
  assign _02357_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22504" *) _04639_ : wt4_actv_data[935:928];
  assign _02356_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22494" *) _04638_ : wt4_actv_data[927:920];
  assign _02355_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22484" *) _04637_ : wt4_actv_data[919:912];
  assign _02354_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22474" *) _04636_ : wt4_actv_data[911:904];
  assign _02353_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22464" *) _04635_ : wt4_actv_data[903:896];
  assign _02352_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22454" *) _04634_ : wt4_actv_data[895:888];
  assign _02351_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22444" *) _04633_ : wt4_actv_data[887:880];
  assign _02349_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22434" *) _04632_ : wt4_actv_data[879:872];
  assign _02348_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22424" *) _04631_ : wt4_actv_data[871:864];
  assign _02347_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22414" *) _04630_ : wt4_actv_data[863:856];
  assign _02346_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22404" *) _04629_ : wt4_actv_data[855:848];
  assign _02345_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22394" *) _04628_ : wt4_actv_data[847:840];
  assign _02344_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22384" *) _04627_ : wt4_actv_data[839:832];
  assign _02343_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22374" *) _04626_ : wt4_actv_data[831:824];
  assign _02342_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22364" *) _04625_ : wt4_actv_data[823:816];
  assign _02341_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22354" *) _04624_ : wt4_actv_data[815:808];
  assign _02340_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22344" *) _04623_ : wt4_actv_data[807:800];
  assign _02337_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22334" *) _04622_ : wt4_actv_data[799:792];
  assign _02336_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22324" *) _04621_ : wt4_actv_data[791:784];
  assign _02335_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22314" *) _04620_ : wt4_actv_data[783:776];
  assign _02334_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22304" *) _04619_ : wt4_actv_data[775:768];
  assign _02333_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22294" *) _04618_ : wt4_actv_data[767:760];
  assign _02332_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22284" *) _04617_ : wt4_actv_data[759:752];
  assign _02331_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22274" *) _04616_ : wt4_actv_data[751:744];
  assign _02330_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22264" *) _04615_ : wt4_actv_data[743:736];
  assign _02329_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22254" *) _04614_ : wt4_actv_data[735:728];
  assign _02328_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22244" *) _04613_ : wt4_actv_data[727:720];
  assign _02326_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22234" *) _04612_ : wt4_actv_data[719:712];
  assign _02325_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22224" *) _04611_ : wt4_actv_data[711:704];
  assign _02324_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22214" *) _04610_ : wt4_actv_data[703:696];
  assign _02323_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22204" *) _04609_ : wt4_actv_data[695:688];
  assign _02322_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22194" *) _04608_ : wt4_actv_data[687:680];
  assign _02321_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22184" *) _04607_ : wt4_actv_data[679:672];
  assign _02320_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22174" *) _04606_ : wt4_actv_data[671:664];
  assign _02319_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22164" *) _04605_ : wt4_actv_data[663:656];
  assign _02318_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22154" *) _04604_ : wt4_actv_data[655:648];
  assign _02317_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22144" *) _04603_ : wt4_actv_data[647:640];
  assign _02315_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22134" *) _04602_ : wt4_actv_data[639:632];
  assign _02314_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22124" *) _04601_ : wt4_actv_data[631:624];
  assign _02313_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22114" *) _04600_ : wt4_actv_data[623:616];
  assign _02312_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22104" *) _04599_ : wt4_actv_data[615:608];
  assign _02311_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22094" *) _04598_ : wt4_actv_data[607:600];
  assign _02310_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22084" *) _04597_ : wt4_actv_data[599:592];
  assign _02309_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22074" *) _04596_ : wt4_actv_data[591:584];
  assign _02308_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22064" *) _04595_ : wt4_actv_data[583:576];
  assign _02307_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22054" *) _04594_ : wt4_actv_data[575:568];
  assign _02306_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22044" *) _04593_ : wt4_actv_data[567:560];
  assign _02304_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22034" *) _04592_ : wt4_actv_data[559:552];
  assign _02303_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22024" *) _04591_ : wt4_actv_data[551:544];
  assign _02302_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22014" *) _04590_ : wt4_actv_data[543:536];
  assign _02301_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22004" *) _04589_ : wt4_actv_data[535:528];
  assign _02300_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21994" *) _04588_ : wt4_actv_data[527:520];
  assign _02299_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21984" *) _04587_ : wt4_actv_data[519:512];
  assign _02298_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21974" *) _04586_ : wt4_actv_data[511:504];
  assign _02297_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21964" *) _04585_ : wt4_actv_data[503:496];
  assign _02296_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21954" *) _04584_ : wt4_actv_data[495:488];
  assign _02295_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21944" *) _04583_ : wt4_actv_data[487:480];
  assign _02293_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21934" *) _04582_ : wt4_actv_data[479:472];
  assign _02292_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21924" *) _04581_ : wt4_actv_data[471:464];
  assign _02291_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21914" *) _04580_ : wt4_actv_data[463:456];
  assign _02290_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21904" *) _04579_ : wt4_actv_data[455:448];
  assign _02289_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21894" *) _04578_ : wt4_actv_data[447:440];
  assign _02288_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21884" *) _04577_ : wt4_actv_data[439:432];
  assign _02287_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21874" *) _04576_ : wt4_actv_data[431:424];
  assign _02286_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21864" *) _04575_ : wt4_actv_data[423:416];
  assign _02285_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21854" *) _04574_ : wt4_actv_data[415:408];
  assign _02284_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21844" *) _04573_ : wt4_actv_data[407:400];
  assign _02282_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21834" *) _04572_ : wt4_actv_data[399:392];
  assign _02281_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21824" *) _04571_ : wt4_actv_data[391:384];
  assign _02280_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21814" *) _04570_ : wt4_actv_data[383:376];
  assign _02279_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21804" *) _04569_ : wt4_actv_data[375:368];
  assign _02278_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21794" *) _04568_ : wt4_actv_data[367:360];
  assign _02277_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21784" *) _04567_ : wt4_actv_data[359:352];
  assign _02276_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21774" *) _04566_ : wt4_actv_data[351:344];
  assign _02275_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21764" *) _04565_ : wt4_actv_data[343:336];
  assign _02274_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21754" *) _04564_ : wt4_actv_data[335:328];
  assign _02273_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21744" *) _04563_ : wt4_actv_data[327:320];
  assign _02271_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21734" *) _04562_ : wt4_actv_data[319:312];
  assign _02270_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21724" *) _04561_ : wt4_actv_data[311:304];
  assign _02269_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21714" *) _04560_ : wt4_actv_data[303:296];
  assign _02268_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21704" *) _04559_ : wt4_actv_data[295:288];
  assign _02267_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21694" *) _04558_ : wt4_actv_data[287:280];
  assign _02266_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21684" *) _04557_ : wt4_actv_data[279:272];
  assign _02265_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21674" *) _04556_ : wt4_actv_data[271:264];
  assign _02264_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21664" *) _04555_ : wt4_actv_data[263:256];
  assign _02263_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21654" *) _04554_ : wt4_actv_data[255:248];
  assign _02262_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21644" *) _04553_ : wt4_actv_data[247:240];
  assign _02260_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21634" *) _04552_ : wt4_actv_data[239:232];
  assign _02259_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21624" *) _04551_ : wt4_actv_data[231:224];
  assign _02258_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21614" *) _04550_ : wt4_actv_data[223:216];
  assign _02257_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21604" *) _04549_ : wt4_actv_data[215:208];
  assign _02256_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21594" *) _04548_ : wt4_actv_data[207:200];
  assign _02255_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21584" *) _04547_ : wt4_actv_data[199:192];
  assign _02254_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21574" *) _04546_ : wt4_actv_data[191:184];
  assign _02253_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21564" *) _04545_ : wt4_actv_data[183:176];
  assign _02252_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21554" *) _04544_ : wt4_actv_data[175:168];
  assign _02251_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21544" *) _04543_ : wt4_actv_data[167:160];
  assign _02249_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21534" *) _04542_ : wt4_actv_data[159:152];
  assign _02248_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21524" *) _04541_ : wt4_actv_data[151:144];
  assign _02247_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21514" *) _04540_ : wt4_actv_data[143:136];
  assign _02246_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21504" *) _04539_ : wt4_actv_data[135:128];
  assign _02245_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21494" *) _04538_ : wt4_actv_data[127:120];
  assign _02244_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21484" *) _04537_ : wt4_actv_data[119:112];
  assign _02243_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21474" *) _04536_ : wt4_actv_data[111:104];
  assign _02242_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21464" *) _04535_ : wt4_actv_data[103:96];
  assign _02361_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21454" *) _04534_ : wt4_actv_data[95:88];
  assign _02350_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21444" *) _04533_ : wt4_actv_data[87:80];
  assign _02338_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21434" *) _04532_ : wt4_actv_data[79:72];
  assign _02327_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21424" *) _04531_ : wt4_actv_data[71:64];
  assign _02316_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21414" *) _04530_ : wt4_actv_data[63:56];
  assign _02305_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21404" *) _04529_ : wt4_actv_data[55:48];
  assign _02294_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21394" *) _04528_ : wt4_actv_data[47:40];
  assign _02283_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21384" *) _04527_ : wt4_actv_data[39:32];
  assign _02272_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21374" *) _04526_ : wt4_actv_data[31:24];
  assign _02261_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21364" *) _04525_ : wt4_actv_data[23:16];
  assign _02250_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21354" *) _04524_ : wt4_actv_data[15:8];
  assign _02339_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21344" *) _04523_ : wt4_actv_data[7:0];
  assign _02367_ = _04522_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21334" *) wt4_sd_nan : wt4_actv_nan;
  assign _02368_ = _04521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21324" *) wt4_sd_nz : wt4_actv_nz;
  assign _01979_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21290" *) _04520_ : wt3_actv_data[1023:1016];
  assign _01978_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21280" *) _04519_ : wt3_actv_data[1015:1008];
  assign _01977_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21270" *) _04518_ : wt3_actv_data[1007:1000];
  assign _02104_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21260" *) _04517_ : wt3_actv_data[999:992];
  assign _02103_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21250" *) _04516_ : wt3_actv_data[991:984];
  assign _02102_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21240" *) _04515_ : wt3_actv_data[983:976];
  assign _02101_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21230" *) _04514_ : wt3_actv_data[975:968];
  assign _02100_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21220" *) _04513_ : wt3_actv_data[967:960];
  assign _02098_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21210" *) _04512_ : wt3_actv_data[959:952];
  assign _02097_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21200" *) _04511_ : wt3_actv_data[951:944];
  assign _02096_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21190" *) _04510_ : wt3_actv_data[943:936];
  assign _02095_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21180" *) _04509_ : wt3_actv_data[935:928];
  assign _02094_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21170" *) _04508_ : wt3_actv_data[927:920];
  assign _02093_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21160" *) _04507_ : wt3_actv_data[919:912];
  assign _02092_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21150" *) _04506_ : wt3_actv_data[911:904];
  assign _02091_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21140" *) _04505_ : wt3_actv_data[903:896];
  assign _02090_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21130" *) _04504_ : wt3_actv_data[895:888];
  assign _02089_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21120" *) _04503_ : wt3_actv_data[887:880];
  assign _02087_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21110" *) _04502_ : wt3_actv_data[879:872];
  assign _02086_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21100" *) _04501_ : wt3_actv_data[871:864];
  assign _02085_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21090" *) _04500_ : wt3_actv_data[863:856];
  assign _02084_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21080" *) _04499_ : wt3_actv_data[855:848];
  assign _02083_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21070" *) _04498_ : wt3_actv_data[847:840];
  assign _02082_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21060" *) _04497_ : wt3_actv_data[839:832];
  assign _02081_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21050" *) _04496_ : wt3_actv_data[831:824];
  assign _02080_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21040" *) _04495_ : wt3_actv_data[823:816];
  assign _02079_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21030" *) _04494_ : wt3_actv_data[815:808];
  assign _02078_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21020" *) _04493_ : wt3_actv_data[807:800];
  assign _02075_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21010" *) _04492_ : wt3_actv_data[799:792];
  assign _02074_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21000" *) _04491_ : wt3_actv_data[791:784];
  assign _02073_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20990" *) _04490_ : wt3_actv_data[783:776];
  assign _02072_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20980" *) _04489_ : wt3_actv_data[775:768];
  assign _02071_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20970" *) _04488_ : wt3_actv_data[767:760];
  assign _02070_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20960" *) _04487_ : wt3_actv_data[759:752];
  assign _02069_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20950" *) _04486_ : wt3_actv_data[751:744];
  assign _02068_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20940" *) _04485_ : wt3_actv_data[743:736];
  assign _02067_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20930" *) _04484_ : wt3_actv_data[735:728];
  assign _02066_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20920" *) _04483_ : wt3_actv_data[727:720];
  assign _02064_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20910" *) _04482_ : wt3_actv_data[719:712];
  assign _02063_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20900" *) _04481_ : wt3_actv_data[711:704];
  assign _02062_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20890" *) _04480_ : wt3_actv_data[703:696];
  assign _02061_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20880" *) _04479_ : wt3_actv_data[695:688];
  assign _02060_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20870" *) _04478_ : wt3_actv_data[687:680];
  assign _02059_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20860" *) _04477_ : wt3_actv_data[679:672];
  assign _02058_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20850" *) _04476_ : wt3_actv_data[671:664];
  assign _02057_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20840" *) _04475_ : wt3_actv_data[663:656];
  assign _02056_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20830" *) _04474_ : wt3_actv_data[655:648];
  assign _02055_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20820" *) _04473_ : wt3_actv_data[647:640];
  assign _02053_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20810" *) _04472_ : wt3_actv_data[639:632];
  assign _02052_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20800" *) _04471_ : wt3_actv_data[631:624];
  assign _02051_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20790" *) _04470_ : wt3_actv_data[623:616];
  assign _02050_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20780" *) _04469_ : wt3_actv_data[615:608];
  assign _02049_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20770" *) _04468_ : wt3_actv_data[607:600];
  assign _02048_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20760" *) _04467_ : wt3_actv_data[599:592];
  assign _02047_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20750" *) _04466_ : wt3_actv_data[591:584];
  assign _02046_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20740" *) _04465_ : wt3_actv_data[583:576];
  assign _02045_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20730" *) _04464_ : wt3_actv_data[575:568];
  assign _02044_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20720" *) _04463_ : wt3_actv_data[567:560];
  assign _02042_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20710" *) _04462_ : wt3_actv_data[559:552];
  assign _02041_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20700" *) _04461_ : wt3_actv_data[551:544];
  assign _02040_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20690" *) _04460_ : wt3_actv_data[543:536];
  assign _02039_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20680" *) _04459_ : wt3_actv_data[535:528];
  assign _02038_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20670" *) _04458_ : wt3_actv_data[527:520];
  assign _02037_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20660" *) _04457_ : wt3_actv_data[519:512];
  assign _02036_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20650" *) _04456_ : wt3_actv_data[511:504];
  assign _02035_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20640" *) _04455_ : wt3_actv_data[503:496];
  assign _02034_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20630" *) _04454_ : wt3_actv_data[495:488];
  assign _02033_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20620" *) _04453_ : wt3_actv_data[487:480];
  assign _02031_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20610" *) _04452_ : wt3_actv_data[479:472];
  assign _02030_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20600" *) _04451_ : wt3_actv_data[471:464];
  assign _02029_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20590" *) _04450_ : wt3_actv_data[463:456];
  assign _02028_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20580" *) _04449_ : wt3_actv_data[455:448];
  assign _02027_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20570" *) _04448_ : wt3_actv_data[447:440];
  assign _02026_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20560" *) _04447_ : wt3_actv_data[439:432];
  assign _02025_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20550" *) _04446_ : wt3_actv_data[431:424];
  assign _02024_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20540" *) _04445_ : wt3_actv_data[423:416];
  assign _02023_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20530" *) _04444_ : wt3_actv_data[415:408];
  assign _02022_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20520" *) _04443_ : wt3_actv_data[407:400];
  assign _02020_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20510" *) _04442_ : wt3_actv_data[399:392];
  assign _02019_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20500" *) _04441_ : wt3_actv_data[391:384];
  assign _02018_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20490" *) _04440_ : wt3_actv_data[383:376];
  assign _02017_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20480" *) _04439_ : wt3_actv_data[375:368];
  assign _02016_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20470" *) _04438_ : wt3_actv_data[367:360];
  assign _02015_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20460" *) _04437_ : wt3_actv_data[359:352];
  assign _02014_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20450" *) _04436_ : wt3_actv_data[351:344];
  assign _02013_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20440" *) _04435_ : wt3_actv_data[343:336];
  assign _02012_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20430" *) _04434_ : wt3_actv_data[335:328];
  assign _02011_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20420" *) _04433_ : wt3_actv_data[327:320];
  assign _02009_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20410" *) _04432_ : wt3_actv_data[319:312];
  assign _02008_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20400" *) _04431_ : wt3_actv_data[311:304];
  assign _02007_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20390" *) _04430_ : wt3_actv_data[303:296];
  assign _02006_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20380" *) _04429_ : wt3_actv_data[295:288];
  assign _02005_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20370" *) _04428_ : wt3_actv_data[287:280];
  assign _02004_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20360" *) _04427_ : wt3_actv_data[279:272];
  assign _02003_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20350" *) _04426_ : wt3_actv_data[271:264];
  assign _02002_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20340" *) _04425_ : wt3_actv_data[263:256];
  assign _02001_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20330" *) _04424_ : wt3_actv_data[255:248];
  assign _02000_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20320" *) _04423_ : wt3_actv_data[247:240];
  assign _01998_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20310" *) _04422_ : wt3_actv_data[239:232];
  assign _01997_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20300" *) _04421_ : wt3_actv_data[231:224];
  assign _01996_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20290" *) _04420_ : wt3_actv_data[223:216];
  assign _01995_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20280" *) _04419_ : wt3_actv_data[215:208];
  assign _01994_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20270" *) _04418_ : wt3_actv_data[207:200];
  assign _01993_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20260" *) _04417_ : wt3_actv_data[199:192];
  assign _01992_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20250" *) _04416_ : wt3_actv_data[191:184];
  assign _01991_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20240" *) _04415_ : wt3_actv_data[183:176];
  assign _01990_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20230" *) _04414_ : wt3_actv_data[175:168];
  assign _01989_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20220" *) _04413_ : wt3_actv_data[167:160];
  assign _01987_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20210" *) _04412_ : wt3_actv_data[159:152];
  assign _01986_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20200" *) _04411_ : wt3_actv_data[151:144];
  assign _01985_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20190" *) _04410_ : wt3_actv_data[143:136];
  assign _01984_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20180" *) _04409_ : wt3_actv_data[135:128];
  assign _01983_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20170" *) _04408_ : wt3_actv_data[127:120];
  assign _01982_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20160" *) _04407_ : wt3_actv_data[119:112];
  assign _01981_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20150" *) _04406_ : wt3_actv_data[111:104];
  assign _01980_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20140" *) _04405_ : wt3_actv_data[103:96];
  assign _02099_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20130" *) _04404_ : wt3_actv_data[95:88];
  assign _02088_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20120" *) _04403_ : wt3_actv_data[87:80];
  assign _02076_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20110" *) _04402_ : wt3_actv_data[79:72];
  assign _02065_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20100" *) _04401_ : wt3_actv_data[71:64];
  assign _02054_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20090" *) _04400_ : wt3_actv_data[63:56];
  assign _02043_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20080" *) _04399_ : wt3_actv_data[55:48];
  assign _02032_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20070" *) _04398_ : wt3_actv_data[47:40];
  assign _02021_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20060" *) _04397_ : wt3_actv_data[39:32];
  assign _02010_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20050" *) _04396_ : wt3_actv_data[31:24];
  assign _01999_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20040" *) _04395_ : wt3_actv_data[23:16];
  assign _01988_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20030" *) _04394_ : wt3_actv_data[15:8];
  assign _02077_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20020" *) _04393_ : wt3_actv_data[7:0];
  assign _02105_ = _04392_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20010" *) wt3_sd_nan : wt3_actv_nan;
  assign _02106_ = _04391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:20000" *) wt3_sd_nz : wt3_actv_nz;
  assign _01717_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19966" *) _04390_ : wt2_actv_data[1023:1016];
  assign _01716_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19956" *) _04389_ : wt2_actv_data[1015:1008];
  assign _01715_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19946" *) _04388_ : wt2_actv_data[1007:1000];
  assign _01842_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19936" *) _04387_ : wt2_actv_data[999:992];
  assign _01841_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19926" *) _04386_ : wt2_actv_data[991:984];
  assign _01840_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19916" *) _04385_ : wt2_actv_data[983:976];
  assign _01839_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19906" *) _04384_ : wt2_actv_data[975:968];
  assign _01838_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19896" *) _04383_ : wt2_actv_data[967:960];
  assign _01836_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19886" *) _04382_ : wt2_actv_data[959:952];
  assign _01835_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19876" *) _04381_ : wt2_actv_data[951:944];
  assign _01834_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19866" *) _04380_ : wt2_actv_data[943:936];
  assign _01833_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19856" *) _04379_ : wt2_actv_data[935:928];
  assign _01832_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19846" *) _04378_ : wt2_actv_data[927:920];
  assign _01831_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19836" *) _04377_ : wt2_actv_data[919:912];
  assign _01830_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19826" *) _04376_ : wt2_actv_data[911:904];
  assign _01829_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19816" *) _04375_ : wt2_actv_data[903:896];
  assign _01828_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19806" *) _04374_ : wt2_actv_data[895:888];
  assign _01827_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19796" *) _04373_ : wt2_actv_data[887:880];
  assign _01825_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19786" *) _04372_ : wt2_actv_data[879:872];
  assign _01824_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19776" *) _04371_ : wt2_actv_data[871:864];
  assign _01823_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19766" *) _04370_ : wt2_actv_data[863:856];
  assign _01822_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19756" *) _04369_ : wt2_actv_data[855:848];
  assign _01821_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19746" *) _04368_ : wt2_actv_data[847:840];
  assign _01820_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19736" *) _04367_ : wt2_actv_data[839:832];
  assign _01819_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19726" *) _04366_ : wt2_actv_data[831:824];
  assign _01818_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19716" *) _04365_ : wt2_actv_data[823:816];
  assign _01817_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19706" *) _04364_ : wt2_actv_data[815:808];
  assign _01816_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19696" *) _04363_ : wt2_actv_data[807:800];
  assign _01813_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19686" *) _04362_ : wt2_actv_data[799:792];
  assign _01812_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19676" *) _04361_ : wt2_actv_data[791:784];
  assign _01811_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19666" *) _04360_ : wt2_actv_data[783:776];
  assign _01810_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19656" *) _04359_ : wt2_actv_data[775:768];
  assign _01809_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19646" *) _04358_ : wt2_actv_data[767:760];
  assign _01808_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19636" *) _04357_ : wt2_actv_data[759:752];
  assign _01807_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19626" *) _04356_ : wt2_actv_data[751:744];
  assign _01806_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19616" *) _04355_ : wt2_actv_data[743:736];
  assign _01805_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19606" *) _04354_ : wt2_actv_data[735:728];
  assign _01804_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19596" *) _04353_ : wt2_actv_data[727:720];
  assign _01802_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19586" *) _04352_ : wt2_actv_data[719:712];
  assign _01801_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19576" *) _04351_ : wt2_actv_data[711:704];
  assign _01800_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19566" *) _04350_ : wt2_actv_data[703:696];
  assign _01799_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19556" *) _04349_ : wt2_actv_data[695:688];
  assign _01798_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19546" *) _04348_ : wt2_actv_data[687:680];
  assign _01797_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19536" *) _04347_ : wt2_actv_data[679:672];
  assign _01796_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19526" *) _04346_ : wt2_actv_data[671:664];
  assign _01795_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19516" *) _04345_ : wt2_actv_data[663:656];
  assign _01794_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19506" *) _04344_ : wt2_actv_data[655:648];
  assign _01793_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19496" *) _04343_ : wt2_actv_data[647:640];
  assign _01791_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19486" *) _04342_ : wt2_actv_data[639:632];
  assign _01790_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19476" *) _04341_ : wt2_actv_data[631:624];
  assign _01789_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19466" *) _04340_ : wt2_actv_data[623:616];
  assign _01788_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19456" *) _04339_ : wt2_actv_data[615:608];
  assign _01787_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19446" *) _04338_ : wt2_actv_data[607:600];
  assign _01786_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19436" *) _04337_ : wt2_actv_data[599:592];
  assign _01785_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19426" *) _04336_ : wt2_actv_data[591:584];
  assign _01784_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19416" *) _04335_ : wt2_actv_data[583:576];
  assign _01783_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19406" *) _04334_ : wt2_actv_data[575:568];
  assign _01782_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19396" *) _04333_ : wt2_actv_data[567:560];
  assign _01780_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19386" *) _04332_ : wt2_actv_data[559:552];
  assign _01779_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19376" *) _04331_ : wt2_actv_data[551:544];
  assign _01778_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19366" *) _04330_ : wt2_actv_data[543:536];
  assign _01777_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19356" *) _04329_ : wt2_actv_data[535:528];
  assign _01776_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19346" *) _04328_ : wt2_actv_data[527:520];
  assign _01775_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19336" *) _04327_ : wt2_actv_data[519:512];
  assign _01774_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19326" *) _04326_ : wt2_actv_data[511:504];
  assign _01773_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19316" *) _04325_ : wt2_actv_data[503:496];
  assign _01772_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19306" *) _04324_ : wt2_actv_data[495:488];
  assign _01771_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19296" *) _04323_ : wt2_actv_data[487:480];
  assign _01769_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19286" *) _04322_ : wt2_actv_data[479:472];
  assign _01768_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19276" *) _04321_ : wt2_actv_data[471:464];
  assign _01767_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19266" *) _04320_ : wt2_actv_data[463:456];
  assign _01766_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19256" *) _04319_ : wt2_actv_data[455:448];
  assign _01765_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19246" *) _04318_ : wt2_actv_data[447:440];
  assign _01764_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19236" *) _04317_ : wt2_actv_data[439:432];
  assign _01763_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19226" *) _04316_ : wt2_actv_data[431:424];
  assign _01762_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19216" *) _04315_ : wt2_actv_data[423:416];
  assign _01761_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19206" *) _04314_ : wt2_actv_data[415:408];
  assign _01760_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19196" *) _04313_ : wt2_actv_data[407:400];
  assign _01758_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19186" *) _04312_ : wt2_actv_data[399:392];
  assign _01757_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19176" *) _04311_ : wt2_actv_data[391:384];
  assign _01756_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19166" *) _04310_ : wt2_actv_data[383:376];
  assign _01755_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19156" *) _04309_ : wt2_actv_data[375:368];
  assign _01754_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19146" *) _04308_ : wt2_actv_data[367:360];
  assign _01753_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19136" *) _04307_ : wt2_actv_data[359:352];
  assign _01752_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19126" *) _04306_ : wt2_actv_data[351:344];
  assign _01751_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19116" *) _04305_ : wt2_actv_data[343:336];
  assign _01750_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19106" *) _04304_ : wt2_actv_data[335:328];
  assign _01749_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19096" *) _04303_ : wt2_actv_data[327:320];
  assign _01747_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19086" *) _04302_ : wt2_actv_data[319:312];
  assign _01746_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19076" *) _04301_ : wt2_actv_data[311:304];
  assign _01745_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19066" *) _04300_ : wt2_actv_data[303:296];
  assign _01744_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19056" *) _04299_ : wt2_actv_data[295:288];
  assign _01743_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19046" *) _04298_ : wt2_actv_data[287:280];
  assign _01742_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19036" *) _04297_ : wt2_actv_data[279:272];
  assign _01741_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19026" *) _04296_ : wt2_actv_data[271:264];
  assign _01740_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19016" *) _04295_ : wt2_actv_data[263:256];
  assign _01739_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19006" *) _04294_ : wt2_actv_data[255:248];
  assign _01738_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18996" *) _04293_ : wt2_actv_data[247:240];
  assign _01736_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18986" *) _04292_ : wt2_actv_data[239:232];
  assign _01735_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18976" *) _04291_ : wt2_actv_data[231:224];
  assign _01734_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18966" *) _04290_ : wt2_actv_data[223:216];
  assign _01733_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18956" *) _04289_ : wt2_actv_data[215:208];
  assign _01732_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18946" *) _04288_ : wt2_actv_data[207:200];
  assign _01731_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18936" *) _04287_ : wt2_actv_data[199:192];
  assign _01730_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18926" *) _04286_ : wt2_actv_data[191:184];
  assign _01729_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18916" *) _04285_ : wt2_actv_data[183:176];
  assign _01728_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18906" *) _04284_ : wt2_actv_data[175:168];
  assign _01727_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18896" *) _04283_ : wt2_actv_data[167:160];
  assign _01725_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18886" *) _04282_ : wt2_actv_data[159:152];
  assign _01724_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18876" *) _04281_ : wt2_actv_data[151:144];
  assign _01723_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18866" *) _04280_ : wt2_actv_data[143:136];
  assign _01722_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18856" *) _04279_ : wt2_actv_data[135:128];
  assign _01721_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18846" *) _04278_ : wt2_actv_data[127:120];
  assign _01720_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18836" *) _04277_ : wt2_actv_data[119:112];
  assign _01719_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18826" *) _04276_ : wt2_actv_data[111:104];
  assign _01718_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18816" *) _04275_ : wt2_actv_data[103:96];
  assign _01837_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18806" *) _04274_ : wt2_actv_data[95:88];
  assign _01826_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18796" *) _04273_ : wt2_actv_data[87:80];
  assign _01814_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18786" *) _04272_ : wt2_actv_data[79:72];
  assign _01803_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18776" *) _04271_ : wt2_actv_data[71:64];
  assign _01792_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18766" *) _04270_ : wt2_actv_data[63:56];
  assign _01781_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18756" *) _04269_ : wt2_actv_data[55:48];
  assign _01770_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18746" *) _04268_ : wt2_actv_data[47:40];
  assign _01759_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18736" *) _04267_ : wt2_actv_data[39:32];
  assign _01748_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18726" *) _04266_ : wt2_actv_data[31:24];
  assign _01737_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18716" *) _04265_ : wt2_actv_data[23:16];
  assign _01726_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18706" *) _04264_ : wt2_actv_data[15:8];
  assign _01815_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18696" *) _04263_ : wt2_actv_data[7:0];
  assign _01843_ = _04262_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18686" *) wt2_sd_nan : wt2_actv_nan;
  assign _01844_ = _04261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18676" *) wt2_sd_nz : wt2_actv_nz;
  assign _01455_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18642" *) _04260_ : wt1_actv_data[1023:1016];
  assign _01454_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18632" *) _04259_ : wt1_actv_data[1015:1008];
  assign _01453_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18622" *) _04258_ : wt1_actv_data[1007:1000];
  assign _01580_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18612" *) _04257_ : wt1_actv_data[999:992];
  assign _01579_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18602" *) _04256_ : wt1_actv_data[991:984];
  assign _01578_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18592" *) _04255_ : wt1_actv_data[983:976];
  assign _01577_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18582" *) _04254_ : wt1_actv_data[975:968];
  assign _01576_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18572" *) _04253_ : wt1_actv_data[967:960];
  assign _01574_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18562" *) _04252_ : wt1_actv_data[959:952];
  assign _01573_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18552" *) _04251_ : wt1_actv_data[951:944];
  assign _01572_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18542" *) _04250_ : wt1_actv_data[943:936];
  assign _01571_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18532" *) _04249_ : wt1_actv_data[935:928];
  assign _01570_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18522" *) _04248_ : wt1_actv_data[927:920];
  assign _01569_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18512" *) _04247_ : wt1_actv_data[919:912];
  assign _01568_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18502" *) _04246_ : wt1_actv_data[911:904];
  assign _01567_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18492" *) _04245_ : wt1_actv_data[903:896];
  assign _01566_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18482" *) _04244_ : wt1_actv_data[895:888];
  assign _01565_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18472" *) _04243_ : wt1_actv_data[887:880];
  assign _01563_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18462" *) _04242_ : wt1_actv_data[879:872];
  assign _01562_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18452" *) _04241_ : wt1_actv_data[871:864];
  assign _01561_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18442" *) _04240_ : wt1_actv_data[863:856];
  assign _01560_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18432" *) _04239_ : wt1_actv_data[855:848];
  assign _01559_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18422" *) _04238_ : wt1_actv_data[847:840];
  assign _01558_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18412" *) _04237_ : wt1_actv_data[839:832];
  assign _01557_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18402" *) _04236_ : wt1_actv_data[831:824];
  assign _01556_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18392" *) _04235_ : wt1_actv_data[823:816];
  assign _01555_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18382" *) _04234_ : wt1_actv_data[815:808];
  assign _01554_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18372" *) _04233_ : wt1_actv_data[807:800];
  assign _01551_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18362" *) _04232_ : wt1_actv_data[799:792];
  assign _01550_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18352" *) _04231_ : wt1_actv_data[791:784];
  assign _01549_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18342" *) _04230_ : wt1_actv_data[783:776];
  assign _01548_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18332" *) _04229_ : wt1_actv_data[775:768];
  assign _01547_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18322" *) _04228_ : wt1_actv_data[767:760];
  assign _01546_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18312" *) _04227_ : wt1_actv_data[759:752];
  assign _01545_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18302" *) _04226_ : wt1_actv_data[751:744];
  assign _01544_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18292" *) _04225_ : wt1_actv_data[743:736];
  assign _01543_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18282" *) _04224_ : wt1_actv_data[735:728];
  assign _01542_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18272" *) _04223_ : wt1_actv_data[727:720];
  assign _01540_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18262" *) _04222_ : wt1_actv_data[719:712];
  assign _01539_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18252" *) _04221_ : wt1_actv_data[711:704];
  assign _01538_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18242" *) _04220_ : wt1_actv_data[703:696];
  assign _01537_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18232" *) _04219_ : wt1_actv_data[695:688];
  assign _01536_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18222" *) _04218_ : wt1_actv_data[687:680];
  assign _01535_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18212" *) _04217_ : wt1_actv_data[679:672];
  assign _01534_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18202" *) _04216_ : wt1_actv_data[671:664];
  assign _01533_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18192" *) _04215_ : wt1_actv_data[663:656];
  assign _01532_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18182" *) _04214_ : wt1_actv_data[655:648];
  assign _01531_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18172" *) _04213_ : wt1_actv_data[647:640];
  assign _01529_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18162" *) _04212_ : wt1_actv_data[639:632];
  assign _01528_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18152" *) _04211_ : wt1_actv_data[631:624];
  assign _01527_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18142" *) _04210_ : wt1_actv_data[623:616];
  assign _01526_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18132" *) _04209_ : wt1_actv_data[615:608];
  assign _01525_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18122" *) _04208_ : wt1_actv_data[607:600];
  assign _01524_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18112" *) _04207_ : wt1_actv_data[599:592];
  assign _01523_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18102" *) _04206_ : wt1_actv_data[591:584];
  assign _01522_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18092" *) _04205_ : wt1_actv_data[583:576];
  assign _01521_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18082" *) _04204_ : wt1_actv_data[575:568];
  assign _01520_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18072" *) _04203_ : wt1_actv_data[567:560];
  assign _01518_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18062" *) _04202_ : wt1_actv_data[559:552];
  assign _01517_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18052" *) _04201_ : wt1_actv_data[551:544];
  assign _01516_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18042" *) _04200_ : wt1_actv_data[543:536];
  assign _01515_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18032" *) _04199_ : wt1_actv_data[535:528];
  assign _01514_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18022" *) _04198_ : wt1_actv_data[527:520];
  assign _01513_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18012" *) _04197_ : wt1_actv_data[519:512];
  assign _01512_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18002" *) _04196_ : wt1_actv_data[511:504];
  assign _01511_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17992" *) _04195_ : wt1_actv_data[503:496];
  assign _01510_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17982" *) _04194_ : wt1_actv_data[495:488];
  assign _01509_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17972" *) _04193_ : wt1_actv_data[487:480];
  assign _01507_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17962" *) _04192_ : wt1_actv_data[479:472];
  assign _01506_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17952" *) _04191_ : wt1_actv_data[471:464];
  assign _01505_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17942" *) _04190_ : wt1_actv_data[463:456];
  assign _01504_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17932" *) _04189_ : wt1_actv_data[455:448];
  assign _01503_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17922" *) _04188_ : wt1_actv_data[447:440];
  assign _01502_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17912" *) _04187_ : wt1_actv_data[439:432];
  assign _01501_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17902" *) _04186_ : wt1_actv_data[431:424];
  assign _01500_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17892" *) _04185_ : wt1_actv_data[423:416];
  assign _01499_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17882" *) _04184_ : wt1_actv_data[415:408];
  assign _01498_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17872" *) _04183_ : wt1_actv_data[407:400];
  assign _01496_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17862" *) _04182_ : wt1_actv_data[399:392];
  assign _01495_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17852" *) _04181_ : wt1_actv_data[391:384];
  assign _01494_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17842" *) _04180_ : wt1_actv_data[383:376];
  assign _01493_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17832" *) _04179_ : wt1_actv_data[375:368];
  assign _01492_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17822" *) _04178_ : wt1_actv_data[367:360];
  assign _01491_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17812" *) _04177_ : wt1_actv_data[359:352];
  assign _01490_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17802" *) _04176_ : wt1_actv_data[351:344];
  assign _01489_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17792" *) _04175_ : wt1_actv_data[343:336];
  assign _01488_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17782" *) _04174_ : wt1_actv_data[335:328];
  assign _01487_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17772" *) _04173_ : wt1_actv_data[327:320];
  assign _01485_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17762" *) _04172_ : wt1_actv_data[319:312];
  assign _01484_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17752" *) _04171_ : wt1_actv_data[311:304];
  assign _01483_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17742" *) _04170_ : wt1_actv_data[303:296];
  assign _01482_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17732" *) _04169_ : wt1_actv_data[295:288];
  assign _01481_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17722" *) _04168_ : wt1_actv_data[287:280];
  assign _01480_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17712" *) _04167_ : wt1_actv_data[279:272];
  assign _01479_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17702" *) _04166_ : wt1_actv_data[271:264];
  assign _01478_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17692" *) _04165_ : wt1_actv_data[263:256];
  assign _01477_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17682" *) _04164_ : wt1_actv_data[255:248];
  assign _01476_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17672" *) _04163_ : wt1_actv_data[247:240];
  assign _01474_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17662" *) _04162_ : wt1_actv_data[239:232];
  assign _01473_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17652" *) _04161_ : wt1_actv_data[231:224];
  assign _01472_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17642" *) _04160_ : wt1_actv_data[223:216];
  assign _01471_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17632" *) _04159_ : wt1_actv_data[215:208];
  assign _01470_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17622" *) _04158_ : wt1_actv_data[207:200];
  assign _01469_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17612" *) _04157_ : wt1_actv_data[199:192];
  assign _01468_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17602" *) _04156_ : wt1_actv_data[191:184];
  assign _01467_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17592" *) _04155_ : wt1_actv_data[183:176];
  assign _01466_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17582" *) _04154_ : wt1_actv_data[175:168];
  assign _01465_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17572" *) _04153_ : wt1_actv_data[167:160];
  assign _01463_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17562" *) _04152_ : wt1_actv_data[159:152];
  assign _01462_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17552" *) _04151_ : wt1_actv_data[151:144];
  assign _01461_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17542" *) _04150_ : wt1_actv_data[143:136];
  assign _01460_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17532" *) _04149_ : wt1_actv_data[135:128];
  assign _01459_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17522" *) _04148_ : wt1_actv_data[127:120];
  assign _01458_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17512" *) _04147_ : wt1_actv_data[119:112];
  assign _01457_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17502" *) _04146_ : wt1_actv_data[111:104];
  assign _01456_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17492" *) _04145_ : wt1_actv_data[103:96];
  assign _01575_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17482" *) _04144_ : wt1_actv_data[95:88];
  assign _01564_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17472" *) _04143_ : wt1_actv_data[87:80];
  assign _01552_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17462" *) _04142_ : wt1_actv_data[79:72];
  assign _01541_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17452" *) _04141_ : wt1_actv_data[71:64];
  assign _01530_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17442" *) _04140_ : wt1_actv_data[63:56];
  assign _01519_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17432" *) _04139_ : wt1_actv_data[55:48];
  assign _01508_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17422" *) _04138_ : wt1_actv_data[47:40];
  assign _01497_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17412" *) _04137_ : wt1_actv_data[39:32];
  assign _01486_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17402" *) _04136_ : wt1_actv_data[31:24];
  assign _01475_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17392" *) _04135_ : wt1_actv_data[23:16];
  assign _01464_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17382" *) _04134_ : wt1_actv_data[15:8];
  assign _01553_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17372" *) _04133_ : wt1_actv_data[7:0];
  assign _01581_ = _04132_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17362" *) wt1_sd_nan : wt1_actv_nan;
  assign _01582_ = _04131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17352" *) wt1_sd_nz : wt1_actv_nz;
  assign _01193_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17318" *) _04130_ : wt0_actv_data[1023:1016];
  assign _01192_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17308" *) _04129_ : wt0_actv_data[1015:1008];
  assign _01191_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17298" *) _04128_ : wt0_actv_data[1007:1000];
  assign _01318_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17288" *) _04127_ : wt0_actv_data[999:992];
  assign _01317_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17278" *) _04126_ : wt0_actv_data[991:984];
  assign _01316_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17268" *) _04125_ : wt0_actv_data[983:976];
  assign _01315_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17258" *) _04124_ : wt0_actv_data[975:968];
  assign _01314_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17248" *) _04123_ : wt0_actv_data[967:960];
  assign _01312_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17238" *) _04122_ : wt0_actv_data[959:952];
  assign _01311_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17228" *) _04121_ : wt0_actv_data[951:944];
  assign _01310_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17218" *) _04120_ : wt0_actv_data[943:936];
  assign _01309_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17208" *) _04119_ : wt0_actv_data[935:928];
  assign _01308_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17198" *) _04118_ : wt0_actv_data[927:920];
  assign _01307_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17188" *) _04117_ : wt0_actv_data[919:912];
  assign _01306_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17178" *) _04116_ : wt0_actv_data[911:904];
  assign _01305_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17168" *) _04115_ : wt0_actv_data[903:896];
  assign _01304_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17158" *) _04114_ : wt0_actv_data[895:888];
  assign _01303_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17148" *) _04113_ : wt0_actv_data[887:880];
  assign _01301_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17138" *) _04112_ : wt0_actv_data[879:872];
  assign _01300_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17128" *) _04111_ : wt0_actv_data[871:864];
  assign _01299_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17118" *) _04110_ : wt0_actv_data[863:856];
  assign _01298_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17108" *) _04109_ : wt0_actv_data[855:848];
  assign _01297_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17098" *) _04108_ : wt0_actv_data[847:840];
  assign _01296_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17088" *) _04107_ : wt0_actv_data[839:832];
  assign _01295_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17078" *) _04106_ : wt0_actv_data[831:824];
  assign _01294_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17068" *) _04105_ : wt0_actv_data[823:816];
  assign _01293_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17058" *) _04104_ : wt0_actv_data[815:808];
  assign _01292_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17048" *) _04103_ : wt0_actv_data[807:800];
  assign _01289_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17038" *) _04102_ : wt0_actv_data[799:792];
  assign _01288_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17028" *) _04101_ : wt0_actv_data[791:784];
  assign _01287_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17018" *) _04100_ : wt0_actv_data[783:776];
  assign _01286_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17008" *) _04099_ : wt0_actv_data[775:768];
  assign _01285_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16998" *) _04098_ : wt0_actv_data[767:760];
  assign _01284_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16988" *) _04097_ : wt0_actv_data[759:752];
  assign _01283_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16978" *) _04096_ : wt0_actv_data[751:744];
  assign _01282_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16968" *) _04095_ : wt0_actv_data[743:736];
  assign _01281_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16958" *) _04094_ : wt0_actv_data[735:728];
  assign _01280_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16948" *) _04093_ : wt0_actv_data[727:720];
  assign _01278_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16938" *) _04092_ : wt0_actv_data[719:712];
  assign _01277_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16928" *) _04091_ : wt0_actv_data[711:704];
  assign _01276_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16918" *) _04090_ : wt0_actv_data[703:696];
  assign _01275_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16908" *) _04089_ : wt0_actv_data[695:688];
  assign _01274_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16898" *) _04088_ : wt0_actv_data[687:680];
  assign _01273_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16888" *) _04087_ : wt0_actv_data[679:672];
  assign _01272_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16878" *) _04086_ : wt0_actv_data[671:664];
  assign _01271_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16868" *) _04085_ : wt0_actv_data[663:656];
  assign _01270_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16858" *) _04084_ : wt0_actv_data[655:648];
  assign _01269_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16848" *) _04083_ : wt0_actv_data[647:640];
  assign _01267_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16838" *) _04082_ : wt0_actv_data[639:632];
  assign _01266_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16828" *) _04081_ : wt0_actv_data[631:624];
  assign _01265_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16818" *) _04080_ : wt0_actv_data[623:616];
  assign _01264_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16808" *) _04079_ : wt0_actv_data[615:608];
  assign _01263_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16798" *) _04078_ : wt0_actv_data[607:600];
  assign _01262_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16788" *) _04077_ : wt0_actv_data[599:592];
  assign _01261_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16778" *) _04076_ : wt0_actv_data[591:584];
  assign _01260_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16768" *) _04075_ : wt0_actv_data[583:576];
  assign _01259_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16758" *) _04074_ : wt0_actv_data[575:568];
  assign _01258_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16748" *) _04073_ : wt0_actv_data[567:560];
  assign _01256_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16738" *) _04072_ : wt0_actv_data[559:552];
  assign _01255_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16728" *) _04071_ : wt0_actv_data[551:544];
  assign _01254_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16718" *) _04070_ : wt0_actv_data[543:536];
  assign _01253_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16708" *) _04069_ : wt0_actv_data[535:528];
  assign _01252_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16698" *) _04068_ : wt0_actv_data[527:520];
  assign _01251_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16688" *) _04067_ : wt0_actv_data[519:512];
  assign _01250_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16678" *) _04066_ : wt0_actv_data[511:504];
  assign _01249_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16668" *) _04065_ : wt0_actv_data[503:496];
  assign _01248_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16658" *) _04064_ : wt0_actv_data[495:488];
  assign _01247_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16648" *) _04063_ : wt0_actv_data[487:480];
  assign _01245_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16638" *) _04062_ : wt0_actv_data[479:472];
  assign _01244_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16628" *) _04061_ : wt0_actv_data[471:464];
  assign _01243_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16618" *) _04060_ : wt0_actv_data[463:456];
  assign _01242_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16608" *) _04059_ : wt0_actv_data[455:448];
  assign _01241_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16598" *) _04058_ : wt0_actv_data[447:440];
  assign _01240_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16588" *) _04057_ : wt0_actv_data[439:432];
  assign _01239_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16578" *) _04056_ : wt0_actv_data[431:424];
  assign _01238_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16568" *) _04055_ : wt0_actv_data[423:416];
  assign _01237_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16558" *) _04054_ : wt0_actv_data[415:408];
  assign _01236_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16548" *) _04053_ : wt0_actv_data[407:400];
  assign _01234_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16538" *) _04052_ : wt0_actv_data[399:392];
  assign _01233_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16528" *) _04051_ : wt0_actv_data[391:384];
  assign _01232_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16518" *) _04050_ : wt0_actv_data[383:376];
  assign _01231_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16508" *) _04049_ : wt0_actv_data[375:368];
  assign _01230_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16498" *) _04048_ : wt0_actv_data[367:360];
  assign _01229_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16488" *) _04047_ : wt0_actv_data[359:352];
  assign _01228_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16478" *) _04046_ : wt0_actv_data[351:344];
  assign _01227_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16468" *) _04045_ : wt0_actv_data[343:336];
  assign _01226_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16458" *) _04044_ : wt0_actv_data[335:328];
  assign _01225_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16448" *) _04043_ : wt0_actv_data[327:320];
  assign _01223_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16438" *) _04042_ : wt0_actv_data[319:312];
  assign _01222_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16428" *) _04041_ : wt0_actv_data[311:304];
  assign _01221_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16418" *) _04040_ : wt0_actv_data[303:296];
  assign _01220_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16408" *) _04039_ : wt0_actv_data[295:288];
  assign _01219_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16398" *) _04038_ : wt0_actv_data[287:280];
  assign _01218_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16388" *) _04037_ : wt0_actv_data[279:272];
  assign _01217_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16378" *) _04036_ : wt0_actv_data[271:264];
  assign _01216_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16368" *) _04035_ : wt0_actv_data[263:256];
  assign _01215_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16358" *) _04034_ : wt0_actv_data[255:248];
  assign _01214_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16348" *) _04033_ : wt0_actv_data[247:240];
  assign _01212_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16338" *) _04032_ : wt0_actv_data[239:232];
  assign _01211_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16328" *) _04031_ : wt0_actv_data[231:224];
  assign _01210_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16318" *) _04030_ : wt0_actv_data[223:216];
  assign _01209_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16308" *) _04029_ : wt0_actv_data[215:208];
  assign _01208_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16298" *) _04028_ : wt0_actv_data[207:200];
  assign _01207_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16288" *) _04027_ : wt0_actv_data[199:192];
  assign _01206_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16278" *) _04026_ : wt0_actv_data[191:184];
  assign _01205_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16268" *) _04025_ : wt0_actv_data[183:176];
  assign _01204_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16258" *) _04024_ : wt0_actv_data[175:168];
  assign _01203_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16248" *) _04023_ : wt0_actv_data[167:160];
  assign _01201_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16238" *) _04022_ : wt0_actv_data[159:152];
  assign _01200_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16228" *) _04021_ : wt0_actv_data[151:144];
  assign _01199_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16218" *) _04020_ : wt0_actv_data[143:136];
  assign _01198_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16208" *) _04019_ : wt0_actv_data[135:128];
  assign _01197_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16198" *) _04018_ : wt0_actv_data[127:120];
  assign _01196_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16188" *) _04017_ : wt0_actv_data[119:112];
  assign _01195_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16178" *) _04016_ : wt0_actv_data[111:104];
  assign _01194_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16168" *) _04015_ : wt0_actv_data[103:96];
  assign _01313_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16158" *) _04014_ : wt0_actv_data[95:88];
  assign _01302_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16148" *) _04013_ : wt0_actv_data[87:80];
  assign _01290_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16138" *) _04012_ : wt0_actv_data[79:72];
  assign _01279_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16128" *) _04011_ : wt0_actv_data[71:64];
  assign _01268_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16118" *) _04010_ : wt0_actv_data[63:56];
  assign _01257_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16108" *) _04009_ : wt0_actv_data[55:48];
  assign _01246_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16098" *) _04008_ : wt0_actv_data[47:40];
  assign _01235_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16088" *) _04007_ : wt0_actv_data[39:32];
  assign _01224_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16078" *) _04006_ : wt0_actv_data[31:24];
  assign _01213_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16068" *) _04005_ : wt0_actv_data[23:16];
  assign _01202_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16058" *) _04004_ : wt0_actv_data[15:8];
  assign _01291_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16048" *) _04003_ : wt0_actv_data[7:0];
  assign _01319_ = _04002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16038" *) wt0_sd_nan : wt0_actv_nan;
  assign _01320_ = _04001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16028" *) wt0_sd_nz : wt0_actv_nz;
  assign _03157_ = _04000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15994" *) wt_pre_data[1023:1016] : wt7_sd_data[1023:1016];
  assign _03156_ = _03999_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15984" *) wt_pre_data[1015:1008] : wt7_sd_data[1015:1008];
  assign _03155_ = _03998_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15974" *) wt_pre_data[1007:1000] : wt7_sd_data[1007:1000];
  assign _03282_ = _03997_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15964" *) wt_pre_data[999:992] : wt7_sd_data[999:992];
  assign _03281_ = _03996_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15954" *) wt_pre_data[991:984] : wt7_sd_data[991:984];
  assign _03280_ = _03995_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15944" *) wt_pre_data[983:976] : wt7_sd_data[983:976];
  assign _03279_ = _03994_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15934" *) wt_pre_data[975:968] : wt7_sd_data[975:968];
  assign _03278_ = _03993_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15924" *) wt_pre_data[967:960] : wt7_sd_data[967:960];
  assign _03276_ = _03992_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15914" *) wt_pre_data[959:952] : wt7_sd_data[959:952];
  assign _03275_ = _03991_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15904" *) wt_pre_data[951:944] : wt7_sd_data[951:944];
  assign _03274_ = _03990_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15894" *) wt_pre_data[943:936] : wt7_sd_data[943:936];
  assign _03273_ = _03989_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15884" *) wt_pre_data[935:928] : wt7_sd_data[935:928];
  assign _03272_ = _03988_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15874" *) wt_pre_data[927:920] : wt7_sd_data[927:920];
  assign _03271_ = _03987_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15864" *) wt_pre_data[919:912] : wt7_sd_data[919:912];
  assign _03270_ = _03986_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15854" *) wt_pre_data[911:904] : wt7_sd_data[911:904];
  assign _03269_ = _03985_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15844" *) wt_pre_data[903:896] : wt7_sd_data[903:896];
  assign _03268_ = _03984_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15834" *) wt_pre_data[895:888] : wt7_sd_data[895:888];
  assign _03267_ = _03983_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15824" *) wt_pre_data[887:880] : wt7_sd_data[887:880];
  assign _03265_ = _03982_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15814" *) wt_pre_data[879:872] : wt7_sd_data[879:872];
  assign _03264_ = _03981_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15804" *) wt_pre_data[871:864] : wt7_sd_data[871:864];
  assign _03263_ = _03980_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15794" *) wt_pre_data[863:856] : wt7_sd_data[863:856];
  assign _03262_ = _03979_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15784" *) wt_pre_data[855:848] : wt7_sd_data[855:848];
  assign _03261_ = _03978_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15774" *) wt_pre_data[847:840] : wt7_sd_data[847:840];
  assign _03260_ = _03977_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15764" *) wt_pre_data[839:832] : wt7_sd_data[839:832];
  assign _03259_ = _03976_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15754" *) wt_pre_data[831:824] : wt7_sd_data[831:824];
  assign _03258_ = _03975_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15744" *) wt_pre_data[823:816] : wt7_sd_data[823:816];
  assign _03257_ = _03974_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15734" *) wt_pre_data[815:808] : wt7_sd_data[815:808];
  assign _03256_ = _03973_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15724" *) wt_pre_data[807:800] : wt7_sd_data[807:800];
  assign _03253_ = _03972_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15714" *) wt_pre_data[799:792] : wt7_sd_data[799:792];
  assign _03252_ = _03971_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15704" *) wt_pre_data[791:784] : wt7_sd_data[791:784];
  assign _03251_ = _03970_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15694" *) wt_pre_data[783:776] : wt7_sd_data[783:776];
  assign _03250_ = _03969_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15684" *) wt_pre_data[775:768] : wt7_sd_data[775:768];
  assign _03249_ = _03968_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15674" *) wt_pre_data[767:760] : wt7_sd_data[767:760];
  assign _03248_ = _03967_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15664" *) wt_pre_data[759:752] : wt7_sd_data[759:752];
  assign _03247_ = _03966_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15654" *) wt_pre_data[751:744] : wt7_sd_data[751:744];
  assign _03246_ = _03965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15644" *) wt_pre_data[743:736] : wt7_sd_data[743:736];
  assign _03245_ = _03964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15634" *) wt_pre_data[735:728] : wt7_sd_data[735:728];
  assign _03244_ = _03963_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15624" *) wt_pre_data[727:720] : wt7_sd_data[727:720];
  assign _03242_ = _03962_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15614" *) wt_pre_data[719:712] : wt7_sd_data[719:712];
  assign _03241_ = _03961_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15604" *) wt_pre_data[711:704] : wt7_sd_data[711:704];
  assign _03240_ = _03960_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15594" *) wt_pre_data[703:696] : wt7_sd_data[703:696];
  assign _03239_ = _03959_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15584" *) wt_pre_data[695:688] : wt7_sd_data[695:688];
  assign _03238_ = _03958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15574" *) wt_pre_data[687:680] : wt7_sd_data[687:680];
  assign _03237_ = _03957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15564" *) wt_pre_data[679:672] : wt7_sd_data[679:672];
  assign _03236_ = _03956_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15554" *) wt_pre_data[671:664] : wt7_sd_data[671:664];
  assign _03235_ = _03955_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15544" *) wt_pre_data[663:656] : wt7_sd_data[663:656];
  assign _03234_ = _03954_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15534" *) wt_pre_data[655:648] : wt7_sd_data[655:648];
  assign _03233_ = _03953_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15524" *) wt_pre_data[647:640] : wt7_sd_data[647:640];
  assign _03231_ = _03952_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15514" *) wt_pre_data[639:632] : wt7_sd_data[639:632];
  assign _03230_ = _03951_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15504" *) wt_pre_data[631:624] : wt7_sd_data[631:624];
  assign _03229_ = _03950_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15494" *) wt_pre_data[623:616] : wt7_sd_data[623:616];
  assign _03228_ = _03949_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15484" *) wt_pre_data[615:608] : wt7_sd_data[615:608];
  assign _03227_ = _03948_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15474" *) wt_pre_data[607:600] : wt7_sd_data[607:600];
  assign _03226_ = _03947_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15464" *) wt_pre_data[599:592] : wt7_sd_data[599:592];
  assign _03225_ = _03946_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15454" *) wt_pre_data[591:584] : wt7_sd_data[591:584];
  assign _03224_ = _03945_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15444" *) wt_pre_data[583:576] : wt7_sd_data[583:576];
  assign _03223_ = _03944_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15434" *) wt_pre_data[575:568] : wt7_sd_data[575:568];
  assign _03222_ = _03943_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15424" *) wt_pre_data[567:560] : wt7_sd_data[567:560];
  assign _03220_ = _03942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15414" *) wt_pre_data[559:552] : wt7_sd_data[559:552];
  assign _03219_ = _03941_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15404" *) wt_pre_data[551:544] : wt7_sd_data[551:544];
  assign _03218_ = _03940_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15394" *) wt_pre_data[543:536] : wt7_sd_data[543:536];
  assign _03217_ = _03939_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15384" *) wt_pre_data[535:528] : wt7_sd_data[535:528];
  assign _03216_ = _03938_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15374" *) wt_pre_data[527:520] : wt7_sd_data[527:520];
  assign _03215_ = _03937_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15364" *) wt_pre_data[519:512] : wt7_sd_data[519:512];
  assign _03214_ = _03936_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15354" *) wt_pre_data[511:504] : wt7_sd_data[511:504];
  assign _03213_ = _03935_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15344" *) wt_pre_data[503:496] : wt7_sd_data[503:496];
  assign _03212_ = _03934_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15334" *) wt_pre_data[495:488] : wt7_sd_data[495:488];
  assign _03211_ = _03933_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15324" *) wt_pre_data[487:480] : wt7_sd_data[487:480];
  assign _03209_ = _03932_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15314" *) wt_pre_data[479:472] : wt7_sd_data[479:472];
  assign _03208_ = _03931_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15304" *) wt_pre_data[471:464] : wt7_sd_data[471:464];
  assign _03207_ = _03930_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15294" *) wt_pre_data[463:456] : wt7_sd_data[463:456];
  assign _03206_ = _03929_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15284" *) wt_pre_data[455:448] : wt7_sd_data[455:448];
  assign _03205_ = _03928_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15274" *) wt_pre_data[447:440] : wt7_sd_data[447:440];
  assign _03204_ = _03927_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15264" *) wt_pre_data[439:432] : wt7_sd_data[439:432];
  assign _03203_ = _03926_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15254" *) wt_pre_data[431:424] : wt7_sd_data[431:424];
  assign _03202_ = _03925_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15244" *) wt_pre_data[423:416] : wt7_sd_data[423:416];
  assign _03201_ = _03924_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15234" *) wt_pre_data[415:408] : wt7_sd_data[415:408];
  assign _03200_ = _03923_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15224" *) wt_pre_data[407:400] : wt7_sd_data[407:400];
  assign _03198_ = _03922_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15214" *) wt_pre_data[399:392] : wt7_sd_data[399:392];
  assign _03197_ = _03921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15204" *) wt_pre_data[391:384] : wt7_sd_data[391:384];
  assign _03196_ = _03920_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15194" *) wt_pre_data[383:376] : wt7_sd_data[383:376];
  assign _03195_ = _03919_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15184" *) wt_pre_data[375:368] : wt7_sd_data[375:368];
  assign _03194_ = _03918_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15174" *) wt_pre_data[367:360] : wt7_sd_data[367:360];
  assign _03193_ = _03917_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15164" *) wt_pre_data[359:352] : wt7_sd_data[359:352];
  assign _03192_ = _03916_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15154" *) wt_pre_data[351:344] : wt7_sd_data[351:344];
  assign _03191_ = _03915_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15144" *) wt_pre_data[343:336] : wt7_sd_data[343:336];
  assign _03190_ = _03914_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15134" *) wt_pre_data[335:328] : wt7_sd_data[335:328];
  assign _03189_ = _03913_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15124" *) wt_pre_data[327:320] : wt7_sd_data[327:320];
  assign _03187_ = _03912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15114" *) wt_pre_data[319:312] : wt7_sd_data[319:312];
  assign _03186_ = _03911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15104" *) wt_pre_data[311:304] : wt7_sd_data[311:304];
  assign _03185_ = _03910_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15094" *) wt_pre_data[303:296] : wt7_sd_data[303:296];
  assign _03184_ = _03909_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15084" *) wt_pre_data[295:288] : wt7_sd_data[295:288];
  assign _03183_ = _03908_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15074" *) wt_pre_data[287:280] : wt7_sd_data[287:280];
  assign _03182_ = _03907_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15064" *) wt_pre_data[279:272] : wt7_sd_data[279:272];
  assign _03181_ = _03906_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15054" *) wt_pre_data[271:264] : wt7_sd_data[271:264];
  assign _03180_ = _03905_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15044" *) wt_pre_data[263:256] : wt7_sd_data[263:256];
  assign _03179_ = _03904_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15034" *) wt_pre_data[255:248] : wt7_sd_data[255:248];
  assign _03178_ = _03903_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15024" *) wt_pre_data[247:240] : wt7_sd_data[247:240];
  assign _03176_ = _03902_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15014" *) wt_pre_data[239:232] : wt7_sd_data[239:232];
  assign _03175_ = _03901_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:15004" *) wt_pre_data[231:224] : wt7_sd_data[231:224];
  assign _03174_ = _03900_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14994" *) wt_pre_data[223:216] : wt7_sd_data[223:216];
  assign _03173_ = _03899_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14984" *) wt_pre_data[215:208] : wt7_sd_data[215:208];
  assign _03172_ = _03898_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14974" *) wt_pre_data[207:200] : wt7_sd_data[207:200];
  assign _03171_ = _03897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14964" *) wt_pre_data[199:192] : wt7_sd_data[199:192];
  assign _03170_ = _03896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14954" *) wt_pre_data[191:184] : wt7_sd_data[191:184];
  assign _03169_ = _03895_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14944" *) wt_pre_data[183:176] : wt7_sd_data[183:176];
  assign _03168_ = _03894_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14934" *) wt_pre_data[175:168] : wt7_sd_data[175:168];
  assign _03167_ = _03893_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14924" *) wt_pre_data[167:160] : wt7_sd_data[167:160];
  assign _03165_ = _03892_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14914" *) wt_pre_data[159:152] : wt7_sd_data[159:152];
  assign _03164_ = _03891_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14904" *) wt_pre_data[151:144] : wt7_sd_data[151:144];
  assign _03163_ = _03890_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14894" *) wt_pre_data[143:136] : wt7_sd_data[143:136];
  assign _03162_ = _03889_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14884" *) wt_pre_data[135:128] : wt7_sd_data[135:128];
  assign _03161_ = _03888_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14874" *) wt_pre_data[127:120] : wt7_sd_data[127:120];
  assign _03160_ = _03887_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14864" *) wt_pre_data[119:112] : wt7_sd_data[119:112];
  assign _03159_ = _03886_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14854" *) wt_pre_data[111:104] : wt7_sd_data[111:104];
  assign _03158_ = _03885_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14844" *) wt_pre_data[103:96] : wt7_sd_data[103:96];
  assign _03277_ = _03884_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14834" *) wt_pre_data[95:88] : wt7_sd_data[95:88];
  assign _03266_ = _03883_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14824" *) wt_pre_data[87:80] : wt7_sd_data[87:80];
  assign _03254_ = _03882_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14814" *) wt_pre_data[79:72] : wt7_sd_data[79:72];
  assign _03243_ = _03881_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14804" *) wt_pre_data[71:64] : wt7_sd_data[71:64];
  assign _03232_ = _03880_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14794" *) wt_pre_data[63:56] : wt7_sd_data[63:56];
  assign _03221_ = _03879_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14784" *) wt_pre_data[55:48] : wt7_sd_data[55:48];
  assign _03210_ = _03878_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14774" *) wt_pre_data[47:40] : wt7_sd_data[47:40];
  assign _03199_ = _03877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14764" *) wt_pre_data[39:32] : wt7_sd_data[39:32];
  assign _03188_ = _03876_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14754" *) wt_pre_data[31:24] : wt7_sd_data[31:24];
  assign _03177_ = _03875_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14744" *) wt_pre_data[23:16] : wt7_sd_data[23:16];
  assign _03166_ = _03874_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14734" *) wt_pre_data[15:8] : wt7_sd_data[15:8];
  assign _03255_ = _03873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14724" *) wt_pre_data[7:0] : wt7_sd_data[7:0];
  assign _03285_ = _03872_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14714" *) wt_pre_nan : wt7_sd_nan;
  assign _03283_ = _03872_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14704" *) wt_pre_exp : wt7_sd_exp;
  assign _03284_ = _03872_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14694" *) wt_pre_mask : wt7_sd_mask;
  assign _03286_ = wt_pre_sel[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14684" *) wt_pre_nz : wt7_sd_nz;
  assign _02895_ = _03871_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14658" *) wt_pre_data[1023:1016] : wt6_sd_data[1023:1016];
  assign _02894_ = _03870_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14648" *) wt_pre_data[1015:1008] : wt6_sd_data[1015:1008];
  assign _02893_ = _03869_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14638" *) wt_pre_data[1007:1000] : wt6_sd_data[1007:1000];
  assign _03020_ = _03868_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14628" *) wt_pre_data[999:992] : wt6_sd_data[999:992];
  assign _03019_ = _03867_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14618" *) wt_pre_data[991:984] : wt6_sd_data[991:984];
  assign _03018_ = _03866_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14608" *) wt_pre_data[983:976] : wt6_sd_data[983:976];
  assign _03017_ = _03865_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14598" *) wt_pre_data[975:968] : wt6_sd_data[975:968];
  assign _03016_ = _03864_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14588" *) wt_pre_data[967:960] : wt6_sd_data[967:960];
  assign _03014_ = _03863_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14578" *) wt_pre_data[959:952] : wt6_sd_data[959:952];
  assign _03013_ = _03862_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14568" *) wt_pre_data[951:944] : wt6_sd_data[951:944];
  assign _03012_ = _03861_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14558" *) wt_pre_data[943:936] : wt6_sd_data[943:936];
  assign _03011_ = _03860_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14548" *) wt_pre_data[935:928] : wt6_sd_data[935:928];
  assign _03010_ = _03859_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14538" *) wt_pre_data[927:920] : wt6_sd_data[927:920];
  assign _03009_ = _03858_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14528" *) wt_pre_data[919:912] : wt6_sd_data[919:912];
  assign _03008_ = _03857_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14518" *) wt_pre_data[911:904] : wt6_sd_data[911:904];
  assign _03007_ = _03856_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14508" *) wt_pre_data[903:896] : wt6_sd_data[903:896];
  assign _03006_ = _03855_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14498" *) wt_pre_data[895:888] : wt6_sd_data[895:888];
  assign _03005_ = _03854_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14488" *) wt_pre_data[887:880] : wt6_sd_data[887:880];
  assign _03003_ = _03853_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14478" *) wt_pre_data[879:872] : wt6_sd_data[879:872];
  assign _03002_ = _03852_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14468" *) wt_pre_data[871:864] : wt6_sd_data[871:864];
  assign _03001_ = _03851_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14458" *) wt_pre_data[863:856] : wt6_sd_data[863:856];
  assign _03000_ = _03850_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14448" *) wt_pre_data[855:848] : wt6_sd_data[855:848];
  assign _02999_ = _03849_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14438" *) wt_pre_data[847:840] : wt6_sd_data[847:840];
  assign _02998_ = _03848_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14428" *) wt_pre_data[839:832] : wt6_sd_data[839:832];
  assign _02997_ = _03847_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14418" *) wt_pre_data[831:824] : wt6_sd_data[831:824];
  assign _02996_ = _03846_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14408" *) wt_pre_data[823:816] : wt6_sd_data[823:816];
  assign _02995_ = _03845_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14398" *) wt_pre_data[815:808] : wt6_sd_data[815:808];
  assign _02994_ = _03844_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14388" *) wt_pre_data[807:800] : wt6_sd_data[807:800];
  assign _02991_ = _03843_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14378" *) wt_pre_data[799:792] : wt6_sd_data[799:792];
  assign _02990_ = _03842_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14368" *) wt_pre_data[791:784] : wt6_sd_data[791:784];
  assign _02989_ = _03841_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14358" *) wt_pre_data[783:776] : wt6_sd_data[783:776];
  assign _02988_ = _03840_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14348" *) wt_pre_data[775:768] : wt6_sd_data[775:768];
  assign _02987_ = _03839_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14338" *) wt_pre_data[767:760] : wt6_sd_data[767:760];
  assign _02986_ = _03838_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14328" *) wt_pre_data[759:752] : wt6_sd_data[759:752];
  assign _02985_ = _03837_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14318" *) wt_pre_data[751:744] : wt6_sd_data[751:744];
  assign _02984_ = _03836_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14308" *) wt_pre_data[743:736] : wt6_sd_data[743:736];
  assign _02983_ = _03835_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14298" *) wt_pre_data[735:728] : wt6_sd_data[735:728];
  assign _02982_ = _03834_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14288" *) wt_pre_data[727:720] : wt6_sd_data[727:720];
  assign _02980_ = _03833_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14278" *) wt_pre_data[719:712] : wt6_sd_data[719:712];
  assign _02979_ = _03832_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14268" *) wt_pre_data[711:704] : wt6_sd_data[711:704];
  assign _02978_ = _03831_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14258" *) wt_pre_data[703:696] : wt6_sd_data[703:696];
  assign _02977_ = _03830_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14248" *) wt_pre_data[695:688] : wt6_sd_data[695:688];
  assign _02976_ = _03829_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14238" *) wt_pre_data[687:680] : wt6_sd_data[687:680];
  assign _02975_ = _03828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14228" *) wt_pre_data[679:672] : wt6_sd_data[679:672];
  assign _02974_ = _03827_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14218" *) wt_pre_data[671:664] : wt6_sd_data[671:664];
  assign _02973_ = _03826_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14208" *) wt_pre_data[663:656] : wt6_sd_data[663:656];
  assign _02972_ = _03825_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14198" *) wt_pre_data[655:648] : wt6_sd_data[655:648];
  assign _02971_ = _03824_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14188" *) wt_pre_data[647:640] : wt6_sd_data[647:640];
  assign _02969_ = _03823_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14178" *) wt_pre_data[639:632] : wt6_sd_data[639:632];
  assign _02968_ = _03822_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14168" *) wt_pre_data[631:624] : wt6_sd_data[631:624];
  assign _02967_ = _03821_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14158" *) wt_pre_data[623:616] : wt6_sd_data[623:616];
  assign _02966_ = _03820_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14148" *) wt_pre_data[615:608] : wt6_sd_data[615:608];
  assign _02965_ = _03819_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14138" *) wt_pre_data[607:600] : wt6_sd_data[607:600];
  assign _02964_ = _03818_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14128" *) wt_pre_data[599:592] : wt6_sd_data[599:592];
  assign _02963_ = _03817_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14118" *) wt_pre_data[591:584] : wt6_sd_data[591:584];
  assign _02962_ = _03816_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14108" *) wt_pre_data[583:576] : wt6_sd_data[583:576];
  assign _02961_ = _03815_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14098" *) wt_pre_data[575:568] : wt6_sd_data[575:568];
  assign _02960_ = _03814_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14088" *) wt_pre_data[567:560] : wt6_sd_data[567:560];
  assign _02958_ = _03813_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14078" *) wt_pre_data[559:552] : wt6_sd_data[559:552];
  assign _02957_ = _03812_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14068" *) wt_pre_data[551:544] : wt6_sd_data[551:544];
  assign _02956_ = _03811_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14058" *) wt_pre_data[543:536] : wt6_sd_data[543:536];
  assign _02955_ = _03810_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14048" *) wt_pre_data[535:528] : wt6_sd_data[535:528];
  assign _02954_ = _03809_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14038" *) wt_pre_data[527:520] : wt6_sd_data[527:520];
  assign _02953_ = _03808_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14028" *) wt_pre_data[519:512] : wt6_sd_data[519:512];
  assign _02952_ = _03807_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14018" *) wt_pre_data[511:504] : wt6_sd_data[511:504];
  assign _02951_ = _03806_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14008" *) wt_pre_data[503:496] : wt6_sd_data[503:496];
  assign _02950_ = _03805_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13998" *) wt_pre_data[495:488] : wt6_sd_data[495:488];
  assign _02949_ = _03804_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13988" *) wt_pre_data[487:480] : wt6_sd_data[487:480];
  assign _02947_ = _03803_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13978" *) wt_pre_data[479:472] : wt6_sd_data[479:472];
  assign _02946_ = _03802_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13968" *) wt_pre_data[471:464] : wt6_sd_data[471:464];
  assign _02945_ = _03801_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13958" *) wt_pre_data[463:456] : wt6_sd_data[463:456];
  assign _02944_ = _03800_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13948" *) wt_pre_data[455:448] : wt6_sd_data[455:448];
  assign _02943_ = _03799_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13938" *) wt_pre_data[447:440] : wt6_sd_data[447:440];
  assign _02942_ = _03798_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13928" *) wt_pre_data[439:432] : wt6_sd_data[439:432];
  assign _02941_ = _03797_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13918" *) wt_pre_data[431:424] : wt6_sd_data[431:424];
  assign _02940_ = _03796_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13908" *) wt_pre_data[423:416] : wt6_sd_data[423:416];
  assign _02939_ = _03795_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13898" *) wt_pre_data[415:408] : wt6_sd_data[415:408];
  assign _02938_ = _03794_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13888" *) wt_pre_data[407:400] : wt6_sd_data[407:400];
  assign _02936_ = _03793_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13878" *) wt_pre_data[399:392] : wt6_sd_data[399:392];
  assign _02935_ = _03792_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13868" *) wt_pre_data[391:384] : wt6_sd_data[391:384];
  assign _02934_ = _03791_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13858" *) wt_pre_data[383:376] : wt6_sd_data[383:376];
  assign _02933_ = _03790_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13848" *) wt_pre_data[375:368] : wt6_sd_data[375:368];
  assign _02932_ = _03789_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13838" *) wt_pre_data[367:360] : wt6_sd_data[367:360];
  assign _02931_ = _03788_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13828" *) wt_pre_data[359:352] : wt6_sd_data[359:352];
  assign _02930_ = _03787_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13818" *) wt_pre_data[351:344] : wt6_sd_data[351:344];
  assign _02929_ = _03786_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13808" *) wt_pre_data[343:336] : wt6_sd_data[343:336];
  assign _02928_ = _03785_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13798" *) wt_pre_data[335:328] : wt6_sd_data[335:328];
  assign _02927_ = _03784_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13788" *) wt_pre_data[327:320] : wt6_sd_data[327:320];
  assign _02925_ = _03783_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13778" *) wt_pre_data[319:312] : wt6_sd_data[319:312];
  assign _02924_ = _03782_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13768" *) wt_pre_data[311:304] : wt6_sd_data[311:304];
  assign _02923_ = _03781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13758" *) wt_pre_data[303:296] : wt6_sd_data[303:296];
  assign _02922_ = _03780_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13748" *) wt_pre_data[295:288] : wt6_sd_data[295:288];
  assign _02921_ = _03779_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13738" *) wt_pre_data[287:280] : wt6_sd_data[287:280];
  assign _02920_ = _03778_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13728" *) wt_pre_data[279:272] : wt6_sd_data[279:272];
  assign _02919_ = _03777_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13718" *) wt_pre_data[271:264] : wt6_sd_data[271:264];
  assign _02918_ = _03776_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13708" *) wt_pre_data[263:256] : wt6_sd_data[263:256];
  assign _02917_ = _03775_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13698" *) wt_pre_data[255:248] : wt6_sd_data[255:248];
  assign _02916_ = _03774_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13688" *) wt_pre_data[247:240] : wt6_sd_data[247:240];
  assign _02914_ = _03773_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13678" *) wt_pre_data[239:232] : wt6_sd_data[239:232];
  assign _02913_ = _03772_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13668" *) wt_pre_data[231:224] : wt6_sd_data[231:224];
  assign _02912_ = _03771_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13658" *) wt_pre_data[223:216] : wt6_sd_data[223:216];
  assign _02911_ = _03770_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13648" *) wt_pre_data[215:208] : wt6_sd_data[215:208];
  assign _02910_ = _03769_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13638" *) wt_pre_data[207:200] : wt6_sd_data[207:200];
  assign _02909_ = _03768_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13628" *) wt_pre_data[199:192] : wt6_sd_data[199:192];
  assign _02908_ = _03767_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13618" *) wt_pre_data[191:184] : wt6_sd_data[191:184];
  assign _02907_ = _03766_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13608" *) wt_pre_data[183:176] : wt6_sd_data[183:176];
  assign _02906_ = _03765_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13598" *) wt_pre_data[175:168] : wt6_sd_data[175:168];
  assign _02905_ = _03764_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13588" *) wt_pre_data[167:160] : wt6_sd_data[167:160];
  assign _02903_ = _03763_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13578" *) wt_pre_data[159:152] : wt6_sd_data[159:152];
  assign _02902_ = _03762_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13568" *) wt_pre_data[151:144] : wt6_sd_data[151:144];
  assign _02901_ = _03761_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13558" *) wt_pre_data[143:136] : wt6_sd_data[143:136];
  assign _02900_ = _03760_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13548" *) wt_pre_data[135:128] : wt6_sd_data[135:128];
  assign _02899_ = _03759_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13538" *) wt_pre_data[127:120] : wt6_sd_data[127:120];
  assign _02898_ = _03758_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13528" *) wt_pre_data[119:112] : wt6_sd_data[119:112];
  assign _02897_ = _03757_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13518" *) wt_pre_data[111:104] : wt6_sd_data[111:104];
  assign _02896_ = _03756_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13508" *) wt_pre_data[103:96] : wt6_sd_data[103:96];
  assign _03015_ = _03755_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13498" *) wt_pre_data[95:88] : wt6_sd_data[95:88];
  assign _03004_ = _03754_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13488" *) wt_pre_data[87:80] : wt6_sd_data[87:80];
  assign _02992_ = _03753_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13478" *) wt_pre_data[79:72] : wt6_sd_data[79:72];
  assign _02981_ = _03752_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13468" *) wt_pre_data[71:64] : wt6_sd_data[71:64];
  assign _02970_ = _03751_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13458" *) wt_pre_data[63:56] : wt6_sd_data[63:56];
  assign _02959_ = _03750_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13448" *) wt_pre_data[55:48] : wt6_sd_data[55:48];
  assign _02948_ = _03749_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13438" *) wt_pre_data[47:40] : wt6_sd_data[47:40];
  assign _02937_ = _03748_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13428" *) wt_pre_data[39:32] : wt6_sd_data[39:32];
  assign _02926_ = _03747_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13418" *) wt_pre_data[31:24] : wt6_sd_data[31:24];
  assign _02915_ = _03746_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13408" *) wt_pre_data[23:16] : wt6_sd_data[23:16];
  assign _02904_ = _03745_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13398" *) wt_pre_data[15:8] : wt6_sd_data[15:8];
  assign _02993_ = _03744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13388" *) wt_pre_data[7:0] : wt6_sd_data[7:0];
  assign _03023_ = _03743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13378" *) wt_pre_nan : wt6_sd_nan;
  assign _03021_ = _03743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13368" *) wt_pre_exp : wt6_sd_exp;
  assign _03022_ = _03743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13358" *) wt_pre_mask : wt6_sd_mask;
  assign _03024_ = wt_pre_sel[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13348" *) wt_pre_nz : wt6_sd_nz;
  assign _02633_ = _03742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13322" *) wt_pre_data[1023:1016] : wt5_sd_data[1023:1016];
  assign _02632_ = _03741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13312" *) wt_pre_data[1015:1008] : wt5_sd_data[1015:1008];
  assign _02631_ = _03740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13302" *) wt_pre_data[1007:1000] : wt5_sd_data[1007:1000];
  assign _02758_ = _03739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13292" *) wt_pre_data[999:992] : wt5_sd_data[999:992];
  assign _02757_ = _03738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13282" *) wt_pre_data[991:984] : wt5_sd_data[991:984];
  assign _02756_ = _03737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13272" *) wt_pre_data[983:976] : wt5_sd_data[983:976];
  assign _02755_ = _03736_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13262" *) wt_pre_data[975:968] : wt5_sd_data[975:968];
  assign _02754_ = _03735_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13252" *) wt_pre_data[967:960] : wt5_sd_data[967:960];
  assign _02752_ = _03734_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13242" *) wt_pre_data[959:952] : wt5_sd_data[959:952];
  assign _02751_ = _03733_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13232" *) wt_pre_data[951:944] : wt5_sd_data[951:944];
  assign _02750_ = _03732_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13222" *) wt_pre_data[943:936] : wt5_sd_data[943:936];
  assign _02749_ = _03731_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13212" *) wt_pre_data[935:928] : wt5_sd_data[935:928];
  assign _02748_ = _03730_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13202" *) wt_pre_data[927:920] : wt5_sd_data[927:920];
  assign _02747_ = _03729_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13192" *) wt_pre_data[919:912] : wt5_sd_data[919:912];
  assign _02746_ = _03728_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13182" *) wt_pre_data[911:904] : wt5_sd_data[911:904];
  assign _02745_ = _03727_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13172" *) wt_pre_data[903:896] : wt5_sd_data[903:896];
  assign _02744_ = _03726_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13162" *) wt_pre_data[895:888] : wt5_sd_data[895:888];
  assign _02743_ = _03725_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13152" *) wt_pre_data[887:880] : wt5_sd_data[887:880];
  assign _02741_ = _03724_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13142" *) wt_pre_data[879:872] : wt5_sd_data[879:872];
  assign _02740_ = _03723_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13132" *) wt_pre_data[871:864] : wt5_sd_data[871:864];
  assign _02739_ = _03722_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13122" *) wt_pre_data[863:856] : wt5_sd_data[863:856];
  assign _02738_ = _03721_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13112" *) wt_pre_data[855:848] : wt5_sd_data[855:848];
  assign _02737_ = _03720_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13102" *) wt_pre_data[847:840] : wt5_sd_data[847:840];
  assign _02736_ = _03719_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13092" *) wt_pre_data[839:832] : wt5_sd_data[839:832];
  assign _02735_ = _03718_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13082" *) wt_pre_data[831:824] : wt5_sd_data[831:824];
  assign _02734_ = _03717_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13072" *) wt_pre_data[823:816] : wt5_sd_data[823:816];
  assign _02733_ = _03716_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13062" *) wt_pre_data[815:808] : wt5_sd_data[815:808];
  assign _02732_ = _03715_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13052" *) wt_pre_data[807:800] : wt5_sd_data[807:800];
  assign _02729_ = _03714_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13042" *) wt_pre_data[799:792] : wt5_sd_data[799:792];
  assign _02728_ = _03713_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13032" *) wt_pre_data[791:784] : wt5_sd_data[791:784];
  assign _02727_ = _03712_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13022" *) wt_pre_data[783:776] : wt5_sd_data[783:776];
  assign _02726_ = _03711_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13012" *) wt_pre_data[775:768] : wt5_sd_data[775:768];
  assign _02725_ = _03710_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13002" *) wt_pre_data[767:760] : wt5_sd_data[767:760];
  assign _02724_ = _03709_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12992" *) wt_pre_data[759:752] : wt5_sd_data[759:752];
  assign _02723_ = _03708_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12982" *) wt_pre_data[751:744] : wt5_sd_data[751:744];
  assign _02722_ = _03707_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12972" *) wt_pre_data[743:736] : wt5_sd_data[743:736];
  assign _02721_ = _03706_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12962" *) wt_pre_data[735:728] : wt5_sd_data[735:728];
  assign _02720_ = _03705_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12952" *) wt_pre_data[727:720] : wt5_sd_data[727:720];
  assign _02718_ = _03704_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12942" *) wt_pre_data[719:712] : wt5_sd_data[719:712];
  assign _02717_ = _03703_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12932" *) wt_pre_data[711:704] : wt5_sd_data[711:704];
  assign _02716_ = _03702_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12922" *) wt_pre_data[703:696] : wt5_sd_data[703:696];
  assign _02715_ = _03701_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12912" *) wt_pre_data[695:688] : wt5_sd_data[695:688];
  assign _02714_ = _03700_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12902" *) wt_pre_data[687:680] : wt5_sd_data[687:680];
  assign _02713_ = _03699_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12892" *) wt_pre_data[679:672] : wt5_sd_data[679:672];
  assign _02712_ = _03698_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12882" *) wt_pre_data[671:664] : wt5_sd_data[671:664];
  assign _02711_ = _03697_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12872" *) wt_pre_data[663:656] : wt5_sd_data[663:656];
  assign _02710_ = _03696_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12862" *) wt_pre_data[655:648] : wt5_sd_data[655:648];
  assign _02709_ = _03695_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12852" *) wt_pre_data[647:640] : wt5_sd_data[647:640];
  assign _02707_ = _03694_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12842" *) wt_pre_data[639:632] : wt5_sd_data[639:632];
  assign _02706_ = _03693_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12832" *) wt_pre_data[631:624] : wt5_sd_data[631:624];
  assign _02705_ = _03692_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12822" *) wt_pre_data[623:616] : wt5_sd_data[623:616];
  assign _02704_ = _03691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12812" *) wt_pre_data[615:608] : wt5_sd_data[615:608];
  assign _02703_ = _03690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12802" *) wt_pre_data[607:600] : wt5_sd_data[607:600];
  assign _02702_ = _03689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12792" *) wt_pre_data[599:592] : wt5_sd_data[599:592];
  assign _02701_ = _03688_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12782" *) wt_pre_data[591:584] : wt5_sd_data[591:584];
  assign _02700_ = _03687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12772" *) wt_pre_data[583:576] : wt5_sd_data[583:576];
  assign _02699_ = _03686_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12762" *) wt_pre_data[575:568] : wt5_sd_data[575:568];
  assign _02698_ = _03685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12752" *) wt_pre_data[567:560] : wt5_sd_data[567:560];
  assign _02696_ = _03684_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12742" *) wt_pre_data[559:552] : wt5_sd_data[559:552];
  assign _02695_ = _03683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12732" *) wt_pre_data[551:544] : wt5_sd_data[551:544];
  assign _02694_ = _03682_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12722" *) wt_pre_data[543:536] : wt5_sd_data[543:536];
  assign _02693_ = _03681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12712" *) wt_pre_data[535:528] : wt5_sd_data[535:528];
  assign _02692_ = _03680_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12702" *) wt_pre_data[527:520] : wt5_sd_data[527:520];
  assign _02691_ = _03679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12692" *) wt_pre_data[519:512] : wt5_sd_data[519:512];
  assign _02690_ = _03678_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12682" *) wt_pre_data[511:504] : wt5_sd_data[511:504];
  assign _02689_ = _03677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12672" *) wt_pre_data[503:496] : wt5_sd_data[503:496];
  assign _02688_ = _03676_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12662" *) wt_pre_data[495:488] : wt5_sd_data[495:488];
  assign _02687_ = _03675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12652" *) wt_pre_data[487:480] : wt5_sd_data[487:480];
  assign _02685_ = _03674_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12642" *) wt_pre_data[479:472] : wt5_sd_data[479:472];
  assign _02684_ = _03673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12632" *) wt_pre_data[471:464] : wt5_sd_data[471:464];
  assign _02683_ = _03672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12622" *) wt_pre_data[463:456] : wt5_sd_data[463:456];
  assign _02682_ = _03671_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12612" *) wt_pre_data[455:448] : wt5_sd_data[455:448];
  assign _02681_ = _03670_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12602" *) wt_pre_data[447:440] : wt5_sd_data[447:440];
  assign _02680_ = _03669_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12592" *) wt_pre_data[439:432] : wt5_sd_data[439:432];
  assign _02679_ = _03668_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12582" *) wt_pre_data[431:424] : wt5_sd_data[431:424];
  assign _02678_ = _03667_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12572" *) wt_pre_data[423:416] : wt5_sd_data[423:416];
  assign _02677_ = _03666_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12562" *) wt_pre_data[415:408] : wt5_sd_data[415:408];
  assign _02676_ = _03665_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12552" *) wt_pre_data[407:400] : wt5_sd_data[407:400];
  assign _02674_ = _03664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12542" *) wt_pre_data[399:392] : wt5_sd_data[399:392];
  assign _02673_ = _03663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12532" *) wt_pre_data[391:384] : wt5_sd_data[391:384];
  assign _02672_ = _03662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12522" *) wt_pre_data[383:376] : wt5_sd_data[383:376];
  assign _02671_ = _03661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12512" *) wt_pre_data[375:368] : wt5_sd_data[375:368];
  assign _02670_ = _03660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12502" *) wt_pre_data[367:360] : wt5_sd_data[367:360];
  assign _02669_ = _03659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12492" *) wt_pre_data[359:352] : wt5_sd_data[359:352];
  assign _02668_ = _03658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12482" *) wt_pre_data[351:344] : wt5_sd_data[351:344];
  assign _02667_ = _03657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12472" *) wt_pre_data[343:336] : wt5_sd_data[343:336];
  assign _02666_ = _03656_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12462" *) wt_pre_data[335:328] : wt5_sd_data[335:328];
  assign _02665_ = _03655_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12452" *) wt_pre_data[327:320] : wt5_sd_data[327:320];
  assign _02663_ = _03654_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12442" *) wt_pre_data[319:312] : wt5_sd_data[319:312];
  assign _02662_ = _03653_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12432" *) wt_pre_data[311:304] : wt5_sd_data[311:304];
  assign _02661_ = _03652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12422" *) wt_pre_data[303:296] : wt5_sd_data[303:296];
  assign _02660_ = _03651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12412" *) wt_pre_data[295:288] : wt5_sd_data[295:288];
  assign _02659_ = _03650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12402" *) wt_pre_data[287:280] : wt5_sd_data[287:280];
  assign _02658_ = _03649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12392" *) wt_pre_data[279:272] : wt5_sd_data[279:272];
  assign _02657_ = _03648_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12382" *) wt_pre_data[271:264] : wt5_sd_data[271:264];
  assign _02656_ = _03647_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12372" *) wt_pre_data[263:256] : wt5_sd_data[263:256];
  assign _02655_ = _03646_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12362" *) wt_pre_data[255:248] : wt5_sd_data[255:248];
  assign _02654_ = _03645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12352" *) wt_pre_data[247:240] : wt5_sd_data[247:240];
  assign _02652_ = _03644_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12342" *) wt_pre_data[239:232] : wt5_sd_data[239:232];
  assign _02651_ = _03643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12332" *) wt_pre_data[231:224] : wt5_sd_data[231:224];
  assign _02650_ = _03642_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12322" *) wt_pre_data[223:216] : wt5_sd_data[223:216];
  assign _02649_ = _03641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12312" *) wt_pre_data[215:208] : wt5_sd_data[215:208];
  assign _02648_ = _03640_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12302" *) wt_pre_data[207:200] : wt5_sd_data[207:200];
  assign _02647_ = _03639_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12292" *) wt_pre_data[199:192] : wt5_sd_data[199:192];
  assign _02646_ = _03638_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12282" *) wt_pre_data[191:184] : wt5_sd_data[191:184];
  assign _02645_ = _03637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12272" *) wt_pre_data[183:176] : wt5_sd_data[183:176];
  assign _02644_ = _03636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12262" *) wt_pre_data[175:168] : wt5_sd_data[175:168];
  assign _02643_ = _03635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12252" *) wt_pre_data[167:160] : wt5_sd_data[167:160];
  assign _02641_ = _03634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12242" *) wt_pre_data[159:152] : wt5_sd_data[159:152];
  assign _02640_ = _03633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12232" *) wt_pre_data[151:144] : wt5_sd_data[151:144];
  assign _02639_ = _03632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12222" *) wt_pre_data[143:136] : wt5_sd_data[143:136];
  assign _02638_ = _03631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12212" *) wt_pre_data[135:128] : wt5_sd_data[135:128];
  assign _02637_ = _03630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12202" *) wt_pre_data[127:120] : wt5_sd_data[127:120];
  assign _02636_ = _03629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12192" *) wt_pre_data[119:112] : wt5_sd_data[119:112];
  assign _02635_ = _03628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12182" *) wt_pre_data[111:104] : wt5_sd_data[111:104];
  assign _02634_ = _03627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12172" *) wt_pre_data[103:96] : wt5_sd_data[103:96];
  assign _02753_ = _03626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12162" *) wt_pre_data[95:88] : wt5_sd_data[95:88];
  assign _02742_ = _03625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12152" *) wt_pre_data[87:80] : wt5_sd_data[87:80];
  assign _02730_ = _03624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12142" *) wt_pre_data[79:72] : wt5_sd_data[79:72];
  assign _02719_ = _03623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12132" *) wt_pre_data[71:64] : wt5_sd_data[71:64];
  assign _02708_ = _03622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12122" *) wt_pre_data[63:56] : wt5_sd_data[63:56];
  assign _02697_ = _03621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12112" *) wt_pre_data[55:48] : wt5_sd_data[55:48];
  assign _02686_ = _03620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12102" *) wt_pre_data[47:40] : wt5_sd_data[47:40];
  assign _02675_ = _03619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12092" *) wt_pre_data[39:32] : wt5_sd_data[39:32];
  assign _02664_ = _03618_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12082" *) wt_pre_data[31:24] : wt5_sd_data[31:24];
  assign _02653_ = _03617_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12072" *) wt_pre_data[23:16] : wt5_sd_data[23:16];
  assign _02642_ = _03616_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12062" *) wt_pre_data[15:8] : wt5_sd_data[15:8];
  assign _02731_ = _03615_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12052" *) wt_pre_data[7:0] : wt5_sd_data[7:0];
  assign _02761_ = _03614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12042" *) wt_pre_nan : wt5_sd_nan;
  assign _02759_ = _03614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12032" *) wt_pre_exp : wt5_sd_exp;
  assign _02760_ = _03614_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12022" *) wt_pre_mask : wt5_sd_mask;
  assign _02762_ = wt_pre_sel[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12012" *) wt_pre_nz : wt5_sd_nz;
  assign _02371_ = _03613_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11986" *) wt_pre_data[1023:1016] : wt4_sd_data[1023:1016];
  assign _02370_ = _03612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11976" *) wt_pre_data[1015:1008] : wt4_sd_data[1015:1008];
  assign _02369_ = _03611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11966" *) wt_pre_data[1007:1000] : wt4_sd_data[1007:1000];
  assign _02496_ = _03610_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11956" *) wt_pre_data[999:992] : wt4_sd_data[999:992];
  assign _02495_ = _03609_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11946" *) wt_pre_data[991:984] : wt4_sd_data[991:984];
  assign _02494_ = _03608_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11936" *) wt_pre_data[983:976] : wt4_sd_data[983:976];
  assign _02493_ = _03607_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11926" *) wt_pre_data[975:968] : wt4_sd_data[975:968];
  assign _02492_ = _03606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11916" *) wt_pre_data[967:960] : wt4_sd_data[967:960];
  assign _02490_ = _03605_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11906" *) wt_pre_data[959:952] : wt4_sd_data[959:952];
  assign _02489_ = _03604_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11896" *) wt_pre_data[951:944] : wt4_sd_data[951:944];
  assign _02488_ = _03603_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11886" *) wt_pre_data[943:936] : wt4_sd_data[943:936];
  assign _02487_ = _03602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11876" *) wt_pre_data[935:928] : wt4_sd_data[935:928];
  assign _02486_ = _03601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11866" *) wt_pre_data[927:920] : wt4_sd_data[927:920];
  assign _02485_ = _03600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11856" *) wt_pre_data[919:912] : wt4_sd_data[919:912];
  assign _02484_ = _03599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11846" *) wt_pre_data[911:904] : wt4_sd_data[911:904];
  assign _02483_ = _03598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11836" *) wt_pre_data[903:896] : wt4_sd_data[903:896];
  assign _02482_ = _03597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11826" *) wt_pre_data[895:888] : wt4_sd_data[895:888];
  assign _02481_ = _03596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11816" *) wt_pre_data[887:880] : wt4_sd_data[887:880];
  assign _02479_ = _03595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11806" *) wt_pre_data[879:872] : wt4_sd_data[879:872];
  assign _02478_ = _03594_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11796" *) wt_pre_data[871:864] : wt4_sd_data[871:864];
  assign _02477_ = _03593_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11786" *) wt_pre_data[863:856] : wt4_sd_data[863:856];
  assign _02476_ = _03592_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11776" *) wt_pre_data[855:848] : wt4_sd_data[855:848];
  assign _02475_ = _03591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11766" *) wt_pre_data[847:840] : wt4_sd_data[847:840];
  assign _02474_ = _03590_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11756" *) wt_pre_data[839:832] : wt4_sd_data[839:832];
  assign _02473_ = _03589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11746" *) wt_pre_data[831:824] : wt4_sd_data[831:824];
  assign _02472_ = _03588_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11736" *) wt_pre_data[823:816] : wt4_sd_data[823:816];
  assign _02471_ = _03587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11726" *) wt_pre_data[815:808] : wt4_sd_data[815:808];
  assign _02470_ = _03586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11716" *) wt_pre_data[807:800] : wt4_sd_data[807:800];
  assign _02467_ = _03585_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11706" *) wt_pre_data[799:792] : wt4_sd_data[799:792];
  assign _02466_ = _03584_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11696" *) wt_pre_data[791:784] : wt4_sd_data[791:784];
  assign _02465_ = _03583_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11686" *) wt_pre_data[783:776] : wt4_sd_data[783:776];
  assign _02464_ = _03582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11676" *) wt_pre_data[775:768] : wt4_sd_data[775:768];
  assign _02463_ = _03581_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11666" *) wt_pre_data[767:760] : wt4_sd_data[767:760];
  assign _02462_ = _03580_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11656" *) wt_pre_data[759:752] : wt4_sd_data[759:752];
  assign _02461_ = _03579_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11646" *) wt_pre_data[751:744] : wt4_sd_data[751:744];
  assign _02460_ = _03578_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11636" *) wt_pre_data[743:736] : wt4_sd_data[743:736];
  assign _02459_ = _03577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11626" *) wt_pre_data[735:728] : wt4_sd_data[735:728];
  assign _02458_ = _03576_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11616" *) wt_pre_data[727:720] : wt4_sd_data[727:720];
  assign _02456_ = _03575_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11606" *) wt_pre_data[719:712] : wt4_sd_data[719:712];
  assign _02455_ = _03574_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11596" *) wt_pre_data[711:704] : wt4_sd_data[711:704];
  assign _02454_ = _03573_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11586" *) wt_pre_data[703:696] : wt4_sd_data[703:696];
  assign _02453_ = _03572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11576" *) wt_pre_data[695:688] : wt4_sd_data[695:688];
  assign _02452_ = _03571_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11566" *) wt_pre_data[687:680] : wt4_sd_data[687:680];
  assign _02451_ = _03570_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11556" *) wt_pre_data[679:672] : wt4_sd_data[679:672];
  assign _02450_ = _03569_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11546" *) wt_pre_data[671:664] : wt4_sd_data[671:664];
  assign _02449_ = _03568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11536" *) wt_pre_data[663:656] : wt4_sd_data[663:656];
  assign _02448_ = _03567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11526" *) wt_pre_data[655:648] : wt4_sd_data[655:648];
  assign _02447_ = _03566_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11516" *) wt_pre_data[647:640] : wt4_sd_data[647:640];
  assign _02445_ = _03565_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11506" *) wt_pre_data[639:632] : wt4_sd_data[639:632];
  assign _02444_ = _03564_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11496" *) wt_pre_data[631:624] : wt4_sd_data[631:624];
  assign _02443_ = _03563_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11486" *) wt_pre_data[623:616] : wt4_sd_data[623:616];
  assign _02442_ = _03562_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11476" *) wt_pre_data[615:608] : wt4_sd_data[615:608];
  assign _02441_ = _03561_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11466" *) wt_pre_data[607:600] : wt4_sd_data[607:600];
  assign _02440_ = _03560_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11456" *) wt_pre_data[599:592] : wt4_sd_data[599:592];
  assign _02439_ = _03559_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11446" *) wt_pre_data[591:584] : wt4_sd_data[591:584];
  assign _02438_ = _03558_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11436" *) wt_pre_data[583:576] : wt4_sd_data[583:576];
  assign _02437_ = _03557_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11426" *) wt_pre_data[575:568] : wt4_sd_data[575:568];
  assign _02436_ = _03556_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11416" *) wt_pre_data[567:560] : wt4_sd_data[567:560];
  assign _02434_ = _03555_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11406" *) wt_pre_data[559:552] : wt4_sd_data[559:552];
  assign _02433_ = _03554_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11396" *) wt_pre_data[551:544] : wt4_sd_data[551:544];
  assign _02432_ = _03553_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11386" *) wt_pre_data[543:536] : wt4_sd_data[543:536];
  assign _02431_ = _03552_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11376" *) wt_pre_data[535:528] : wt4_sd_data[535:528];
  assign _02430_ = _03551_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11366" *) wt_pre_data[527:520] : wt4_sd_data[527:520];
  assign _02429_ = _03550_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11356" *) wt_pre_data[519:512] : wt4_sd_data[519:512];
  assign _02428_ = _03549_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11346" *) wt_pre_data[511:504] : wt4_sd_data[511:504];
  assign _02427_ = _03548_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11336" *) wt_pre_data[503:496] : wt4_sd_data[503:496];
  assign _02426_ = _03547_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11326" *) wt_pre_data[495:488] : wt4_sd_data[495:488];
  assign _02425_ = _03546_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11316" *) wt_pre_data[487:480] : wt4_sd_data[487:480];
  assign _02423_ = _03545_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11306" *) wt_pre_data[479:472] : wt4_sd_data[479:472];
  assign _02422_ = _03544_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11296" *) wt_pre_data[471:464] : wt4_sd_data[471:464];
  assign _02421_ = _03543_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11286" *) wt_pre_data[463:456] : wt4_sd_data[463:456];
  assign _02420_ = _03542_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11276" *) wt_pre_data[455:448] : wt4_sd_data[455:448];
  assign _02419_ = _03541_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11266" *) wt_pre_data[447:440] : wt4_sd_data[447:440];
  assign _02418_ = _03540_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11256" *) wt_pre_data[439:432] : wt4_sd_data[439:432];
  assign _02417_ = _03539_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11246" *) wt_pre_data[431:424] : wt4_sd_data[431:424];
  assign _02416_ = _03538_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11236" *) wt_pre_data[423:416] : wt4_sd_data[423:416];
  assign _02415_ = _03537_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11226" *) wt_pre_data[415:408] : wt4_sd_data[415:408];
  assign _02414_ = _03536_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11216" *) wt_pre_data[407:400] : wt4_sd_data[407:400];
  assign _02412_ = _03535_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11206" *) wt_pre_data[399:392] : wt4_sd_data[399:392];
  assign _02411_ = _03534_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11196" *) wt_pre_data[391:384] : wt4_sd_data[391:384];
  assign _02410_ = _03533_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11186" *) wt_pre_data[383:376] : wt4_sd_data[383:376];
  assign _02409_ = _03532_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11176" *) wt_pre_data[375:368] : wt4_sd_data[375:368];
  assign _02408_ = _03531_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11166" *) wt_pre_data[367:360] : wt4_sd_data[367:360];
  assign _02407_ = _03530_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11156" *) wt_pre_data[359:352] : wt4_sd_data[359:352];
  assign _02406_ = _03529_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11146" *) wt_pre_data[351:344] : wt4_sd_data[351:344];
  assign _02405_ = _03528_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11136" *) wt_pre_data[343:336] : wt4_sd_data[343:336];
  assign _02404_ = _03527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11126" *) wt_pre_data[335:328] : wt4_sd_data[335:328];
  assign _02403_ = _03526_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11116" *) wt_pre_data[327:320] : wt4_sd_data[327:320];
  assign _02401_ = _03525_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11106" *) wt_pre_data[319:312] : wt4_sd_data[319:312];
  assign _02400_ = _03524_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11096" *) wt_pre_data[311:304] : wt4_sd_data[311:304];
  assign _02399_ = _03523_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11086" *) wt_pre_data[303:296] : wt4_sd_data[303:296];
  assign _02398_ = _03522_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11076" *) wt_pre_data[295:288] : wt4_sd_data[295:288];
  assign _02397_ = _03521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11066" *) wt_pre_data[287:280] : wt4_sd_data[287:280];
  assign _02396_ = _03520_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11056" *) wt_pre_data[279:272] : wt4_sd_data[279:272];
  assign _02395_ = _03519_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11046" *) wt_pre_data[271:264] : wt4_sd_data[271:264];
  assign _02394_ = _03518_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11036" *) wt_pre_data[263:256] : wt4_sd_data[263:256];
  assign _02393_ = _03517_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11026" *) wt_pre_data[255:248] : wt4_sd_data[255:248];
  assign _02392_ = _03516_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11016" *) wt_pre_data[247:240] : wt4_sd_data[247:240];
  assign _02390_ = _03515_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:11006" *) wt_pre_data[239:232] : wt4_sd_data[239:232];
  assign _02389_ = _03514_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10996" *) wt_pre_data[231:224] : wt4_sd_data[231:224];
  assign _02388_ = _03513_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10986" *) wt_pre_data[223:216] : wt4_sd_data[223:216];
  assign _02387_ = _03512_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10976" *) wt_pre_data[215:208] : wt4_sd_data[215:208];
  assign _02386_ = _03511_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10966" *) wt_pre_data[207:200] : wt4_sd_data[207:200];
  assign _02385_ = _03510_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10956" *) wt_pre_data[199:192] : wt4_sd_data[199:192];
  assign _02384_ = _03509_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10946" *) wt_pre_data[191:184] : wt4_sd_data[191:184];
  assign _02383_ = _03508_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10936" *) wt_pre_data[183:176] : wt4_sd_data[183:176];
  assign _02382_ = _03507_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10926" *) wt_pre_data[175:168] : wt4_sd_data[175:168];
  assign _02381_ = _03506_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10916" *) wt_pre_data[167:160] : wt4_sd_data[167:160];
  assign _02379_ = _03505_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10906" *) wt_pre_data[159:152] : wt4_sd_data[159:152];
  assign _02378_ = _03504_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10896" *) wt_pre_data[151:144] : wt4_sd_data[151:144];
  assign _02377_ = _03503_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10886" *) wt_pre_data[143:136] : wt4_sd_data[143:136];
  assign _02376_ = _03502_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10876" *) wt_pre_data[135:128] : wt4_sd_data[135:128];
  assign _02375_ = _03501_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10866" *) wt_pre_data[127:120] : wt4_sd_data[127:120];
  assign _02374_ = _03500_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10856" *) wt_pre_data[119:112] : wt4_sd_data[119:112];
  assign _02373_ = _03499_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10846" *) wt_pre_data[111:104] : wt4_sd_data[111:104];
  assign _02372_ = _03498_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10836" *) wt_pre_data[103:96] : wt4_sd_data[103:96];
  assign _02491_ = _03497_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10826" *) wt_pre_data[95:88] : wt4_sd_data[95:88];
  assign _02480_ = _03496_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10816" *) wt_pre_data[87:80] : wt4_sd_data[87:80];
  assign _02468_ = _03495_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10806" *) wt_pre_data[79:72] : wt4_sd_data[79:72];
  assign _02457_ = _03494_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10796" *) wt_pre_data[71:64] : wt4_sd_data[71:64];
  assign _02446_ = _03493_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10786" *) wt_pre_data[63:56] : wt4_sd_data[63:56];
  assign _02435_ = _03492_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10776" *) wt_pre_data[55:48] : wt4_sd_data[55:48];
  assign _02424_ = _03491_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10766" *) wt_pre_data[47:40] : wt4_sd_data[47:40];
  assign _02413_ = _03490_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10756" *) wt_pre_data[39:32] : wt4_sd_data[39:32];
  assign _02402_ = _03489_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10746" *) wt_pre_data[31:24] : wt4_sd_data[31:24];
  assign _02391_ = _03488_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10736" *) wt_pre_data[23:16] : wt4_sd_data[23:16];
  assign _02380_ = _03487_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10726" *) wt_pre_data[15:8] : wt4_sd_data[15:8];
  assign _02469_ = _03486_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10716" *) wt_pre_data[7:0] : wt4_sd_data[7:0];
  assign _02499_ = _03485_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10706" *) wt_pre_nan : wt4_sd_nan;
  assign _02497_ = _03485_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10696" *) wt_pre_exp : wt4_sd_exp;
  assign _02498_ = _03485_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10686" *) wt_pre_mask : wt4_sd_mask;
  assign _02500_ = wt_pre_sel[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10676" *) wt_pre_nz : wt4_sd_nz;
  assign _02109_ = _03484_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10650" *) wt_pre_data[1023:1016] : wt3_sd_data[1023:1016];
  assign _02108_ = _03483_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10640" *) wt_pre_data[1015:1008] : wt3_sd_data[1015:1008];
  assign _02107_ = _03482_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10630" *) wt_pre_data[1007:1000] : wt3_sd_data[1007:1000];
  assign _02234_ = _03481_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10620" *) wt_pre_data[999:992] : wt3_sd_data[999:992];
  assign _02233_ = _03480_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10610" *) wt_pre_data[991:984] : wt3_sd_data[991:984];
  assign _02232_ = _03479_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10600" *) wt_pre_data[983:976] : wt3_sd_data[983:976];
  assign _02231_ = _03478_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10590" *) wt_pre_data[975:968] : wt3_sd_data[975:968];
  assign _02230_ = _03477_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10580" *) wt_pre_data[967:960] : wt3_sd_data[967:960];
  assign _02228_ = _03476_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10570" *) wt_pre_data[959:952] : wt3_sd_data[959:952];
  assign _02227_ = _03475_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10560" *) wt_pre_data[951:944] : wt3_sd_data[951:944];
  assign _02226_ = _03474_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10550" *) wt_pre_data[943:936] : wt3_sd_data[943:936];
  assign _02225_ = _03473_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10540" *) wt_pre_data[935:928] : wt3_sd_data[935:928];
  assign _02224_ = _03472_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10530" *) wt_pre_data[927:920] : wt3_sd_data[927:920];
  assign _02223_ = _03471_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10520" *) wt_pre_data[919:912] : wt3_sd_data[919:912];
  assign _02222_ = _03470_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10510" *) wt_pre_data[911:904] : wt3_sd_data[911:904];
  assign _02221_ = _03469_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10500" *) wt_pre_data[903:896] : wt3_sd_data[903:896];
  assign _02220_ = _03468_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10490" *) wt_pre_data[895:888] : wt3_sd_data[895:888];
  assign _02219_ = _03467_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10480" *) wt_pre_data[887:880] : wt3_sd_data[887:880];
  assign _02217_ = _03466_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10470" *) wt_pre_data[879:872] : wt3_sd_data[879:872];
  assign _02216_ = _03465_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10460" *) wt_pre_data[871:864] : wt3_sd_data[871:864];
  assign _02215_ = _03464_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10450" *) wt_pre_data[863:856] : wt3_sd_data[863:856];
  assign _02214_ = _03463_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10440" *) wt_pre_data[855:848] : wt3_sd_data[855:848];
  assign _02213_ = _03462_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10430" *) wt_pre_data[847:840] : wt3_sd_data[847:840];
  assign _02212_ = _03461_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10420" *) wt_pre_data[839:832] : wt3_sd_data[839:832];
  assign _02211_ = _03460_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10410" *) wt_pre_data[831:824] : wt3_sd_data[831:824];
  assign _02210_ = _03459_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10400" *) wt_pre_data[823:816] : wt3_sd_data[823:816];
  assign _02209_ = _03458_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10390" *) wt_pre_data[815:808] : wt3_sd_data[815:808];
  assign _02208_ = _03457_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10380" *) wt_pre_data[807:800] : wt3_sd_data[807:800];
  assign _02205_ = _03456_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10370" *) wt_pre_data[799:792] : wt3_sd_data[799:792];
  assign _02204_ = _03455_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10360" *) wt_pre_data[791:784] : wt3_sd_data[791:784];
  assign _02203_ = _03454_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10350" *) wt_pre_data[783:776] : wt3_sd_data[783:776];
  assign _02202_ = _03453_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10340" *) wt_pre_data[775:768] : wt3_sd_data[775:768];
  assign _02201_ = _03452_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10330" *) wt_pre_data[767:760] : wt3_sd_data[767:760];
  assign _02200_ = _03451_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10320" *) wt_pre_data[759:752] : wt3_sd_data[759:752];
  assign _02199_ = _03450_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10310" *) wt_pre_data[751:744] : wt3_sd_data[751:744];
  assign _02198_ = _03449_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10300" *) wt_pre_data[743:736] : wt3_sd_data[743:736];
  assign _02197_ = _03448_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10290" *) wt_pre_data[735:728] : wt3_sd_data[735:728];
  assign _02196_ = _03447_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10280" *) wt_pre_data[727:720] : wt3_sd_data[727:720];
  assign _02194_ = _03446_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10270" *) wt_pre_data[719:712] : wt3_sd_data[719:712];
  assign _02193_ = _03445_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10260" *) wt_pre_data[711:704] : wt3_sd_data[711:704];
  assign _02192_ = _03444_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10250" *) wt_pre_data[703:696] : wt3_sd_data[703:696];
  assign _02191_ = _03443_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10240" *) wt_pre_data[695:688] : wt3_sd_data[695:688];
  assign _02190_ = _03442_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10230" *) wt_pre_data[687:680] : wt3_sd_data[687:680];
  assign _02189_ = _03441_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10220" *) wt_pre_data[679:672] : wt3_sd_data[679:672];
  assign _02188_ = _03440_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10210" *) wt_pre_data[671:664] : wt3_sd_data[671:664];
  assign _02187_ = _03439_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10200" *) wt_pre_data[663:656] : wt3_sd_data[663:656];
  assign _02186_ = _03438_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10190" *) wt_pre_data[655:648] : wt3_sd_data[655:648];
  assign _02185_ = _03437_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10180" *) wt_pre_data[647:640] : wt3_sd_data[647:640];
  assign _02183_ = _03436_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10170" *) wt_pre_data[639:632] : wt3_sd_data[639:632];
  assign _02182_ = _03435_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10160" *) wt_pre_data[631:624] : wt3_sd_data[631:624];
  assign _02181_ = _03434_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10150" *) wt_pre_data[623:616] : wt3_sd_data[623:616];
  assign _02180_ = _03433_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10140" *) wt_pre_data[615:608] : wt3_sd_data[615:608];
  assign _02179_ = _03432_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10130" *) wt_pre_data[607:600] : wt3_sd_data[607:600];
  assign _02178_ = _03431_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10120" *) wt_pre_data[599:592] : wt3_sd_data[599:592];
  assign _02177_ = _03430_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10110" *) wt_pre_data[591:584] : wt3_sd_data[591:584];
  assign _02176_ = _03429_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10100" *) wt_pre_data[583:576] : wt3_sd_data[583:576];
  assign _02175_ = _03428_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10090" *) wt_pre_data[575:568] : wt3_sd_data[575:568];
  assign _02174_ = _03427_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10080" *) wt_pre_data[567:560] : wt3_sd_data[567:560];
  assign _02172_ = _03426_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10070" *) wt_pre_data[559:552] : wt3_sd_data[559:552];
  assign _02171_ = _03425_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10060" *) wt_pre_data[551:544] : wt3_sd_data[551:544];
  assign _02170_ = _03424_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10050" *) wt_pre_data[543:536] : wt3_sd_data[543:536];
  assign _02169_ = _03423_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10040" *) wt_pre_data[535:528] : wt3_sd_data[535:528];
  assign _02168_ = _03422_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10030" *) wt_pre_data[527:520] : wt3_sd_data[527:520];
  assign _02167_ = _03421_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10020" *) wt_pre_data[519:512] : wt3_sd_data[519:512];
  assign _02166_ = _03420_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10010" *) wt_pre_data[511:504] : wt3_sd_data[511:504];
  assign _02165_ = _03419_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10000" *) wt_pre_data[503:496] : wt3_sd_data[503:496];
  assign _02164_ = _06278_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9990" *) wt_pre_data[495:488] : wt3_sd_data[495:488];
  assign _02163_ = _06277_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9980" *) wt_pre_data[487:480] : wt3_sd_data[487:480];
  assign _02161_ = _06276_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9970" *) wt_pre_data[479:472] : wt3_sd_data[479:472];
  assign _02160_ = _06275_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9960" *) wt_pre_data[471:464] : wt3_sd_data[471:464];
  assign _02159_ = _06274_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9950" *) wt_pre_data[463:456] : wt3_sd_data[463:456];
  assign _02158_ = _06273_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9940" *) wt_pre_data[455:448] : wt3_sd_data[455:448];
  assign _02157_ = _06272_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9930" *) wt_pre_data[447:440] : wt3_sd_data[447:440];
  assign _02156_ = _06271_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9920" *) wt_pre_data[439:432] : wt3_sd_data[439:432];
  assign _02155_ = _06270_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9910" *) wt_pre_data[431:424] : wt3_sd_data[431:424];
  assign _02154_ = _06269_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9900" *) wt_pre_data[423:416] : wt3_sd_data[423:416];
  assign _02153_ = _06268_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9890" *) wt_pre_data[415:408] : wt3_sd_data[415:408];
  assign _02152_ = _06267_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9880" *) wt_pre_data[407:400] : wt3_sd_data[407:400];
  assign _02150_ = _06266_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9870" *) wt_pre_data[399:392] : wt3_sd_data[399:392];
  assign _02149_ = _06265_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9860" *) wt_pre_data[391:384] : wt3_sd_data[391:384];
  assign _02148_ = _06264_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9850" *) wt_pre_data[383:376] : wt3_sd_data[383:376];
  assign _02147_ = _06263_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9840" *) wt_pre_data[375:368] : wt3_sd_data[375:368];
  assign _02146_ = _06262_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9830" *) wt_pre_data[367:360] : wt3_sd_data[367:360];
  assign _02145_ = _06261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9820" *) wt_pre_data[359:352] : wt3_sd_data[359:352];
  assign _02144_ = _06260_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9810" *) wt_pre_data[351:344] : wt3_sd_data[351:344];
  assign _02143_ = _06259_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9800" *) wt_pre_data[343:336] : wt3_sd_data[343:336];
  assign _02142_ = _06258_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9790" *) wt_pre_data[335:328] : wt3_sd_data[335:328];
  assign _02141_ = _06257_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9780" *) wt_pre_data[327:320] : wt3_sd_data[327:320];
  assign _02139_ = _06256_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9770" *) wt_pre_data[319:312] : wt3_sd_data[319:312];
  assign _02138_ = _06255_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9760" *) wt_pre_data[311:304] : wt3_sd_data[311:304];
  assign _02137_ = _06254_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9750" *) wt_pre_data[303:296] : wt3_sd_data[303:296];
  assign _02136_ = _06253_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9740" *) wt_pre_data[295:288] : wt3_sd_data[295:288];
  assign _02135_ = _06252_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9730" *) wt_pre_data[287:280] : wt3_sd_data[287:280];
  assign _02134_ = _06251_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9720" *) wt_pre_data[279:272] : wt3_sd_data[279:272];
  assign _02133_ = _06250_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9710" *) wt_pre_data[271:264] : wt3_sd_data[271:264];
  assign _02132_ = _06249_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9700" *) wt_pre_data[263:256] : wt3_sd_data[263:256];
  assign _02131_ = _06248_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9690" *) wt_pre_data[255:248] : wt3_sd_data[255:248];
  assign _02130_ = _06247_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9680" *) wt_pre_data[247:240] : wt3_sd_data[247:240];
  assign _02128_ = _06246_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9670" *) wt_pre_data[239:232] : wt3_sd_data[239:232];
  assign _02127_ = _06245_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9660" *) wt_pre_data[231:224] : wt3_sd_data[231:224];
  assign _02126_ = _06244_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9650" *) wt_pre_data[223:216] : wt3_sd_data[223:216];
  assign _02125_ = _06243_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9640" *) wt_pre_data[215:208] : wt3_sd_data[215:208];
  assign _02124_ = _06242_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9630" *) wt_pre_data[207:200] : wt3_sd_data[207:200];
  assign _02123_ = _06241_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9620" *) wt_pre_data[199:192] : wt3_sd_data[199:192];
  assign _02122_ = _06240_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9610" *) wt_pre_data[191:184] : wt3_sd_data[191:184];
  assign _02121_ = _06239_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9600" *) wt_pre_data[183:176] : wt3_sd_data[183:176];
  assign _02120_ = _06238_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9590" *) wt_pre_data[175:168] : wt3_sd_data[175:168];
  assign _02119_ = _06237_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9580" *) wt_pre_data[167:160] : wt3_sd_data[167:160];
  assign _02117_ = _06236_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9570" *) wt_pre_data[159:152] : wt3_sd_data[159:152];
  assign _02116_ = _06235_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9560" *) wt_pre_data[151:144] : wt3_sd_data[151:144];
  assign _02115_ = _06234_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9550" *) wt_pre_data[143:136] : wt3_sd_data[143:136];
  assign _02114_ = _06233_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9540" *) wt_pre_data[135:128] : wt3_sd_data[135:128];
  assign _02113_ = _06232_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9530" *) wt_pre_data[127:120] : wt3_sd_data[127:120];
  assign _02112_ = _06231_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9520" *) wt_pre_data[119:112] : wt3_sd_data[119:112];
  assign _02111_ = _06230_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9510" *) wt_pre_data[111:104] : wt3_sd_data[111:104];
  assign _02110_ = _06229_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9500" *) wt_pre_data[103:96] : wt3_sd_data[103:96];
  assign _02229_ = _06228_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9490" *) wt_pre_data[95:88] : wt3_sd_data[95:88];
  assign _02218_ = _06227_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9480" *) wt_pre_data[87:80] : wt3_sd_data[87:80];
  assign _02206_ = _06226_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9470" *) wt_pre_data[79:72] : wt3_sd_data[79:72];
  assign _02195_ = _06225_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9460" *) wt_pre_data[71:64] : wt3_sd_data[71:64];
  assign _02184_ = _06224_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9450" *) wt_pre_data[63:56] : wt3_sd_data[63:56];
  assign _02173_ = _06223_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9440" *) wt_pre_data[55:48] : wt3_sd_data[55:48];
  assign _02162_ = _06222_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9430" *) wt_pre_data[47:40] : wt3_sd_data[47:40];
  assign _02151_ = _06221_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9420" *) wt_pre_data[39:32] : wt3_sd_data[39:32];
  assign _02140_ = _06220_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9410" *) wt_pre_data[31:24] : wt3_sd_data[31:24];
  assign _02129_ = _06219_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9400" *) wt_pre_data[23:16] : wt3_sd_data[23:16];
  assign _02118_ = _06218_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9390" *) wt_pre_data[15:8] : wt3_sd_data[15:8];
  assign _02207_ = _06217_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9380" *) wt_pre_data[7:0] : wt3_sd_data[7:0];
  assign _02237_ = _06216_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9370" *) wt_pre_nan : wt3_sd_nan;
  assign _02235_ = _06216_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9360" *) wt_pre_exp : wt3_sd_exp;
  assign _02236_ = _06216_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9350" *) wt_pre_mask : wt3_sd_mask;
  assign _02238_ = wt_pre_sel[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9340" *) wt_pre_nz : wt3_sd_nz;
  assign _01847_ = _06215_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9314" *) wt_pre_data[1023:1016] : wt2_sd_data[1023:1016];
  assign _01846_ = _06214_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9304" *) wt_pre_data[1015:1008] : wt2_sd_data[1015:1008];
  assign _01845_ = _06213_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9294" *) wt_pre_data[1007:1000] : wt2_sd_data[1007:1000];
  assign _01972_ = _06212_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9284" *) wt_pre_data[999:992] : wt2_sd_data[999:992];
  assign _01971_ = _06211_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9274" *) wt_pre_data[991:984] : wt2_sd_data[991:984];
  assign _01970_ = _06210_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9264" *) wt_pre_data[983:976] : wt2_sd_data[983:976];
  assign _01969_ = _06209_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9254" *) wt_pre_data[975:968] : wt2_sd_data[975:968];
  assign _01968_ = _06208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9244" *) wt_pre_data[967:960] : wt2_sd_data[967:960];
  assign _01966_ = _06207_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9234" *) wt_pre_data[959:952] : wt2_sd_data[959:952];
  assign _01965_ = _06206_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9224" *) wt_pre_data[951:944] : wt2_sd_data[951:944];
  assign _01964_ = _06205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9214" *) wt_pre_data[943:936] : wt2_sd_data[943:936];
  assign _01963_ = _06204_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9204" *) wt_pre_data[935:928] : wt2_sd_data[935:928];
  assign _01962_ = _06203_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9194" *) wt_pre_data[927:920] : wt2_sd_data[927:920];
  assign _01961_ = _06202_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9184" *) wt_pre_data[919:912] : wt2_sd_data[919:912];
  assign _01960_ = _06201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9174" *) wt_pre_data[911:904] : wt2_sd_data[911:904];
  assign _01959_ = _06200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9164" *) wt_pre_data[903:896] : wt2_sd_data[903:896];
  assign _01958_ = _06199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9154" *) wt_pre_data[895:888] : wt2_sd_data[895:888];
  assign _01957_ = _06198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9144" *) wt_pre_data[887:880] : wt2_sd_data[887:880];
  assign _01955_ = _06197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9134" *) wt_pre_data[879:872] : wt2_sd_data[879:872];
  assign _01954_ = _06196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9124" *) wt_pre_data[871:864] : wt2_sd_data[871:864];
  assign _01953_ = _06195_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9114" *) wt_pre_data[863:856] : wt2_sd_data[863:856];
  assign _01952_ = _06194_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9104" *) wt_pre_data[855:848] : wt2_sd_data[855:848];
  assign _01951_ = _06193_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9094" *) wt_pre_data[847:840] : wt2_sd_data[847:840];
  assign _01950_ = _06192_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9084" *) wt_pre_data[839:832] : wt2_sd_data[839:832];
  assign _01949_ = _06191_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9074" *) wt_pre_data[831:824] : wt2_sd_data[831:824];
  assign _01948_ = _06190_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9064" *) wt_pre_data[823:816] : wt2_sd_data[823:816];
  assign _01947_ = _06189_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9054" *) wt_pre_data[815:808] : wt2_sd_data[815:808];
  assign _01946_ = _06188_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9044" *) wt_pre_data[807:800] : wt2_sd_data[807:800];
  assign _01943_ = _06187_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9034" *) wt_pre_data[799:792] : wt2_sd_data[799:792];
  assign _01942_ = _06186_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9024" *) wt_pre_data[791:784] : wt2_sd_data[791:784];
  assign _01941_ = _06185_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9014" *) wt_pre_data[783:776] : wt2_sd_data[783:776];
  assign _01940_ = _06184_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9004" *) wt_pre_data[775:768] : wt2_sd_data[775:768];
  assign _01939_ = _06183_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8994" *) wt_pre_data[767:760] : wt2_sd_data[767:760];
  assign _01938_ = _06182_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8984" *) wt_pre_data[759:752] : wt2_sd_data[759:752];
  assign _01937_ = _06181_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8974" *) wt_pre_data[751:744] : wt2_sd_data[751:744];
  assign _01936_ = _06180_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8964" *) wt_pre_data[743:736] : wt2_sd_data[743:736];
  assign _01935_ = _06179_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8954" *) wt_pre_data[735:728] : wt2_sd_data[735:728];
  assign _01934_ = _06178_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8944" *) wt_pre_data[727:720] : wt2_sd_data[727:720];
  assign _01932_ = _06177_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8934" *) wt_pre_data[719:712] : wt2_sd_data[719:712];
  assign _01931_ = _06176_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8924" *) wt_pre_data[711:704] : wt2_sd_data[711:704];
  assign _01930_ = _06175_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8914" *) wt_pre_data[703:696] : wt2_sd_data[703:696];
  assign _01929_ = _06174_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8904" *) wt_pre_data[695:688] : wt2_sd_data[695:688];
  assign _01928_ = _06173_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8894" *) wt_pre_data[687:680] : wt2_sd_data[687:680];
  assign _01927_ = _06172_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8884" *) wt_pre_data[679:672] : wt2_sd_data[679:672];
  assign _01926_ = _06171_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8874" *) wt_pre_data[671:664] : wt2_sd_data[671:664];
  assign _01925_ = _06170_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8864" *) wt_pre_data[663:656] : wt2_sd_data[663:656];
  assign _01924_ = _06169_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8854" *) wt_pre_data[655:648] : wt2_sd_data[655:648];
  assign _01923_ = _06168_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8844" *) wt_pre_data[647:640] : wt2_sd_data[647:640];
  assign _01921_ = _06167_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8834" *) wt_pre_data[639:632] : wt2_sd_data[639:632];
  assign _01920_ = _06166_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8824" *) wt_pre_data[631:624] : wt2_sd_data[631:624];
  assign _01919_ = _06165_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8814" *) wt_pre_data[623:616] : wt2_sd_data[623:616];
  assign _01918_ = _06164_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8804" *) wt_pre_data[615:608] : wt2_sd_data[615:608];
  assign _01917_ = _06163_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8794" *) wt_pre_data[607:600] : wt2_sd_data[607:600];
  assign _01916_ = _06162_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8784" *) wt_pre_data[599:592] : wt2_sd_data[599:592];
  assign _01915_ = _06161_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8774" *) wt_pre_data[591:584] : wt2_sd_data[591:584];
  assign _01914_ = _06160_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8764" *) wt_pre_data[583:576] : wt2_sd_data[583:576];
  assign _01913_ = _06159_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8754" *) wt_pre_data[575:568] : wt2_sd_data[575:568];
  assign _01912_ = _06158_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8744" *) wt_pre_data[567:560] : wt2_sd_data[567:560];
  assign _01910_ = _06157_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8734" *) wt_pre_data[559:552] : wt2_sd_data[559:552];
  assign _01909_ = _06156_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8724" *) wt_pre_data[551:544] : wt2_sd_data[551:544];
  assign _01908_ = _06155_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8714" *) wt_pre_data[543:536] : wt2_sd_data[543:536];
  assign _01907_ = _06154_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8704" *) wt_pre_data[535:528] : wt2_sd_data[535:528];
  assign _01906_ = _06153_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8694" *) wt_pre_data[527:520] : wt2_sd_data[527:520];
  assign _01905_ = _06152_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8684" *) wt_pre_data[519:512] : wt2_sd_data[519:512];
  assign _01904_ = _06151_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8674" *) wt_pre_data[511:504] : wt2_sd_data[511:504];
  assign _01903_ = _06150_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8664" *) wt_pre_data[503:496] : wt2_sd_data[503:496];
  assign _01902_ = _06149_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8654" *) wt_pre_data[495:488] : wt2_sd_data[495:488];
  assign _01901_ = _06148_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8644" *) wt_pre_data[487:480] : wt2_sd_data[487:480];
  assign _01899_ = _06147_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8634" *) wt_pre_data[479:472] : wt2_sd_data[479:472];
  assign _01898_ = _06146_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8624" *) wt_pre_data[471:464] : wt2_sd_data[471:464];
  assign _01897_ = _06145_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8614" *) wt_pre_data[463:456] : wt2_sd_data[463:456];
  assign _01896_ = _06144_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8604" *) wt_pre_data[455:448] : wt2_sd_data[455:448];
  assign _01895_ = _06143_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8594" *) wt_pre_data[447:440] : wt2_sd_data[447:440];
  assign _01894_ = _06142_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8584" *) wt_pre_data[439:432] : wt2_sd_data[439:432];
  assign _01893_ = _06141_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8574" *) wt_pre_data[431:424] : wt2_sd_data[431:424];
  assign _01892_ = _06140_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8564" *) wt_pre_data[423:416] : wt2_sd_data[423:416];
  assign _01891_ = _06139_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8554" *) wt_pre_data[415:408] : wt2_sd_data[415:408];
  assign _01890_ = _06138_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8544" *) wt_pre_data[407:400] : wt2_sd_data[407:400];
  assign _01888_ = _06137_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8534" *) wt_pre_data[399:392] : wt2_sd_data[399:392];
  assign _01887_ = _06136_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8524" *) wt_pre_data[391:384] : wt2_sd_data[391:384];
  assign _01886_ = _06135_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8514" *) wt_pre_data[383:376] : wt2_sd_data[383:376];
  assign _01885_ = _06134_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8504" *) wt_pre_data[375:368] : wt2_sd_data[375:368];
  assign _01884_ = _06133_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8494" *) wt_pre_data[367:360] : wt2_sd_data[367:360];
  assign _01883_ = _06132_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8484" *) wt_pre_data[359:352] : wt2_sd_data[359:352];
  assign _01882_ = _06131_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8474" *) wt_pre_data[351:344] : wt2_sd_data[351:344];
  assign _01881_ = _06130_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8464" *) wt_pre_data[343:336] : wt2_sd_data[343:336];
  assign _01880_ = _06129_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8454" *) wt_pre_data[335:328] : wt2_sd_data[335:328];
  assign _01879_ = _06128_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8444" *) wt_pre_data[327:320] : wt2_sd_data[327:320];
  assign _01877_ = _06127_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8434" *) wt_pre_data[319:312] : wt2_sd_data[319:312];
  assign _01876_ = _06126_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8424" *) wt_pre_data[311:304] : wt2_sd_data[311:304];
  assign _01875_ = _06125_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8414" *) wt_pre_data[303:296] : wt2_sd_data[303:296];
  assign _01874_ = _06124_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8404" *) wt_pre_data[295:288] : wt2_sd_data[295:288];
  assign _01873_ = _06123_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8394" *) wt_pre_data[287:280] : wt2_sd_data[287:280];
  assign _01872_ = _06122_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8384" *) wt_pre_data[279:272] : wt2_sd_data[279:272];
  assign _01871_ = _06121_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8374" *) wt_pre_data[271:264] : wt2_sd_data[271:264];
  assign _01870_ = _06120_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8364" *) wt_pre_data[263:256] : wt2_sd_data[263:256];
  assign _01869_ = _06119_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8354" *) wt_pre_data[255:248] : wt2_sd_data[255:248];
  assign _01868_ = _06118_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8344" *) wt_pre_data[247:240] : wt2_sd_data[247:240];
  assign _01866_ = _06117_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8334" *) wt_pre_data[239:232] : wt2_sd_data[239:232];
  assign _01865_ = _06116_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8324" *) wt_pre_data[231:224] : wt2_sd_data[231:224];
  assign _01864_ = _06115_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8314" *) wt_pre_data[223:216] : wt2_sd_data[223:216];
  assign _01863_ = _06114_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8304" *) wt_pre_data[215:208] : wt2_sd_data[215:208];
  assign _01862_ = _06113_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8294" *) wt_pre_data[207:200] : wt2_sd_data[207:200];
  assign _01861_ = _06112_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8284" *) wt_pre_data[199:192] : wt2_sd_data[199:192];
  assign _01860_ = _06111_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8274" *) wt_pre_data[191:184] : wt2_sd_data[191:184];
  assign _01859_ = _06110_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8264" *) wt_pre_data[183:176] : wt2_sd_data[183:176];
  assign _01858_ = _06109_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8254" *) wt_pre_data[175:168] : wt2_sd_data[175:168];
  assign _01857_ = _06108_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8244" *) wt_pre_data[167:160] : wt2_sd_data[167:160];
  assign _01855_ = _06107_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8234" *) wt_pre_data[159:152] : wt2_sd_data[159:152];
  assign _01854_ = _06106_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8224" *) wt_pre_data[151:144] : wt2_sd_data[151:144];
  assign _01853_ = _06105_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8214" *) wt_pre_data[143:136] : wt2_sd_data[143:136];
  assign _01852_ = _06104_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8204" *) wt_pre_data[135:128] : wt2_sd_data[135:128];
  assign _01851_ = _06103_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8194" *) wt_pre_data[127:120] : wt2_sd_data[127:120];
  assign _01850_ = _06102_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8184" *) wt_pre_data[119:112] : wt2_sd_data[119:112];
  assign _01849_ = _06101_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8174" *) wt_pre_data[111:104] : wt2_sd_data[111:104];
  assign _01848_ = _06100_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8164" *) wt_pre_data[103:96] : wt2_sd_data[103:96];
  assign _01967_ = _06099_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8154" *) wt_pre_data[95:88] : wt2_sd_data[95:88];
  assign _01956_ = _06098_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8144" *) wt_pre_data[87:80] : wt2_sd_data[87:80];
  assign _01944_ = _06097_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8134" *) wt_pre_data[79:72] : wt2_sd_data[79:72];
  assign _01933_ = _06096_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8124" *) wt_pre_data[71:64] : wt2_sd_data[71:64];
  assign _01922_ = _06095_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8114" *) wt_pre_data[63:56] : wt2_sd_data[63:56];
  assign _01911_ = _06094_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8104" *) wt_pre_data[55:48] : wt2_sd_data[55:48];
  assign _01900_ = _06093_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8094" *) wt_pre_data[47:40] : wt2_sd_data[47:40];
  assign _01889_ = _06092_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8084" *) wt_pre_data[39:32] : wt2_sd_data[39:32];
  assign _01878_ = _06091_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8074" *) wt_pre_data[31:24] : wt2_sd_data[31:24];
  assign _01867_ = _06090_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8064" *) wt_pre_data[23:16] : wt2_sd_data[23:16];
  assign _01856_ = _06089_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8054" *) wt_pre_data[15:8] : wt2_sd_data[15:8];
  assign _01945_ = _06088_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8044" *) wt_pre_data[7:0] : wt2_sd_data[7:0];
  assign _01975_ = _06087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8034" *) wt_pre_nan : wt2_sd_nan;
  assign _01973_ = _06087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8024" *) wt_pre_exp : wt2_sd_exp;
  assign _01974_ = _06087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8014" *) wt_pre_mask : wt2_sd_mask;
  assign _01976_ = wt_pre_sel[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:8004" *) wt_pre_nz : wt2_sd_nz;
  assign _01585_ = _06086_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7978" *) wt_pre_data[1023:1016] : wt1_sd_data[1023:1016];
  assign _01584_ = _06085_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7968" *) wt_pre_data[1015:1008] : wt1_sd_data[1015:1008];
  assign _01583_ = _06084_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7958" *) wt_pre_data[1007:1000] : wt1_sd_data[1007:1000];
  assign _01710_ = _06083_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7948" *) wt_pre_data[999:992] : wt1_sd_data[999:992];
  assign _01709_ = _06082_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7938" *) wt_pre_data[991:984] : wt1_sd_data[991:984];
  assign _01708_ = _06081_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7928" *) wt_pre_data[983:976] : wt1_sd_data[983:976];
  assign _01707_ = _06080_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7918" *) wt_pre_data[975:968] : wt1_sd_data[975:968];
  assign _01706_ = _06079_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7908" *) wt_pre_data[967:960] : wt1_sd_data[967:960];
  assign _01704_ = _06078_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7898" *) wt_pre_data[959:952] : wt1_sd_data[959:952];
  assign _01703_ = _06077_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7888" *) wt_pre_data[951:944] : wt1_sd_data[951:944];
  assign _01702_ = _06076_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7878" *) wt_pre_data[943:936] : wt1_sd_data[943:936];
  assign _01701_ = _06075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7868" *) wt_pre_data[935:928] : wt1_sd_data[935:928];
  assign _01700_ = _06074_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7858" *) wt_pre_data[927:920] : wt1_sd_data[927:920];
  assign _01699_ = _06073_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7848" *) wt_pre_data[919:912] : wt1_sd_data[919:912];
  assign _01698_ = _06072_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7838" *) wt_pre_data[911:904] : wt1_sd_data[911:904];
  assign _01697_ = _06071_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7828" *) wt_pre_data[903:896] : wt1_sd_data[903:896];
  assign _01696_ = _06070_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7818" *) wt_pre_data[895:888] : wt1_sd_data[895:888];
  assign _01695_ = _06069_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7808" *) wt_pre_data[887:880] : wt1_sd_data[887:880];
  assign _01693_ = _06068_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7798" *) wt_pre_data[879:872] : wt1_sd_data[879:872];
  assign _01692_ = _06067_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7788" *) wt_pre_data[871:864] : wt1_sd_data[871:864];
  assign _01691_ = _06066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7778" *) wt_pre_data[863:856] : wt1_sd_data[863:856];
  assign _01690_ = _06065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7768" *) wt_pre_data[855:848] : wt1_sd_data[855:848];
  assign _01689_ = _06064_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7758" *) wt_pre_data[847:840] : wt1_sd_data[847:840];
  assign _01688_ = _06063_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7748" *) wt_pre_data[839:832] : wt1_sd_data[839:832];
  assign _01687_ = _06062_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7738" *) wt_pre_data[831:824] : wt1_sd_data[831:824];
  assign _01686_ = _06061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7728" *) wt_pre_data[823:816] : wt1_sd_data[823:816];
  assign _01685_ = _06060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7718" *) wt_pre_data[815:808] : wt1_sd_data[815:808];
  assign _01684_ = _06059_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7708" *) wt_pre_data[807:800] : wt1_sd_data[807:800];
  assign _01681_ = _06058_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7698" *) wt_pre_data[799:792] : wt1_sd_data[799:792];
  assign _01680_ = _06057_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7688" *) wt_pre_data[791:784] : wt1_sd_data[791:784];
  assign _01679_ = _06056_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7678" *) wt_pre_data[783:776] : wt1_sd_data[783:776];
  assign _01678_ = _06055_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7668" *) wt_pre_data[775:768] : wt1_sd_data[775:768];
  assign _01677_ = _06054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7658" *) wt_pre_data[767:760] : wt1_sd_data[767:760];
  assign _01676_ = _06053_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7648" *) wt_pre_data[759:752] : wt1_sd_data[759:752];
  assign _01675_ = _06052_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7638" *) wt_pre_data[751:744] : wt1_sd_data[751:744];
  assign _01674_ = _06051_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7628" *) wt_pre_data[743:736] : wt1_sd_data[743:736];
  assign _01673_ = _06050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7618" *) wt_pre_data[735:728] : wt1_sd_data[735:728];
  assign _01672_ = _06049_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7608" *) wt_pre_data[727:720] : wt1_sd_data[727:720];
  assign _01670_ = _06048_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7598" *) wt_pre_data[719:712] : wt1_sd_data[719:712];
  assign _01669_ = _06047_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7588" *) wt_pre_data[711:704] : wt1_sd_data[711:704];
  assign _01668_ = _06046_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7578" *) wt_pre_data[703:696] : wt1_sd_data[703:696];
  assign _01667_ = _06045_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7568" *) wt_pre_data[695:688] : wt1_sd_data[695:688];
  assign _01666_ = _06044_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7558" *) wt_pre_data[687:680] : wt1_sd_data[687:680];
  assign _01665_ = _06043_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7548" *) wt_pre_data[679:672] : wt1_sd_data[679:672];
  assign _01664_ = _06042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7538" *) wt_pre_data[671:664] : wt1_sd_data[671:664];
  assign _01663_ = _06041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7528" *) wt_pre_data[663:656] : wt1_sd_data[663:656];
  assign _01662_ = _06040_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7518" *) wt_pre_data[655:648] : wt1_sd_data[655:648];
  assign _01661_ = _06039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7508" *) wt_pre_data[647:640] : wt1_sd_data[647:640];
  assign _01659_ = _06038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7498" *) wt_pre_data[639:632] : wt1_sd_data[639:632];
  assign _01658_ = _06037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7488" *) wt_pre_data[631:624] : wt1_sd_data[631:624];
  assign _01657_ = _06036_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7478" *) wt_pre_data[623:616] : wt1_sd_data[623:616];
  assign _01656_ = _06035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7468" *) wt_pre_data[615:608] : wt1_sd_data[615:608];
  assign _01655_ = _06034_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7458" *) wt_pre_data[607:600] : wt1_sd_data[607:600];
  assign _01654_ = _06033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7448" *) wt_pre_data[599:592] : wt1_sd_data[599:592];
  assign _01653_ = _06032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7438" *) wt_pre_data[591:584] : wt1_sd_data[591:584];
  assign _01652_ = _06031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7428" *) wt_pre_data[583:576] : wt1_sd_data[583:576];
  assign _01651_ = _06030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7418" *) wt_pre_data[575:568] : wt1_sd_data[575:568];
  assign _01650_ = _06029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7408" *) wt_pre_data[567:560] : wt1_sd_data[567:560];
  assign _01648_ = _06028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7398" *) wt_pre_data[559:552] : wt1_sd_data[559:552];
  assign _01647_ = _06027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7388" *) wt_pre_data[551:544] : wt1_sd_data[551:544];
  assign _01646_ = _06026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7378" *) wt_pre_data[543:536] : wt1_sd_data[543:536];
  assign _01645_ = _06025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7368" *) wt_pre_data[535:528] : wt1_sd_data[535:528];
  assign _01644_ = _06024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7358" *) wt_pre_data[527:520] : wt1_sd_data[527:520];
  assign _01643_ = _06023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7348" *) wt_pre_data[519:512] : wt1_sd_data[519:512];
  assign _01642_ = _06022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7338" *) wt_pre_data[511:504] : wt1_sd_data[511:504];
  assign _01641_ = _06021_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7328" *) wt_pre_data[503:496] : wt1_sd_data[503:496];
  assign _01640_ = _06020_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7318" *) wt_pre_data[495:488] : wt1_sd_data[495:488];
  assign _01639_ = _06019_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7308" *) wt_pre_data[487:480] : wt1_sd_data[487:480];
  assign _01637_ = _06018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7298" *) wt_pre_data[479:472] : wt1_sd_data[479:472];
  assign _01636_ = _06017_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7288" *) wt_pre_data[471:464] : wt1_sd_data[471:464];
  assign _01635_ = _06016_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7278" *) wt_pre_data[463:456] : wt1_sd_data[463:456];
  assign _01634_ = _06015_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7268" *) wt_pre_data[455:448] : wt1_sd_data[455:448];
  assign _01633_ = _06014_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7258" *) wt_pre_data[447:440] : wt1_sd_data[447:440];
  assign _01632_ = _06013_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7248" *) wt_pre_data[439:432] : wt1_sd_data[439:432];
  assign _01631_ = _06012_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7238" *) wt_pre_data[431:424] : wt1_sd_data[431:424];
  assign _01630_ = _06011_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7228" *) wt_pre_data[423:416] : wt1_sd_data[423:416];
  assign _01629_ = _06010_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7218" *) wt_pre_data[415:408] : wt1_sd_data[415:408];
  assign _01628_ = _06009_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7208" *) wt_pre_data[407:400] : wt1_sd_data[407:400];
  assign _01626_ = _06008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7198" *) wt_pre_data[399:392] : wt1_sd_data[399:392];
  assign _01625_ = _06007_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7188" *) wt_pre_data[391:384] : wt1_sd_data[391:384];
  assign _01624_ = _06006_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7178" *) wt_pre_data[383:376] : wt1_sd_data[383:376];
  assign _01623_ = _06005_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7168" *) wt_pre_data[375:368] : wt1_sd_data[375:368];
  assign _01622_ = _06004_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7158" *) wt_pre_data[367:360] : wt1_sd_data[367:360];
  assign _01621_ = _06003_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7148" *) wt_pre_data[359:352] : wt1_sd_data[359:352];
  assign _01620_ = _06002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7138" *) wt_pre_data[351:344] : wt1_sd_data[351:344];
  assign _01619_ = _06001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7128" *) wt_pre_data[343:336] : wt1_sd_data[343:336];
  assign _01618_ = _06000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7118" *) wt_pre_data[335:328] : wt1_sd_data[335:328];
  assign _01617_ = _05999_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7108" *) wt_pre_data[327:320] : wt1_sd_data[327:320];
  assign _01615_ = _05998_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7098" *) wt_pre_data[319:312] : wt1_sd_data[319:312];
  assign _01614_ = _05997_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7088" *) wt_pre_data[311:304] : wt1_sd_data[311:304];
  assign _01613_ = _05996_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7078" *) wt_pre_data[303:296] : wt1_sd_data[303:296];
  assign _01612_ = _05995_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7068" *) wt_pre_data[295:288] : wt1_sd_data[295:288];
  assign _01611_ = _05994_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7058" *) wt_pre_data[287:280] : wt1_sd_data[287:280];
  assign _01610_ = _05993_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7048" *) wt_pre_data[279:272] : wt1_sd_data[279:272];
  assign _01609_ = _05992_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7038" *) wt_pre_data[271:264] : wt1_sd_data[271:264];
  assign _01608_ = _05991_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7028" *) wt_pre_data[263:256] : wt1_sd_data[263:256];
  assign _01607_ = _05990_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7018" *) wt_pre_data[255:248] : wt1_sd_data[255:248];
  assign _01606_ = _05989_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7008" *) wt_pre_data[247:240] : wt1_sd_data[247:240];
  assign _01604_ = _05988_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6998" *) wt_pre_data[239:232] : wt1_sd_data[239:232];
  assign _01603_ = _05987_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6988" *) wt_pre_data[231:224] : wt1_sd_data[231:224];
  assign _01602_ = _05986_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6978" *) wt_pre_data[223:216] : wt1_sd_data[223:216];
  assign _01601_ = _05985_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6968" *) wt_pre_data[215:208] : wt1_sd_data[215:208];
  assign _01600_ = _05984_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6958" *) wt_pre_data[207:200] : wt1_sd_data[207:200];
  assign _01599_ = _05983_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6948" *) wt_pre_data[199:192] : wt1_sd_data[199:192];
  assign _01598_ = _05982_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6938" *) wt_pre_data[191:184] : wt1_sd_data[191:184];
  assign _01597_ = _05981_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6928" *) wt_pre_data[183:176] : wt1_sd_data[183:176];
  assign _01596_ = _05980_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6918" *) wt_pre_data[175:168] : wt1_sd_data[175:168];
  assign _01595_ = _05979_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6908" *) wt_pre_data[167:160] : wt1_sd_data[167:160];
  assign _01593_ = _05978_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6898" *) wt_pre_data[159:152] : wt1_sd_data[159:152];
  assign _01592_ = _05977_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6888" *) wt_pre_data[151:144] : wt1_sd_data[151:144];
  assign _01591_ = _05976_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6878" *) wt_pre_data[143:136] : wt1_sd_data[143:136];
  assign _01590_ = _05975_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6868" *) wt_pre_data[135:128] : wt1_sd_data[135:128];
  assign _01589_ = _05974_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6858" *) wt_pre_data[127:120] : wt1_sd_data[127:120];
  assign _01588_ = _05973_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6848" *) wt_pre_data[119:112] : wt1_sd_data[119:112];
  assign _01587_ = _05972_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6838" *) wt_pre_data[111:104] : wt1_sd_data[111:104];
  assign _01586_ = _05971_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6828" *) wt_pre_data[103:96] : wt1_sd_data[103:96];
  assign _01705_ = _05970_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6818" *) wt_pre_data[95:88] : wt1_sd_data[95:88];
  assign _01694_ = _05969_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6808" *) wt_pre_data[87:80] : wt1_sd_data[87:80];
  assign _01682_ = _05968_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6798" *) wt_pre_data[79:72] : wt1_sd_data[79:72];
  assign _01671_ = _05967_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6788" *) wt_pre_data[71:64] : wt1_sd_data[71:64];
  assign _01660_ = _05966_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6778" *) wt_pre_data[63:56] : wt1_sd_data[63:56];
  assign _01649_ = _05965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6768" *) wt_pre_data[55:48] : wt1_sd_data[55:48];
  assign _01638_ = _05964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6758" *) wt_pre_data[47:40] : wt1_sd_data[47:40];
  assign _01627_ = _05963_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6748" *) wt_pre_data[39:32] : wt1_sd_data[39:32];
  assign _01616_ = _05962_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6738" *) wt_pre_data[31:24] : wt1_sd_data[31:24];
  assign _01605_ = _05961_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6728" *) wt_pre_data[23:16] : wt1_sd_data[23:16];
  assign _01594_ = _05960_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6718" *) wt_pre_data[15:8] : wt1_sd_data[15:8];
  assign _01683_ = _05959_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6708" *) wt_pre_data[7:0] : wt1_sd_data[7:0];
  assign _01713_ = _05958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6698" *) wt_pre_nan : wt1_sd_nan;
  assign _01711_ = _05958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6688" *) wt_pre_exp : wt1_sd_exp;
  assign _01712_ = _05958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6678" *) wt_pre_mask : wt1_sd_mask;
  assign _01714_ = wt_pre_sel[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6668" *) wt_pre_nz : wt1_sd_nz;
  assign _01323_ = _05957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6642" *) wt_pre_data[1023:1016] : wt0_sd_data[1023:1016];
  assign _01322_ = _05956_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6632" *) wt_pre_data[1015:1008] : wt0_sd_data[1015:1008];
  assign _01321_ = _05955_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6622" *) wt_pre_data[1007:1000] : wt0_sd_data[1007:1000];
  assign _01448_ = _05954_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6612" *) wt_pre_data[999:992] : wt0_sd_data[999:992];
  assign _01447_ = _05953_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6602" *) wt_pre_data[991:984] : wt0_sd_data[991:984];
  assign _01446_ = _05952_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6592" *) wt_pre_data[983:976] : wt0_sd_data[983:976];
  assign _01445_ = _05951_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6582" *) wt_pre_data[975:968] : wt0_sd_data[975:968];
  assign _01444_ = _05950_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6572" *) wt_pre_data[967:960] : wt0_sd_data[967:960];
  assign _01442_ = _05949_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6562" *) wt_pre_data[959:952] : wt0_sd_data[959:952];
  assign _01441_ = _05948_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6552" *) wt_pre_data[951:944] : wt0_sd_data[951:944];
  assign _01440_ = _05947_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6542" *) wt_pre_data[943:936] : wt0_sd_data[943:936];
  assign _01439_ = _05946_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6532" *) wt_pre_data[935:928] : wt0_sd_data[935:928];
  assign _01438_ = _05945_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6522" *) wt_pre_data[927:920] : wt0_sd_data[927:920];
  assign _01437_ = _05944_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6512" *) wt_pre_data[919:912] : wt0_sd_data[919:912];
  assign _01436_ = _05943_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6502" *) wt_pre_data[911:904] : wt0_sd_data[911:904];
  assign _01435_ = _05942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6492" *) wt_pre_data[903:896] : wt0_sd_data[903:896];
  assign _01434_ = _05941_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6482" *) wt_pre_data[895:888] : wt0_sd_data[895:888];
  assign _01433_ = _05940_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6472" *) wt_pre_data[887:880] : wt0_sd_data[887:880];
  assign _01431_ = _05939_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6462" *) wt_pre_data[879:872] : wt0_sd_data[879:872];
  assign _01430_ = _05938_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6452" *) wt_pre_data[871:864] : wt0_sd_data[871:864];
  assign _01429_ = _05937_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6442" *) wt_pre_data[863:856] : wt0_sd_data[863:856];
  assign _01428_ = _05936_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6432" *) wt_pre_data[855:848] : wt0_sd_data[855:848];
  assign _01427_ = _05935_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6422" *) wt_pre_data[847:840] : wt0_sd_data[847:840];
  assign _01426_ = _05934_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6412" *) wt_pre_data[839:832] : wt0_sd_data[839:832];
  assign _01425_ = _05933_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6402" *) wt_pre_data[831:824] : wt0_sd_data[831:824];
  assign _01424_ = _05932_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6392" *) wt_pre_data[823:816] : wt0_sd_data[823:816];
  assign _01423_ = _05931_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6382" *) wt_pre_data[815:808] : wt0_sd_data[815:808];
  assign _01422_ = _05930_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6372" *) wt_pre_data[807:800] : wt0_sd_data[807:800];
  assign _01419_ = _05929_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6362" *) wt_pre_data[799:792] : wt0_sd_data[799:792];
  assign _01418_ = _05928_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6352" *) wt_pre_data[791:784] : wt0_sd_data[791:784];
  assign _01417_ = _05927_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6342" *) wt_pre_data[783:776] : wt0_sd_data[783:776];
  assign _01416_ = _05926_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6332" *) wt_pre_data[775:768] : wt0_sd_data[775:768];
  assign _01415_ = _05925_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6322" *) wt_pre_data[767:760] : wt0_sd_data[767:760];
  assign _01414_ = _05924_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6312" *) wt_pre_data[759:752] : wt0_sd_data[759:752];
  assign _01413_ = _05923_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6302" *) wt_pre_data[751:744] : wt0_sd_data[751:744];
  assign _01412_ = _05922_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6292" *) wt_pre_data[743:736] : wt0_sd_data[743:736];
  assign _01411_ = _05921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6282" *) wt_pre_data[735:728] : wt0_sd_data[735:728];
  assign _01410_ = _05920_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6272" *) wt_pre_data[727:720] : wt0_sd_data[727:720];
  assign _01408_ = _05919_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6262" *) wt_pre_data[719:712] : wt0_sd_data[719:712];
  assign _01407_ = _05918_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6252" *) wt_pre_data[711:704] : wt0_sd_data[711:704];
  assign _01406_ = _05917_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6242" *) wt_pre_data[703:696] : wt0_sd_data[703:696];
  assign _01405_ = _05916_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6232" *) wt_pre_data[695:688] : wt0_sd_data[695:688];
  assign _01404_ = _05915_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6222" *) wt_pre_data[687:680] : wt0_sd_data[687:680];
  assign _01403_ = _05914_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6212" *) wt_pre_data[679:672] : wt0_sd_data[679:672];
  assign _01402_ = _05913_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6202" *) wt_pre_data[671:664] : wt0_sd_data[671:664];
  assign _01401_ = _05912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6192" *) wt_pre_data[663:656] : wt0_sd_data[663:656];
  assign _01400_ = _05911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6182" *) wt_pre_data[655:648] : wt0_sd_data[655:648];
  assign _01399_ = _05910_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6172" *) wt_pre_data[647:640] : wt0_sd_data[647:640];
  assign _01397_ = _05909_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6162" *) wt_pre_data[639:632] : wt0_sd_data[639:632];
  assign _01396_ = _05908_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6152" *) wt_pre_data[631:624] : wt0_sd_data[631:624];
  assign _01395_ = _05907_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6142" *) wt_pre_data[623:616] : wt0_sd_data[623:616];
  assign _01394_ = _05906_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6132" *) wt_pre_data[615:608] : wt0_sd_data[615:608];
  assign _01393_ = _05905_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6122" *) wt_pre_data[607:600] : wt0_sd_data[607:600];
  assign _01392_ = _05904_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6112" *) wt_pre_data[599:592] : wt0_sd_data[599:592];
  assign _01391_ = _05903_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6102" *) wt_pre_data[591:584] : wt0_sd_data[591:584];
  assign _01390_ = _05902_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6092" *) wt_pre_data[583:576] : wt0_sd_data[583:576];
  assign _01389_ = _05901_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6082" *) wt_pre_data[575:568] : wt0_sd_data[575:568];
  assign _01388_ = _05900_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6072" *) wt_pre_data[567:560] : wt0_sd_data[567:560];
  assign _01386_ = _05899_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6062" *) wt_pre_data[559:552] : wt0_sd_data[559:552];
  assign _01385_ = _05898_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6052" *) wt_pre_data[551:544] : wt0_sd_data[551:544];
  assign _01384_ = _05897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6042" *) wt_pre_data[543:536] : wt0_sd_data[543:536];
  assign _01383_ = _05896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6032" *) wt_pre_data[535:528] : wt0_sd_data[535:528];
  assign _01382_ = _05895_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6022" *) wt_pre_data[527:520] : wt0_sd_data[527:520];
  assign _01381_ = _05894_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6012" *) wt_pre_data[519:512] : wt0_sd_data[519:512];
  assign _01380_ = _05893_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6002" *) wt_pre_data[511:504] : wt0_sd_data[511:504];
  assign _01379_ = _05892_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5992" *) wt_pre_data[503:496] : wt0_sd_data[503:496];
  assign _01378_ = _05891_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5982" *) wt_pre_data[495:488] : wt0_sd_data[495:488];
  assign _01377_ = _05890_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5972" *) wt_pre_data[487:480] : wt0_sd_data[487:480];
  assign _01375_ = _05889_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5962" *) wt_pre_data[479:472] : wt0_sd_data[479:472];
  assign _01374_ = _05888_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5952" *) wt_pre_data[471:464] : wt0_sd_data[471:464];
  assign _01373_ = _05887_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5942" *) wt_pre_data[463:456] : wt0_sd_data[463:456];
  assign _01372_ = _05886_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5932" *) wt_pre_data[455:448] : wt0_sd_data[455:448];
  assign _01371_ = _05885_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5922" *) wt_pre_data[447:440] : wt0_sd_data[447:440];
  assign _01370_ = _05884_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5912" *) wt_pre_data[439:432] : wt0_sd_data[439:432];
  assign _01369_ = _05883_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5902" *) wt_pre_data[431:424] : wt0_sd_data[431:424];
  assign _01368_ = _05882_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5892" *) wt_pre_data[423:416] : wt0_sd_data[423:416];
  assign _01367_ = _05881_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5882" *) wt_pre_data[415:408] : wt0_sd_data[415:408];
  assign _01366_ = _05880_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5872" *) wt_pre_data[407:400] : wt0_sd_data[407:400];
  assign _01364_ = _05879_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5862" *) wt_pre_data[399:392] : wt0_sd_data[399:392];
  assign _01363_ = _05878_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5852" *) wt_pre_data[391:384] : wt0_sd_data[391:384];
  assign _01362_ = _05877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5842" *) wt_pre_data[383:376] : wt0_sd_data[383:376];
  assign _01361_ = _05876_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5832" *) wt_pre_data[375:368] : wt0_sd_data[375:368];
  assign _01360_ = _05875_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5822" *) wt_pre_data[367:360] : wt0_sd_data[367:360];
  assign _01359_ = _05874_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5812" *) wt_pre_data[359:352] : wt0_sd_data[359:352];
  assign _01358_ = _05873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5802" *) wt_pre_data[351:344] : wt0_sd_data[351:344];
  assign _01357_ = _05872_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5792" *) wt_pre_data[343:336] : wt0_sd_data[343:336];
  assign _01356_ = _05871_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5782" *) wt_pre_data[335:328] : wt0_sd_data[335:328];
  assign _01355_ = _05870_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5772" *) wt_pre_data[327:320] : wt0_sd_data[327:320];
  assign _01353_ = _05869_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5762" *) wt_pre_data[319:312] : wt0_sd_data[319:312];
  assign _01352_ = _05868_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5752" *) wt_pre_data[311:304] : wt0_sd_data[311:304];
  assign _01351_ = _05867_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5742" *) wt_pre_data[303:296] : wt0_sd_data[303:296];
  assign _01350_ = _05866_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5732" *) wt_pre_data[295:288] : wt0_sd_data[295:288];
  assign _01349_ = _05865_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5722" *) wt_pre_data[287:280] : wt0_sd_data[287:280];
  assign _01348_ = _05864_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5712" *) wt_pre_data[279:272] : wt0_sd_data[279:272];
  assign _01347_ = _05863_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5702" *) wt_pre_data[271:264] : wt0_sd_data[271:264];
  assign _01346_ = _05862_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5692" *) wt_pre_data[263:256] : wt0_sd_data[263:256];
  assign _01345_ = _05861_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5682" *) wt_pre_data[255:248] : wt0_sd_data[255:248];
  assign _01344_ = _05860_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5672" *) wt_pre_data[247:240] : wt0_sd_data[247:240];
  assign _01342_ = _05859_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5662" *) wt_pre_data[239:232] : wt0_sd_data[239:232];
  assign _01341_ = _05858_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5652" *) wt_pre_data[231:224] : wt0_sd_data[231:224];
  assign _01340_ = _05857_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5642" *) wt_pre_data[223:216] : wt0_sd_data[223:216];
  assign _01339_ = _05856_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5632" *) wt_pre_data[215:208] : wt0_sd_data[215:208];
  assign _01338_ = _05855_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5622" *) wt_pre_data[207:200] : wt0_sd_data[207:200];
  assign _01337_ = _05854_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5612" *) wt_pre_data[199:192] : wt0_sd_data[199:192];
  assign _01336_ = _05853_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5602" *) wt_pre_data[191:184] : wt0_sd_data[191:184];
  assign _01335_ = _05852_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5592" *) wt_pre_data[183:176] : wt0_sd_data[183:176];
  assign _01334_ = _05851_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5582" *) wt_pre_data[175:168] : wt0_sd_data[175:168];
  assign _01333_ = _05850_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5572" *) wt_pre_data[167:160] : wt0_sd_data[167:160];
  assign _01331_ = _05849_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5562" *) wt_pre_data[159:152] : wt0_sd_data[159:152];
  assign _01330_ = _05848_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5552" *) wt_pre_data[151:144] : wt0_sd_data[151:144];
  assign _01329_ = _05847_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5542" *) wt_pre_data[143:136] : wt0_sd_data[143:136];
  assign _01328_ = _05846_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5532" *) wt_pre_data[135:128] : wt0_sd_data[135:128];
  assign _01327_ = _05845_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5522" *) wt_pre_data[127:120] : wt0_sd_data[127:120];
  assign _01326_ = _05844_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5512" *) wt_pre_data[119:112] : wt0_sd_data[119:112];
  assign _01325_ = _05843_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5502" *) wt_pre_data[111:104] : wt0_sd_data[111:104];
  assign _01324_ = _05842_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5492" *) wt_pre_data[103:96] : wt0_sd_data[103:96];
  assign _01443_ = _05841_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5482" *) wt_pre_data[95:88] : wt0_sd_data[95:88];
  assign _01432_ = _05840_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5472" *) wt_pre_data[87:80] : wt0_sd_data[87:80];
  assign _01420_ = _05839_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5462" *) wt_pre_data[79:72] : wt0_sd_data[79:72];
  assign _01409_ = _05838_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5452" *) wt_pre_data[71:64] : wt0_sd_data[71:64];
  assign _01398_ = _05837_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5442" *) wt_pre_data[63:56] : wt0_sd_data[63:56];
  assign _01387_ = _05836_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5432" *) wt_pre_data[55:48] : wt0_sd_data[55:48];
  assign _01376_ = _05835_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5422" *) wt_pre_data[47:40] : wt0_sd_data[47:40];
  assign _01365_ = _05834_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5412" *) wt_pre_data[39:32] : wt0_sd_data[39:32];
  assign _01354_ = _05833_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5402" *) wt_pre_data[31:24] : wt0_sd_data[31:24];
  assign _01343_ = _05832_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5392" *) wt_pre_data[23:16] : wt0_sd_data[23:16];
  assign _01332_ = _05831_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5382" *) wt_pre_data[15:8] : wt0_sd_data[15:8];
  assign _01421_ = _05830_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5372" *) wt_pre_data[7:0] : wt0_sd_data[7:0];
  assign _01451_ = _05829_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5362" *) wt_pre_nan : wt0_sd_nan;
  assign _01449_ = _05829_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5352" *) wt_pre_exp : wt0_sd_exp;
  assign _01450_ = _05829_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5342" *) wt_pre_mask : wt0_sd_mask;
  assign _01452_ = wt_pre_sel[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5332" *) wt_pre_nz : wt0_sd_nz;
  assign _03289_ = _05828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5303" *) wt_pre_data_w[1023:1016] : wt_pre_data[1023:1016];
  assign _03288_ = _05827_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5293" *) wt_pre_data_w[1015:1008] : wt_pre_data[1015:1008];
  assign _03287_ = _05826_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5283" *) wt_pre_data_w[1007:1000] : wt_pre_data[1007:1000];
  assign _03414_ = _05825_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5273" *) wt_pre_data_w[999:992] : wt_pre_data[999:992];
  assign _03413_ = _05824_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5263" *) wt_pre_data_w[991:984] : wt_pre_data[991:984];
  assign _03412_ = _05823_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5253" *) wt_pre_data_w[983:976] : wt_pre_data[983:976];
  assign _03411_ = _05822_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5243" *) wt_pre_data_w[975:968] : wt_pre_data[975:968];
  assign _03410_ = _05821_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5233" *) wt_pre_data_w[967:960] : wt_pre_data[967:960];
  assign _03408_ = _05820_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5223" *) wt_pre_data_w[959:952] : wt_pre_data[959:952];
  assign _03407_ = _05819_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5213" *) wt_pre_data_w[951:944] : wt_pre_data[951:944];
  assign _03406_ = _05818_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5203" *) wt_pre_data_w[943:936] : wt_pre_data[943:936];
  assign _03405_ = _05817_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5193" *) wt_pre_data_w[935:928] : wt_pre_data[935:928];
  assign _03404_ = _05816_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5183" *) wt_pre_data_w[927:920] : wt_pre_data[927:920];
  assign _03403_ = _05815_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5173" *) wt_pre_data_w[919:912] : wt_pre_data[919:912];
  assign _03402_ = _05814_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5163" *) wt_pre_data_w[911:904] : wt_pre_data[911:904];
  assign _03401_ = _05813_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5153" *) wt_pre_data_w[903:896] : wt_pre_data[903:896];
  assign _03400_ = _05812_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5143" *) wt_pre_data_w[895:888] : wt_pre_data[895:888];
  assign _03399_ = _05811_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5133" *) wt_pre_data_w[887:880] : wt_pre_data[887:880];
  assign _03397_ = _05810_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5123" *) wt_pre_data_w[879:872] : wt_pre_data[879:872];
  assign _03396_ = _05809_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5113" *) wt_pre_data_w[871:864] : wt_pre_data[871:864];
  assign _03395_ = _05808_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5103" *) wt_pre_data_w[863:856] : wt_pre_data[863:856];
  assign _03394_ = _05807_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5093" *) wt_pre_data_w[855:848] : wt_pre_data[855:848];
  assign _03393_ = _05806_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5083" *) wt_pre_data_w[847:840] : wt_pre_data[847:840];
  assign _03392_ = _05805_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5073" *) wt_pre_data_w[839:832] : wt_pre_data[839:832];
  assign _03391_ = _05804_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5063" *) wt_pre_data_w[831:824] : wt_pre_data[831:824];
  assign _03390_ = _05803_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5053" *) wt_pre_data_w[823:816] : wt_pre_data[823:816];
  assign _03389_ = _05802_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5043" *) wt_pre_data_w[815:808] : wt_pre_data[815:808];
  assign _03388_ = _05801_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5033" *) wt_pre_data_w[807:800] : wt_pre_data[807:800];
  assign _03385_ = _05800_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5023" *) wt_pre_data_w[799:792] : wt_pre_data[799:792];
  assign _03384_ = _05799_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5013" *) wt_pre_data_w[791:784] : wt_pre_data[791:784];
  assign _03383_ = _05798_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5003" *) wt_pre_data_w[783:776] : wt_pre_data[783:776];
  assign _03382_ = _05797_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4993" *) wt_pre_data_w[775:768] : wt_pre_data[775:768];
  assign _03381_ = _05796_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4983" *) wt_pre_data_w[767:760] : wt_pre_data[767:760];
  assign _03380_ = _05795_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4973" *) wt_pre_data_w[759:752] : wt_pre_data[759:752];
  assign _03379_ = _05794_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4963" *) wt_pre_data_w[751:744] : wt_pre_data[751:744];
  assign _03378_ = _05793_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4953" *) wt_pre_data_w[743:736] : wt_pre_data[743:736];
  assign _03377_ = _05792_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4943" *) wt_pre_data_w[735:728] : wt_pre_data[735:728];
  assign _03376_ = _05791_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4933" *) wt_pre_data_w[727:720] : wt_pre_data[727:720];
  assign _03374_ = _05790_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4923" *) wt_pre_data_w[719:712] : wt_pre_data[719:712];
  assign _03373_ = _05789_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4913" *) wt_pre_data_w[711:704] : wt_pre_data[711:704];
  assign _03372_ = _05788_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4903" *) wt_pre_data_w[703:696] : wt_pre_data[703:696];
  assign _03371_ = _05787_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4893" *) wt_pre_data_w[695:688] : wt_pre_data[695:688];
  assign _03370_ = _05786_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4883" *) wt_pre_data_w[687:680] : wt_pre_data[687:680];
  assign _03369_ = _05785_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4873" *) wt_pre_data_w[679:672] : wt_pre_data[679:672];
  assign _03368_ = _05784_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4863" *) wt_pre_data_w[671:664] : wt_pre_data[671:664];
  assign _03367_ = _05783_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4853" *) wt_pre_data_w[663:656] : wt_pre_data[663:656];
  assign _03366_ = _05782_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4843" *) wt_pre_data_w[655:648] : wt_pre_data[655:648];
  assign _03365_ = _05781_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4833" *) wt_pre_data_w[647:640] : wt_pre_data[647:640];
  assign _03363_ = _05780_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4823" *) wt_pre_data_w[639:632] : wt_pre_data[639:632];
  assign _03362_ = _05779_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4813" *) wt_pre_data_w[631:624] : wt_pre_data[631:624];
  assign _03361_ = _05778_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4803" *) wt_pre_data_w[623:616] : wt_pre_data[623:616];
  assign _03360_ = _05777_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4793" *) wt_pre_data_w[615:608] : wt_pre_data[615:608];
  assign _03359_ = _05776_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4783" *) wt_pre_data_w[607:600] : wt_pre_data[607:600];
  assign _03358_ = _05775_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4773" *) wt_pre_data_w[599:592] : wt_pre_data[599:592];
  assign _03357_ = _05774_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4763" *) wt_pre_data_w[591:584] : wt_pre_data[591:584];
  assign _03356_ = _05773_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4753" *) wt_pre_data_w[583:576] : wt_pre_data[583:576];
  assign _03355_ = _05772_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4743" *) wt_pre_data_w[575:568] : wt_pre_data[575:568];
  assign _03354_ = _05771_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4733" *) wt_pre_data_w[567:560] : wt_pre_data[567:560];
  assign _03352_ = _05770_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4723" *) wt_pre_data_w[559:552] : wt_pre_data[559:552];
  assign _03351_ = _05769_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4713" *) wt_pre_data_w[551:544] : wt_pre_data[551:544];
  assign _03350_ = _05768_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4703" *) wt_pre_data_w[543:536] : wt_pre_data[543:536];
  assign _03349_ = _05767_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4693" *) wt_pre_data_w[535:528] : wt_pre_data[535:528];
  assign _03348_ = _05766_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4683" *) wt_pre_data_w[527:520] : wt_pre_data[527:520];
  assign _03347_ = _05765_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4673" *) wt_pre_data_w[519:512] : wt_pre_data[519:512];
  assign _03346_ = _05764_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4663" *) wt_pre_data_w[511:504] : wt_pre_data[511:504];
  assign _03345_ = _05763_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4653" *) wt_pre_data_w[503:496] : wt_pre_data[503:496];
  assign _03344_ = _05762_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4643" *) wt_pre_data_w[495:488] : wt_pre_data[495:488];
  assign _03343_ = _05761_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4633" *) wt_pre_data_w[487:480] : wt_pre_data[487:480];
  assign _03341_ = _05760_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4623" *) wt_pre_data_w[479:472] : wt_pre_data[479:472];
  assign _03340_ = _05759_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4613" *) wt_pre_data_w[471:464] : wt_pre_data[471:464];
  assign _03339_ = _05758_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4603" *) wt_pre_data_w[463:456] : wt_pre_data[463:456];
  assign _03338_ = _05757_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4593" *) wt_pre_data_w[455:448] : wt_pre_data[455:448];
  assign _03337_ = _05756_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4583" *) wt_pre_data_w[447:440] : wt_pre_data[447:440];
  assign _03336_ = _05755_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4573" *) wt_pre_data_w[439:432] : wt_pre_data[439:432];
  assign _03335_ = _05754_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4563" *) wt_pre_data_w[431:424] : wt_pre_data[431:424];
  assign _03334_ = _05753_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4553" *) wt_pre_data_w[423:416] : wt_pre_data[423:416];
  assign _03333_ = _05752_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4543" *) wt_pre_data_w[415:408] : wt_pre_data[415:408];
  assign _03332_ = _05751_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4533" *) wt_pre_data_w[407:400] : wt_pre_data[407:400];
  assign _03330_ = _05750_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4523" *) wt_pre_data_w[399:392] : wt_pre_data[399:392];
  assign _03329_ = _05749_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4513" *) wt_pre_data_w[391:384] : wt_pre_data[391:384];
  assign _03328_ = _05748_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4503" *) wt_pre_data_w[383:376] : wt_pre_data[383:376];
  assign _03327_ = _05747_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4493" *) wt_pre_data_w[375:368] : wt_pre_data[375:368];
  assign _03326_ = _05746_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4483" *) wt_pre_data_w[367:360] : wt_pre_data[367:360];
  assign _03325_ = _05745_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4473" *) wt_pre_data_w[359:352] : wt_pre_data[359:352];
  assign _03324_ = _05744_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4463" *) wt_pre_data_w[351:344] : wt_pre_data[351:344];
  assign _03323_ = _05743_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4453" *) wt_pre_data_w[343:336] : wt_pre_data[343:336];
  assign _03322_ = _05742_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4443" *) wt_pre_data_w[335:328] : wt_pre_data[335:328];
  assign _03321_ = _05741_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4433" *) wt_pre_data_w[327:320] : wt_pre_data[327:320];
  assign _03319_ = _05740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4423" *) wt_pre_data_w[319:312] : wt_pre_data[319:312];
  assign _03318_ = _05739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4413" *) wt_pre_data_w[311:304] : wt_pre_data[311:304];
  assign _03317_ = _05738_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4403" *) wt_pre_data_w[303:296] : wt_pre_data[303:296];
  assign _03316_ = _05737_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4393" *) wt_pre_data_w[295:288] : wt_pre_data[295:288];
  assign _03315_ = _05736_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4383" *) wt_pre_data_w[287:280] : wt_pre_data[287:280];
  assign _03314_ = _05735_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4373" *) wt_pre_data_w[279:272] : wt_pre_data[279:272];
  assign _03313_ = _05734_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4363" *) wt_pre_data_w[271:264] : wt_pre_data[271:264];
  assign _03312_ = _05733_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4353" *) wt_pre_data_w[263:256] : wt_pre_data[263:256];
  assign _03311_ = _05732_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4343" *) wt_pre_data_w[255:248] : wt_pre_data[255:248];
  assign _03310_ = _05731_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4333" *) wt_pre_data_w[247:240] : wt_pre_data[247:240];
  assign _03308_ = _05730_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4323" *) wt_pre_data_w[239:232] : wt_pre_data[239:232];
  assign _03307_ = _05729_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4313" *) wt_pre_data_w[231:224] : wt_pre_data[231:224];
  assign _03306_ = _05728_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4303" *) wt_pre_data_w[223:216] : wt_pre_data[223:216];
  assign _03305_ = _05727_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4293" *) wt_pre_data_w[215:208] : wt_pre_data[215:208];
  assign _03304_ = _05726_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4283" *) wt_pre_data_w[207:200] : wt_pre_data[207:200];
  assign _03303_ = _05725_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4273" *) wt_pre_data_w[199:192] : wt_pre_data[199:192];
  assign _03302_ = _05724_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4263" *) wt_pre_data_w[191:184] : wt_pre_data[191:184];
  assign _03301_ = _05723_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4253" *) wt_pre_data_w[183:176] : wt_pre_data[183:176];
  assign _03300_ = _05722_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4243" *) wt_pre_data_w[175:168] : wt_pre_data[175:168];
  assign _03299_ = _05721_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4233" *) wt_pre_data_w[167:160] : wt_pre_data[167:160];
  assign _03297_ = _05720_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4223" *) wt_pre_data_w[159:152] : wt_pre_data[159:152];
  assign _03296_ = _05719_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4213" *) wt_pre_data_w[151:144] : wt_pre_data[151:144];
  assign _03295_ = _05718_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4203" *) wt_pre_data_w[143:136] : wt_pre_data[143:136];
  assign _03294_ = _05717_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4193" *) wt_pre_data_w[135:128] : wt_pre_data[135:128];
  assign _03293_ = _05716_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4183" *) wt_pre_data_w[127:120] : wt_pre_data[127:120];
  assign _03292_ = _05715_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4173" *) wt_pre_data_w[119:112] : wt_pre_data[119:112];
  assign _03291_ = _05714_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4163" *) wt_pre_data_w[111:104] : wt_pre_data[111:104];
  assign _03290_ = _05713_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4153" *) wt_pre_data_w[103:96] : wt_pre_data[103:96];
  assign _03409_ = _05712_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4143" *) wt_pre_data_w[95:88] : wt_pre_data[95:88];
  assign _03398_ = _05711_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4133" *) wt_pre_data_w[87:80] : wt_pre_data[87:80];
  assign _03386_ = _05710_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4123" *) wt_pre_data_w[79:72] : wt_pre_data[79:72];
  assign _03375_ = _05709_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4113" *) wt_pre_data_w[71:64] : wt_pre_data[71:64];
  assign _03364_ = _05708_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4103" *) wt_pre_data_w[63:56] : wt_pre_data[63:56];
  assign _03353_ = _05707_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4093" *) wt_pre_data_w[55:48] : wt_pre_data[55:48];
  assign _03342_ = _05706_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4083" *) wt_pre_data_w[47:40] : wt_pre_data[47:40];
  assign _03331_ = _05705_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4073" *) wt_pre_data_w[39:32] : wt_pre_data[39:32];
  assign _03320_ = _05704_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4063" *) wt_pre_data_w[31:24] : wt_pre_data[31:24];
  assign _03309_ = _05703_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4053" *) wt_pre_data_w[23:16] : wt_pre_data[23:16];
  assign _03298_ = _05702_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4043" *) wt_pre_data_w[15:8] : wt_pre_data[15:8];
  assign _03387_ = _05701_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4033" *) wt_pre_data_w[7:0] : wt_pre_data[7:0];
  assign _03417_ = _05700_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4023" *) in_wt_nan : wt_pre_nan;
  assign _03415_ = _05700_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4013" *) wt_pre_exp_w : wt_pre_exp;
  assign _03416_ = _05700_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:4003" *) { wt_pre_nz_w[126], wt_pre_nz_w[124], wt_pre_nz_w[122], wt_pre_nz_w[120], wt_pre_nz_w[118], wt_pre_nz_w[116], wt_pre_nz_w[114], wt_pre_nz_w[112], wt_pre_nz_w[110], wt_pre_nz_w[108], wt_pre_nz_w[106], wt_pre_nz_w[104], wt_pre_nz_w[102], wt_pre_nz_w[100], wt_pre_nz_w[98], wt_pre_nz_w[96], wt_pre_nz_w[94], wt_pre_nz_w[92], wt_pre_nz_w[90], wt_pre_nz_w[88], wt_pre_nz_w[86], wt_pre_nz_w[84], wt_pre_nz_w[82], wt_pre_nz_w[80], wt_pre_nz_w[78], wt_pre_nz_w[76], wt_pre_nz_w[74], wt_pre_nz_w[72], wt_pre_nz_w[70], wt_pre_nz_w[68], wt_pre_nz_w[66], wt_pre_nz_w[64], wt_pre_nz_w[62], wt_pre_nz_w[60], wt_pre_nz_w[58], wt_pre_nz_w[56], wt_pre_nz_w[54], wt_pre_nz_w[52], wt_pre_nz_w[50], wt_pre_nz_w[48], wt_pre_nz_w[46], wt_pre_nz_w[44], wt_pre_nz_w[42], wt_pre_nz_w[40], wt_pre_nz_w[38], wt_pre_nz_w[36], wt_pre_nz_w[34], wt_pre_nz_w[32], wt_pre_nz_w[30], wt_pre_nz_w[28], wt_pre_nz_w[26], wt_pre_nz_w[24], wt_pre_nz_w[22], wt_pre_nz_w[20], wt_pre_nz_w[18], wt_pre_nz_w[16], wt_pre_nz_w[14], wt_pre_nz_w[12], wt_pre_nz_w[10], wt_pre_nz_w[8], wt_pre_nz_w[6], wt_pre_nz_w[4], wt_pre_nz_w[2], wt_pre_nz_w[0] } : wt_pre_mask;
  assign _03418_ = in_wt_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3993" *) wt_pre_nz_w : wt_pre_nz;
  assign _00001_ = cfg_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1848" *) { cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16, cfg_is_int16 } : cfg_is_int16_d1;
  assign _00000_ = cfg_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1787" *) { cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16 } : cfg_is_fp16_d1;
  assign _00002_ = cfg_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:1726" *) { cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8, cfg_is_int8 } : cfg_is_int8_d1;
  assign _07947_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *) { in_wt_data127[2], in_wt_data127[3], in_wt_data127[4], in_wt_data127[5], in_wt_data127[6] };
  assign _07948_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *) { in_wt_data125[2], in_wt_data125[3], in_wt_data125[4], in_wt_data125[5], in_wt_data125[6] };
  assign _07949_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *) { in_wt_data123[2], in_wt_data123[3], in_wt_data123[4], in_wt_data123[5], in_wt_data123[6] };
  assign _07950_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *) { in_wt_data121[2], in_wt_data121[3], in_wt_data121[4], in_wt_data121[5], in_wt_data121[6] };
  assign _07951_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *) { in_wt_data119[2], in_wt_data119[3], in_wt_data119[4], in_wt_data119[5], in_wt_data119[6] };
  assign _07952_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *) { in_wt_data117[2], in_wt_data117[3], in_wt_data117[4], in_wt_data117[5], in_wt_data117[6] };
  assign _07953_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *) { in_wt_data115[2], in_wt_data115[3], in_wt_data115[4], in_wt_data115[5], in_wt_data115[6] };
  assign _07954_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *) { in_wt_data113[2], in_wt_data113[3], in_wt_data113[4], in_wt_data113[5], in_wt_data113[6] };
  assign _07955_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *) { in_wt_data111[2], in_wt_data111[3], in_wt_data111[4], in_wt_data111[5], in_wt_data111[6] };
  assign _07956_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *) { in_wt_data109[2], in_wt_data109[3], in_wt_data109[4], in_wt_data109[5], in_wt_data109[6] };
  assign _07957_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *) { in_wt_data107[2], in_wt_data107[3], in_wt_data107[4], in_wt_data107[5], in_wt_data107[6] };
  assign _07958_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *) { in_wt_data105[2], in_wt_data105[3], in_wt_data105[4], in_wt_data105[5], in_wt_data105[6] };
  assign _07959_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *) { in_wt_data103[2], in_wt_data103[3], in_wt_data103[4], in_wt_data103[5], in_wt_data103[6] };
  assign _07960_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *) { in_wt_data101[2], in_wt_data101[3], in_wt_data101[4], in_wt_data101[5], in_wt_data101[6] };
  assign _07961_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *) { in_wt_data99[2], in_wt_data99[3], in_wt_data99[4], in_wt_data99[5], in_wt_data99[6] };
  assign _07962_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *) { in_wt_data97[2], in_wt_data97[3], in_wt_data97[4], in_wt_data97[5], in_wt_data97[6] };
  assign _07963_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *) { in_wt_data95[2], in_wt_data95[3], in_wt_data95[4], in_wt_data95[5], in_wt_data95[6] };
  assign _07964_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *) { in_wt_data93[2], in_wt_data93[3], in_wt_data93[4], in_wt_data93[5], in_wt_data93[6] };
  assign _07965_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *) { in_wt_data91[2], in_wt_data91[3], in_wt_data91[4], in_wt_data91[5], in_wt_data91[6] };
  assign _07966_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *) { in_wt_data89[2], in_wt_data89[3], in_wt_data89[4], in_wt_data89[5], in_wt_data89[6] };
  assign _07967_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *) { in_wt_data87[2], in_wt_data87[3], in_wt_data87[4], in_wt_data87[5], in_wt_data87[6] };
  assign _07968_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *) { in_wt_data85[2], in_wt_data85[3], in_wt_data85[4], in_wt_data85[5], in_wt_data85[6] };
  assign _07969_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *) { in_wt_data83[2], in_wt_data83[3], in_wt_data83[4], in_wt_data83[5], in_wt_data83[6] };
  assign _07970_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *) { in_wt_data81[2], in_wt_data81[3], in_wt_data81[4], in_wt_data81[5], in_wt_data81[6] };
  assign _07971_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *) { in_wt_data79[2], in_wt_data79[3], in_wt_data79[4], in_wt_data79[5], in_wt_data79[6] };
  assign _07972_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *) { in_wt_data77[2], in_wt_data77[3], in_wt_data77[4], in_wt_data77[5], in_wt_data77[6] };
  assign _07973_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *) { in_wt_data75[2], in_wt_data75[3], in_wt_data75[4], in_wt_data75[5], in_wt_data75[6] };
  assign _07974_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *) { in_wt_data73[2], in_wt_data73[3], in_wt_data73[4], in_wt_data73[5], in_wt_data73[6] };
  assign _07975_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *) { in_wt_data71[2], in_wt_data71[3], in_wt_data71[4], in_wt_data71[5], in_wt_data71[6] };
  assign _07976_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *) { in_wt_data69[2], in_wt_data69[3], in_wt_data69[4], in_wt_data69[5], in_wt_data69[6] };
  assign _07977_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *) { in_wt_data67[2], in_wt_data67[3], in_wt_data67[4], in_wt_data67[5], in_wt_data67[6] };
  assign _07978_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *) { in_wt_data65[2], in_wt_data65[3], in_wt_data65[4], in_wt_data65[5], in_wt_data65[6] };
  assign _07979_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *) { in_wt_data63[2], in_wt_data63[3], in_wt_data63[4], in_wt_data63[5], in_wt_data63[6] };
  assign _07980_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *) { in_wt_data61[2], in_wt_data61[3], in_wt_data61[4], in_wt_data61[5], in_wt_data61[6] };
  assign _07981_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *) { in_wt_data59[2], in_wt_data59[3], in_wt_data59[4], in_wt_data59[5], in_wt_data59[6] };
  assign _07982_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *) { in_wt_data57[2], in_wt_data57[3], in_wt_data57[4], in_wt_data57[5], in_wt_data57[6] };
  assign _07983_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *) { in_wt_data55[2], in_wt_data55[3], in_wt_data55[4], in_wt_data55[5], in_wt_data55[6] };
  assign _07984_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *) { in_wt_data53[2], in_wt_data53[3], in_wt_data53[4], in_wt_data53[5], in_wt_data53[6] };
  assign _07985_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *) { in_wt_data51[2], in_wt_data51[3], in_wt_data51[4], in_wt_data51[5], in_wt_data51[6] };
  assign _07986_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *) { in_wt_data49[2], in_wt_data49[3], in_wt_data49[4], in_wt_data49[5], in_wt_data49[6] };
  assign _07987_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *) { in_wt_data47[2], in_wt_data47[3], in_wt_data47[4], in_wt_data47[5], in_wt_data47[6] };
  assign _07988_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *) { in_wt_data45[2], in_wt_data45[3], in_wt_data45[4], in_wt_data45[5], in_wt_data45[6] };
  assign _07989_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *) { in_wt_data43[2], in_wt_data43[3], in_wt_data43[4], in_wt_data43[5], in_wt_data43[6] };
  assign _07990_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *) { in_wt_data41[2], in_wt_data41[3], in_wt_data41[4], in_wt_data41[5], in_wt_data41[6] };
  assign _07991_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *) { in_wt_data39[2], in_wt_data39[3], in_wt_data39[4], in_wt_data39[5], in_wt_data39[6] };
  assign _07992_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *) { in_wt_data37[2], in_wt_data37[3], in_wt_data37[4], in_wt_data37[5], in_wt_data37[6] };
  assign _07993_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *) { in_wt_data35[2], in_wt_data35[3], in_wt_data35[4], in_wt_data35[5], in_wt_data35[6] };
  assign _07994_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *) { in_wt_data33[2], in_wt_data33[3], in_wt_data33[4], in_wt_data33[5], in_wt_data33[6] };
  assign _07995_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *) { in_wt_data31[2], in_wt_data31[3], in_wt_data31[4], in_wt_data31[5], in_wt_data31[6] };
  assign _07996_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *) { in_wt_data29[2], in_wt_data29[3], in_wt_data29[4], in_wt_data29[5], in_wt_data29[6] };
  assign _07997_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *) { in_wt_data27[2], in_wt_data27[3], in_wt_data27[4], in_wt_data27[5], in_wt_data27[6] };
  assign _07998_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *) { in_wt_data25[2], in_wt_data25[3], in_wt_data25[4], in_wt_data25[5], in_wt_data25[6] };
  assign _07999_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *) { in_wt_data23[2], in_wt_data23[3], in_wt_data23[4], in_wt_data23[5], in_wt_data23[6] };
  assign _08000_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *) { in_wt_data21[2], in_wt_data21[3], in_wt_data21[4], in_wt_data21[5], in_wt_data21[6] };
  assign _08001_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *) { in_wt_data19[2], in_wt_data19[3], in_wt_data19[4], in_wt_data19[5], in_wt_data19[6] };
  assign _08002_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *) { in_wt_data17[2], in_wt_data17[3], in_wt_data17[4], in_wt_data17[5], in_wt_data17[6] };
  assign _08003_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *) { in_wt_data15[2], in_wt_data15[3], in_wt_data15[4], in_wt_data15[5], in_wt_data15[6] };
  assign _08004_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *) { in_wt_data13[2], in_wt_data13[3], in_wt_data13[4], in_wt_data13[5], in_wt_data13[6] };
  assign _08005_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *) { in_wt_data11[2], in_wt_data11[3], in_wt_data11[4], in_wt_data11[5], in_wt_data11[6] };
  assign _08006_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *) { in_wt_data9[2], in_wt_data9[3], in_wt_data9[4], in_wt_data9[5], in_wt_data9[6] };
  assign _08007_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *) { in_wt_data7[2], in_wt_data7[3], in_wt_data7[4], in_wt_data7[5], in_wt_data7[6] };
  assign _08008_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *) { in_wt_data5[2], in_wt_data5[3], in_wt_data5[4], in_wt_data5[5], in_wt_data5[6] };
  assign _08009_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *) { in_wt_data3[2], in_wt_data3[3], in_wt_data3[4], in_wt_data3[5], in_wt_data3[6] };
  assign _08010_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *) { in_wt_data1[2], in_wt_data1[3], in_wt_data1[4], in_wt_data1[5], in_wt_data1[6] };
  assign _08011_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *) { in_dat_data127[2], in_dat_data127[3], in_dat_data127[4], in_dat_data127[5], in_dat_data127[6] };
  assign _08012_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *) { in_dat_data125[2], in_dat_data125[3], in_dat_data125[4], in_dat_data125[5], in_dat_data125[6] };
  assign _08013_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *) { in_dat_data123[2], in_dat_data123[3], in_dat_data123[4], in_dat_data123[5], in_dat_data123[6] };
  assign _08014_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *) { in_dat_data121[2], in_dat_data121[3], in_dat_data121[4], in_dat_data121[5], in_dat_data121[6] };
  assign _08015_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *) { in_dat_data119[2], in_dat_data119[3], in_dat_data119[4], in_dat_data119[5], in_dat_data119[6] };
  assign _08016_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *) { in_dat_data117[2], in_dat_data117[3], in_dat_data117[4], in_dat_data117[5], in_dat_data117[6] };
  assign _08017_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *) { in_dat_data115[2], in_dat_data115[3], in_dat_data115[4], in_dat_data115[5], in_dat_data115[6] };
  assign _08018_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *) { in_dat_data113[2], in_dat_data113[3], in_dat_data113[4], in_dat_data113[5], in_dat_data113[6] };
  assign _08019_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *) { in_dat_data111[2], in_dat_data111[3], in_dat_data111[4], in_dat_data111[5], in_dat_data111[6] };
  assign _08020_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *) { in_dat_data109[2], in_dat_data109[3], in_dat_data109[4], in_dat_data109[5], in_dat_data109[6] };
  assign _08021_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *) { in_dat_data107[2], in_dat_data107[3], in_dat_data107[4], in_dat_data107[5], in_dat_data107[6] };
  assign _08022_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *) { in_dat_data105[2], in_dat_data105[3], in_dat_data105[4], in_dat_data105[5], in_dat_data105[6] };
  assign _08023_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *) { in_dat_data103[2], in_dat_data103[3], in_dat_data103[4], in_dat_data103[5], in_dat_data103[6] };
  assign _08024_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *) { in_dat_data101[2], in_dat_data101[3], in_dat_data101[4], in_dat_data101[5], in_dat_data101[6] };
  assign _08025_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *) { in_dat_data99[2], in_dat_data99[3], in_dat_data99[4], in_dat_data99[5], in_dat_data99[6] };
  assign _08026_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *) { in_dat_data97[2], in_dat_data97[3], in_dat_data97[4], in_dat_data97[5], in_dat_data97[6] };
  assign _08027_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *) { in_dat_data95[2], in_dat_data95[3], in_dat_data95[4], in_dat_data95[5], in_dat_data95[6] };
  assign _08028_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *) { in_dat_data93[2], in_dat_data93[3], in_dat_data93[4], in_dat_data93[5], in_dat_data93[6] };
  assign _08029_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *) { in_dat_data91[2], in_dat_data91[3], in_dat_data91[4], in_dat_data91[5], in_dat_data91[6] };
  assign _08030_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *) { in_dat_data89[2], in_dat_data89[3], in_dat_data89[4], in_dat_data89[5], in_dat_data89[6] };
  assign _08031_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *) { in_dat_data87[2], in_dat_data87[3], in_dat_data87[4], in_dat_data87[5], in_dat_data87[6] };
  assign _08032_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *) { in_dat_data85[2], in_dat_data85[3], in_dat_data85[4], in_dat_data85[5], in_dat_data85[6] };
  assign _08033_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *) { in_dat_data83[2], in_dat_data83[3], in_dat_data83[4], in_dat_data83[5], in_dat_data83[6] };
  assign _08034_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *) { in_dat_data81[2], in_dat_data81[3], in_dat_data81[4], in_dat_data81[5], in_dat_data81[6] };
  assign _08035_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *) { in_dat_data79[2], in_dat_data79[3], in_dat_data79[4], in_dat_data79[5], in_dat_data79[6] };
  assign _08036_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *) { in_dat_data77[2], in_dat_data77[3], in_dat_data77[4], in_dat_data77[5], in_dat_data77[6] };
  assign _08037_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *) { in_dat_data75[2], in_dat_data75[3], in_dat_data75[4], in_dat_data75[5], in_dat_data75[6] };
  assign _08038_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *) { in_dat_data73[2], in_dat_data73[3], in_dat_data73[4], in_dat_data73[5], in_dat_data73[6] };
  assign _08039_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *) { in_dat_data71[2], in_dat_data71[3], in_dat_data71[4], in_dat_data71[5], in_dat_data71[6] };
  assign _08040_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *) { in_dat_data69[2], in_dat_data69[3], in_dat_data69[4], in_dat_data69[5], in_dat_data69[6] };
  assign _08041_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *) { in_dat_data67[2], in_dat_data67[3], in_dat_data67[4], in_dat_data67[5], in_dat_data67[6] };
  assign _08042_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *) { in_dat_data65[2], in_dat_data65[3], in_dat_data65[4], in_dat_data65[5], in_dat_data65[6] };
  assign _08043_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *) { in_dat_data63[2], in_dat_data63[3], in_dat_data63[4], in_dat_data63[5], in_dat_data63[6] };
  assign _08044_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *) { in_dat_data61[2], in_dat_data61[3], in_dat_data61[4], in_dat_data61[5], in_dat_data61[6] };
  assign _08045_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *) { in_dat_data59[2], in_dat_data59[3], in_dat_data59[4], in_dat_data59[5], in_dat_data59[6] };
  assign _08046_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *) { in_dat_data57[2], in_dat_data57[3], in_dat_data57[4], in_dat_data57[5], in_dat_data57[6] };
  assign _08047_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *) { in_dat_data55[2], in_dat_data55[3], in_dat_data55[4], in_dat_data55[5], in_dat_data55[6] };
  assign _08048_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *) { in_dat_data53[2], in_dat_data53[3], in_dat_data53[4], in_dat_data53[5], in_dat_data53[6] };
  assign _08049_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *) { in_dat_data51[2], in_dat_data51[3], in_dat_data51[4], in_dat_data51[5], in_dat_data51[6] };
  assign _08050_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *) { in_dat_data49[2], in_dat_data49[3], in_dat_data49[4], in_dat_data49[5], in_dat_data49[6] };
  assign _08051_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *) { in_dat_data47[2], in_dat_data47[3], in_dat_data47[4], in_dat_data47[5], in_dat_data47[6] };
  assign _08052_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *) { in_dat_data45[2], in_dat_data45[3], in_dat_data45[4], in_dat_data45[5], in_dat_data45[6] };
  assign _08053_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *) { in_dat_data43[2], in_dat_data43[3], in_dat_data43[4], in_dat_data43[5], in_dat_data43[6] };
  assign _08054_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *) { in_dat_data41[2], in_dat_data41[3], in_dat_data41[4], in_dat_data41[5], in_dat_data41[6] };
  assign _08055_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *) { in_dat_data39[2], in_dat_data39[3], in_dat_data39[4], in_dat_data39[5], in_dat_data39[6] };
  assign _08056_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *) { in_dat_data37[2], in_dat_data37[3], in_dat_data37[4], in_dat_data37[5], in_dat_data37[6] };
  assign _08057_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *) { in_dat_data35[2], in_dat_data35[3], in_dat_data35[4], in_dat_data35[5], in_dat_data35[6] };
  assign _08058_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *) { in_dat_data33[2], in_dat_data33[3], in_dat_data33[4], in_dat_data33[5], in_dat_data33[6] };
  assign _08059_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *) { in_dat_data31[2], in_dat_data31[3], in_dat_data31[4], in_dat_data31[5], in_dat_data31[6] };
  assign _08060_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *) { in_dat_data29[2], in_dat_data29[3], in_dat_data29[4], in_dat_data29[5], in_dat_data29[6] };
  assign _08061_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *) { in_dat_data27[2], in_dat_data27[3], in_dat_data27[4], in_dat_data27[5], in_dat_data27[6] };
  assign _08062_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *) { in_dat_data25[2], in_dat_data25[3], in_dat_data25[4], in_dat_data25[5], in_dat_data25[6] };
  assign _08063_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *) { in_dat_data23[2], in_dat_data23[3], in_dat_data23[4], in_dat_data23[5], in_dat_data23[6] };
  assign _08064_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *) { in_dat_data21[2], in_dat_data21[3], in_dat_data21[4], in_dat_data21[5], in_dat_data21[6] };
  assign _08065_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *) { in_dat_data19[2], in_dat_data19[3], in_dat_data19[4], in_dat_data19[5], in_dat_data19[6] };
  assign _08066_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *) { in_dat_data17[2], in_dat_data17[3], in_dat_data17[4], in_dat_data17[5], in_dat_data17[6] };
  assign _08067_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *) { in_dat_data15[2], in_dat_data15[3], in_dat_data15[4], in_dat_data15[5], in_dat_data15[6] };
  assign _08068_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *) { in_dat_data13[2], in_dat_data13[3], in_dat_data13[4], in_dat_data13[5], in_dat_data13[6] };
  assign _08069_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *) { in_dat_data11[2], in_dat_data11[3], in_dat_data11[4], in_dat_data11[5], in_dat_data11[6] };
  assign _08070_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *) { in_dat_data9[2], in_dat_data9[3], in_dat_data9[4], in_dat_data9[5], in_dat_data9[6] };
  assign _08071_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *) { in_dat_data7[2], in_dat_data7[3], in_dat_data7[4], in_dat_data7[5], in_dat_data7[6] };
  assign _08072_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *) { in_dat_data5[2], in_dat_data5[3], in_dat_data5[4], in_dat_data5[5], in_dat_data5[6] };
  assign _08073_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *) { in_dat_data3[2], in_dat_data3[3], in_dat_data3[4], in_dat_data3[5], in_dat_data3[6] };
  assign _08074_ = & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *) { in_dat_data1[2], in_dat_data1[3], in_dat_data1[4], in_dat_data1[5], in_dat_data1[6] };
  assign _08075_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2588" *) { in_wt_data126[0], in_wt_data126[1], in_wt_data126[2], in_wt_data126[3], in_wt_data126[4], in_wt_data126[5], in_wt_data126[6], in_wt_data126[7], in_wt_data127[0], in_wt_data127[1] };
  assign _08076_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2589" *) { in_wt_data124[0], in_wt_data124[1], in_wt_data124[2], in_wt_data124[3], in_wt_data124[4], in_wt_data124[5], in_wt_data124[6], in_wt_data124[7], in_wt_data125[0], in_wt_data125[1] };
  assign _08077_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2590" *) { in_wt_data122[0], in_wt_data122[1], in_wt_data122[2], in_wt_data122[3], in_wt_data122[4], in_wt_data122[5], in_wt_data122[6], in_wt_data122[7], in_wt_data123[0], in_wt_data123[1] };
  assign _08078_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2591" *) { in_wt_data120[0], in_wt_data120[1], in_wt_data120[2], in_wt_data120[3], in_wt_data120[4], in_wt_data120[5], in_wt_data120[6], in_wt_data120[7], in_wt_data121[0], in_wt_data121[1] };
  assign _08079_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2592" *) { in_wt_data118[0], in_wt_data118[1], in_wt_data118[2], in_wt_data118[3], in_wt_data118[4], in_wt_data118[5], in_wt_data118[6], in_wt_data118[7], in_wt_data119[0], in_wt_data119[1] };
  assign _08080_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2593" *) { in_wt_data116[0], in_wt_data116[1], in_wt_data116[2], in_wt_data116[3], in_wt_data116[4], in_wt_data116[5], in_wt_data116[6], in_wt_data116[7], in_wt_data117[0], in_wt_data117[1] };
  assign _08081_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2594" *) { in_wt_data114[0], in_wt_data114[1], in_wt_data114[2], in_wt_data114[3], in_wt_data114[4], in_wt_data114[5], in_wt_data114[6], in_wt_data114[7], in_wt_data115[0], in_wt_data115[1] };
  assign _08082_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2595" *) { in_wt_data112[0], in_wt_data112[1], in_wt_data112[2], in_wt_data112[3], in_wt_data112[4], in_wt_data112[5], in_wt_data112[6], in_wt_data112[7], in_wt_data113[0], in_wt_data113[1] };
  assign _08083_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2596" *) { in_wt_data110[0], in_wt_data110[1], in_wt_data110[2], in_wt_data110[3], in_wt_data110[4], in_wt_data110[5], in_wt_data110[6], in_wt_data110[7], in_wt_data111[0], in_wt_data111[1] };
  assign _08084_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2597" *) { in_wt_data108[0], in_wt_data108[1], in_wt_data108[2], in_wt_data108[3], in_wt_data108[4], in_wt_data108[5], in_wt_data108[6], in_wt_data108[7], in_wt_data109[0], in_wt_data109[1] };
  assign _08085_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2598" *) { in_wt_data106[0], in_wt_data106[1], in_wt_data106[2], in_wt_data106[3], in_wt_data106[4], in_wt_data106[5], in_wt_data106[6], in_wt_data106[7], in_wt_data107[0], in_wt_data107[1] };
  assign _08086_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2599" *) { in_wt_data104[0], in_wt_data104[1], in_wt_data104[2], in_wt_data104[3], in_wt_data104[4], in_wt_data104[5], in_wt_data104[6], in_wt_data104[7], in_wt_data105[0], in_wt_data105[1] };
  assign _08087_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2600" *) { in_wt_data102[0], in_wt_data102[1], in_wt_data102[2], in_wt_data102[3], in_wt_data102[4], in_wt_data102[5], in_wt_data102[6], in_wt_data102[7], in_wt_data103[0], in_wt_data103[1] };
  assign _08088_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2601" *) { in_wt_data100[0], in_wt_data100[1], in_wt_data100[2], in_wt_data100[3], in_wt_data100[4], in_wt_data100[5], in_wt_data100[6], in_wt_data100[7], in_wt_data101[0], in_wt_data101[1] };
  assign _08089_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2602" *) { in_wt_data98[0], in_wt_data98[1], in_wt_data98[2], in_wt_data98[3], in_wt_data98[4], in_wt_data98[5], in_wt_data98[6], in_wt_data98[7], in_wt_data99[0], in_wt_data99[1] };
  assign _08090_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2603" *) { in_wt_data96[0], in_wt_data96[1], in_wt_data96[2], in_wt_data96[3], in_wt_data96[4], in_wt_data96[5], in_wt_data96[6], in_wt_data96[7], in_wt_data97[0], in_wt_data97[1] };
  assign _08091_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2604" *) { in_wt_data94[0], in_wt_data94[1], in_wt_data94[2], in_wt_data94[3], in_wt_data94[4], in_wt_data94[5], in_wt_data94[6], in_wt_data94[7], in_wt_data95[0], in_wt_data95[1] };
  assign _08092_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2605" *) { in_wt_data92[0], in_wt_data92[1], in_wt_data92[2], in_wt_data92[3], in_wt_data92[4], in_wt_data92[5], in_wt_data92[6], in_wt_data92[7], in_wt_data93[0], in_wt_data93[1] };
  assign _08093_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2606" *) { in_wt_data90[0], in_wt_data90[1], in_wt_data90[2], in_wt_data90[3], in_wt_data90[4], in_wt_data90[5], in_wt_data90[6], in_wt_data90[7], in_wt_data91[0], in_wt_data91[1] };
  assign _08094_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2607" *) { in_wt_data88[0], in_wt_data88[1], in_wt_data88[2], in_wt_data88[3], in_wt_data88[4], in_wt_data88[5], in_wt_data88[6], in_wt_data88[7], in_wt_data89[0], in_wt_data89[1] };
  assign _08095_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2608" *) { in_wt_data86[0], in_wt_data86[1], in_wt_data86[2], in_wt_data86[3], in_wt_data86[4], in_wt_data86[5], in_wt_data86[6], in_wt_data86[7], in_wt_data87[0], in_wt_data87[1] };
  assign _08096_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2609" *) { in_wt_data84[0], in_wt_data84[1], in_wt_data84[2], in_wt_data84[3], in_wt_data84[4], in_wt_data84[5], in_wt_data84[6], in_wt_data84[7], in_wt_data85[0], in_wt_data85[1] };
  assign _08097_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2610" *) { in_wt_data82[0], in_wt_data82[1], in_wt_data82[2], in_wt_data82[3], in_wt_data82[4], in_wt_data82[5], in_wt_data82[6], in_wt_data82[7], in_wt_data83[0], in_wt_data83[1] };
  assign _08098_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2611" *) { in_wt_data80[0], in_wt_data80[1], in_wt_data80[2], in_wt_data80[3], in_wt_data80[4], in_wt_data80[5], in_wt_data80[6], in_wt_data80[7], in_wt_data81[0], in_wt_data81[1] };
  assign _08099_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2612" *) { in_wt_data78[0], in_wt_data78[1], in_wt_data78[2], in_wt_data78[3], in_wt_data78[4], in_wt_data78[5], in_wt_data78[6], in_wt_data78[7], in_wt_data79[0], in_wt_data79[1] };
  assign _08100_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2613" *) { in_wt_data76[0], in_wt_data76[1], in_wt_data76[2], in_wt_data76[3], in_wt_data76[4], in_wt_data76[5], in_wt_data76[6], in_wt_data76[7], in_wt_data77[0], in_wt_data77[1] };
  assign _08101_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2614" *) { in_wt_data74[0], in_wt_data74[1], in_wt_data74[2], in_wt_data74[3], in_wt_data74[4], in_wt_data74[5], in_wt_data74[6], in_wt_data74[7], in_wt_data75[0], in_wt_data75[1] };
  assign _08102_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2615" *) { in_wt_data72[0], in_wt_data72[1], in_wt_data72[2], in_wt_data72[3], in_wt_data72[4], in_wt_data72[5], in_wt_data72[6], in_wt_data72[7], in_wt_data73[0], in_wt_data73[1] };
  assign _08103_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2616" *) { in_wt_data70[0], in_wt_data70[1], in_wt_data70[2], in_wt_data70[3], in_wt_data70[4], in_wt_data70[5], in_wt_data70[6], in_wt_data70[7], in_wt_data71[0], in_wt_data71[1] };
  assign _08104_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2617" *) { in_wt_data68[0], in_wt_data68[1], in_wt_data68[2], in_wt_data68[3], in_wt_data68[4], in_wt_data68[5], in_wt_data68[6], in_wt_data68[7], in_wt_data69[0], in_wt_data69[1] };
  assign _08105_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2618" *) { in_wt_data66[0], in_wt_data66[1], in_wt_data66[2], in_wt_data66[3], in_wt_data66[4], in_wt_data66[5], in_wt_data66[6], in_wt_data66[7], in_wt_data67[0], in_wt_data67[1] };
  assign _08106_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2619" *) { in_wt_data64[0], in_wt_data64[1], in_wt_data64[2], in_wt_data64[3], in_wt_data64[4], in_wt_data64[5], in_wt_data64[6], in_wt_data64[7], in_wt_data65[0], in_wt_data65[1] };
  assign _08107_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2620" *) { in_wt_data62[0], in_wt_data62[1], in_wt_data62[2], in_wt_data62[3], in_wt_data62[4], in_wt_data62[5], in_wt_data62[6], in_wt_data62[7], in_wt_data63[0], in_wt_data63[1] };
  assign _08108_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2621" *) { in_wt_data60[0], in_wt_data60[1], in_wt_data60[2], in_wt_data60[3], in_wt_data60[4], in_wt_data60[5], in_wt_data60[6], in_wt_data60[7], in_wt_data61[0], in_wt_data61[1] };
  assign _08109_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2622" *) { in_wt_data58[0], in_wt_data58[1], in_wt_data58[2], in_wt_data58[3], in_wt_data58[4], in_wt_data58[5], in_wt_data58[6], in_wt_data58[7], in_wt_data59[0], in_wt_data59[1] };
  assign _08110_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2623" *) { in_wt_data56[0], in_wt_data56[1], in_wt_data56[2], in_wt_data56[3], in_wt_data56[4], in_wt_data56[5], in_wt_data56[6], in_wt_data56[7], in_wt_data57[0], in_wt_data57[1] };
  assign _08111_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2624" *) { in_wt_data54[0], in_wt_data54[1], in_wt_data54[2], in_wt_data54[3], in_wt_data54[4], in_wt_data54[5], in_wt_data54[6], in_wt_data54[7], in_wt_data55[0], in_wt_data55[1] };
  assign _08112_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2625" *) { in_wt_data52[0], in_wt_data52[1], in_wt_data52[2], in_wt_data52[3], in_wt_data52[4], in_wt_data52[5], in_wt_data52[6], in_wt_data52[7], in_wt_data53[0], in_wt_data53[1] };
  assign _08113_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2626" *) { in_wt_data50[0], in_wt_data50[1], in_wt_data50[2], in_wt_data50[3], in_wt_data50[4], in_wt_data50[5], in_wt_data50[6], in_wt_data50[7], in_wt_data51[0], in_wt_data51[1] };
  assign _08114_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2627" *) { in_wt_data48[0], in_wt_data48[1], in_wt_data48[2], in_wt_data48[3], in_wt_data48[4], in_wt_data48[5], in_wt_data48[6], in_wt_data48[7], in_wt_data49[0], in_wt_data49[1] };
  assign _08115_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2628" *) { in_wt_data46[0], in_wt_data46[1], in_wt_data46[2], in_wt_data46[3], in_wt_data46[4], in_wt_data46[5], in_wt_data46[6], in_wt_data46[7], in_wt_data47[0], in_wt_data47[1] };
  assign _08116_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2629" *) { in_wt_data44[0], in_wt_data44[1], in_wt_data44[2], in_wt_data44[3], in_wt_data44[4], in_wt_data44[5], in_wt_data44[6], in_wt_data44[7], in_wt_data45[0], in_wt_data45[1] };
  assign _08117_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2630" *) { in_wt_data42[0], in_wt_data42[1], in_wt_data42[2], in_wt_data42[3], in_wt_data42[4], in_wt_data42[5], in_wt_data42[6], in_wt_data42[7], in_wt_data43[0], in_wt_data43[1] };
  assign _08118_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2631" *) { in_wt_data40[0], in_wt_data40[1], in_wt_data40[2], in_wt_data40[3], in_wt_data40[4], in_wt_data40[5], in_wt_data40[6], in_wt_data40[7], in_wt_data41[0], in_wt_data41[1] };
  assign _08119_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2632" *) { in_wt_data38[0], in_wt_data38[1], in_wt_data38[2], in_wt_data38[3], in_wt_data38[4], in_wt_data38[5], in_wt_data38[6], in_wt_data38[7], in_wt_data39[0], in_wt_data39[1] };
  assign _08120_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2633" *) { in_wt_data36[0], in_wt_data36[1], in_wt_data36[2], in_wt_data36[3], in_wt_data36[4], in_wt_data36[5], in_wt_data36[6], in_wt_data36[7], in_wt_data37[0], in_wt_data37[1] };
  assign _08121_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2634" *) { in_wt_data34[0], in_wt_data34[1], in_wt_data34[2], in_wt_data34[3], in_wt_data34[4], in_wt_data34[5], in_wt_data34[6], in_wt_data34[7], in_wt_data35[0], in_wt_data35[1] };
  assign _08122_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2635" *) { in_wt_data32[0], in_wt_data32[1], in_wt_data32[2], in_wt_data32[3], in_wt_data32[4], in_wt_data32[5], in_wt_data32[6], in_wt_data32[7], in_wt_data33[0], in_wt_data33[1] };
  assign _08123_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2636" *) { in_wt_data30[0], in_wt_data30[1], in_wt_data30[2], in_wt_data30[3], in_wt_data30[4], in_wt_data30[5], in_wt_data30[6], in_wt_data30[7], in_wt_data31[0], in_wt_data31[1] };
  assign _08124_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2637" *) { in_wt_data28[0], in_wt_data28[1], in_wt_data28[2], in_wt_data28[3], in_wt_data28[4], in_wt_data28[5], in_wt_data28[6], in_wt_data28[7], in_wt_data29[0], in_wt_data29[1] };
  assign _08125_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2638" *) { in_wt_data26[0], in_wt_data26[1], in_wt_data26[2], in_wt_data26[3], in_wt_data26[4], in_wt_data26[5], in_wt_data26[6], in_wt_data26[7], in_wt_data27[0], in_wt_data27[1] };
  assign _08126_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2639" *) { in_wt_data24[0], in_wt_data24[1], in_wt_data24[2], in_wt_data24[3], in_wt_data24[4], in_wt_data24[5], in_wt_data24[6], in_wt_data24[7], in_wt_data25[0], in_wt_data25[1] };
  assign _08127_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2640" *) { in_wt_data22[0], in_wt_data22[1], in_wt_data22[2], in_wt_data22[3], in_wt_data22[4], in_wt_data22[5], in_wt_data22[6], in_wt_data22[7], in_wt_data23[0], in_wt_data23[1] };
  assign _08128_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2641" *) { in_wt_data20[0], in_wt_data20[1], in_wt_data20[2], in_wt_data20[3], in_wt_data20[4], in_wt_data20[5], in_wt_data20[6], in_wt_data20[7], in_wt_data21[0], in_wt_data21[1] };
  assign _08129_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2642" *) { in_wt_data18[0], in_wt_data18[1], in_wt_data18[2], in_wt_data18[3], in_wt_data18[4], in_wt_data18[5], in_wt_data18[6], in_wt_data18[7], in_wt_data19[0], in_wt_data19[1] };
  assign _08130_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2643" *) { in_wt_data16[0], in_wt_data16[1], in_wt_data16[2], in_wt_data16[3], in_wt_data16[4], in_wt_data16[5], in_wt_data16[6], in_wt_data16[7], in_wt_data17[0], in_wt_data17[1] };
  assign _08131_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2644" *) { in_wt_data14[0], in_wt_data14[1], in_wt_data14[2], in_wt_data14[3], in_wt_data14[4], in_wt_data14[5], in_wt_data14[6], in_wt_data14[7], in_wt_data15[0], in_wt_data15[1] };
  assign _08132_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2645" *) { in_wt_data12[0], in_wt_data12[1], in_wt_data12[2], in_wt_data12[3], in_wt_data12[4], in_wt_data12[5], in_wt_data12[6], in_wt_data12[7], in_wt_data13[0], in_wt_data13[1] };
  assign _08133_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2646" *) { in_wt_data10[0], in_wt_data10[1], in_wt_data10[2], in_wt_data10[3], in_wt_data10[4], in_wt_data10[5], in_wt_data10[6], in_wt_data10[7], in_wt_data11[0], in_wt_data11[1] };
  assign _08134_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2647" *) { in_wt_data8[0], in_wt_data8[1], in_wt_data8[2], in_wt_data8[3], in_wt_data8[4], in_wt_data8[5], in_wt_data8[6], in_wt_data8[7], in_wt_data9[0], in_wt_data9[1] };
  assign _08135_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2648" *) { in_wt_data6[0], in_wt_data6[1], in_wt_data6[2], in_wt_data6[3], in_wt_data6[4], in_wt_data6[5], in_wt_data6[6], in_wt_data6[7], in_wt_data7[0], in_wt_data7[1] };
  assign _08136_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2649" *) { in_wt_data4[0], in_wt_data4[1], in_wt_data4[2], in_wt_data4[3], in_wt_data4[4], in_wt_data4[5], in_wt_data4[6], in_wt_data4[7], in_wt_data5[0], in_wt_data5[1] };
  assign _08137_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2650" *) { in_wt_data2[0], in_wt_data2[1], in_wt_data2[2], in_wt_data2[3], in_wt_data2[4], in_wt_data2[5], in_wt_data2[6], in_wt_data2[7], in_wt_data3[0], in_wt_data3[1] };
  assign _08138_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2651" *) { in_wt_data0[0], in_wt_data0[1], in_wt_data0[2], in_wt_data0[3], in_wt_data0[4], in_wt_data0[5], in_wt_data0[6], in_wt_data0[7], in_wt_data1[0], in_wt_data1[1] };
  assign _08139_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2727" *) { in_wt_data127[2], in_wt_data127[3], in_wt_data127[4], in_wt_data127[5], in_wt_data127[6] };
  assign _08140_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2728" *) { in_wt_data125[2], in_wt_data125[3], in_wt_data125[4], in_wt_data125[5], in_wt_data125[6] };
  assign _08141_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2729" *) { in_wt_data123[2], in_wt_data123[3], in_wt_data123[4], in_wt_data123[5], in_wt_data123[6] };
  assign _08142_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2730" *) { in_wt_data121[2], in_wt_data121[3], in_wt_data121[4], in_wt_data121[5], in_wt_data121[6] };
  assign _08143_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2731" *) { in_wt_data119[2], in_wt_data119[3], in_wt_data119[4], in_wt_data119[5], in_wt_data119[6] };
  assign _08144_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2732" *) { in_wt_data117[2], in_wt_data117[3], in_wt_data117[4], in_wt_data117[5], in_wt_data117[6] };
  assign _08145_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2733" *) { in_wt_data115[2], in_wt_data115[3], in_wt_data115[4], in_wt_data115[5], in_wt_data115[6] };
  assign _08146_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2734" *) { in_wt_data113[2], in_wt_data113[3], in_wt_data113[4], in_wt_data113[5], in_wt_data113[6] };
  assign _08147_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2735" *) { in_wt_data111[2], in_wt_data111[3], in_wt_data111[4], in_wt_data111[5], in_wt_data111[6] };
  assign _08148_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2736" *) { in_wt_data109[2], in_wt_data109[3], in_wt_data109[4], in_wt_data109[5], in_wt_data109[6] };
  assign _08149_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2737" *) { in_wt_data107[2], in_wt_data107[3], in_wt_data107[4], in_wt_data107[5], in_wt_data107[6] };
  assign _08150_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2738" *) { in_wt_data105[2], in_wt_data105[3], in_wt_data105[4], in_wt_data105[5], in_wt_data105[6] };
  assign _08151_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2739" *) { in_wt_data103[2], in_wt_data103[3], in_wt_data103[4], in_wt_data103[5], in_wt_data103[6] };
  assign _08152_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2740" *) { in_wt_data101[2], in_wt_data101[3], in_wt_data101[4], in_wt_data101[5], in_wt_data101[6] };
  assign _08153_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2741" *) { in_wt_data99[2], in_wt_data99[3], in_wt_data99[4], in_wt_data99[5], in_wt_data99[6] };
  assign _08154_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2742" *) { in_wt_data97[2], in_wt_data97[3], in_wt_data97[4], in_wt_data97[5], in_wt_data97[6] };
  assign _08155_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2743" *) { in_wt_data95[2], in_wt_data95[3], in_wt_data95[4], in_wt_data95[5], in_wt_data95[6] };
  assign _08156_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2744" *) { in_wt_data93[2], in_wt_data93[3], in_wt_data93[4], in_wt_data93[5], in_wt_data93[6] };
  assign _08157_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2745" *) { in_wt_data91[2], in_wt_data91[3], in_wt_data91[4], in_wt_data91[5], in_wt_data91[6] };
  assign _08158_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2746" *) { in_wt_data89[2], in_wt_data89[3], in_wt_data89[4], in_wt_data89[5], in_wt_data89[6] };
  assign _08159_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2747" *) { in_wt_data87[2], in_wt_data87[3], in_wt_data87[4], in_wt_data87[5], in_wt_data87[6] };
  assign _08160_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2748" *) { in_wt_data85[2], in_wt_data85[3], in_wt_data85[4], in_wt_data85[5], in_wt_data85[6] };
  assign _08161_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2749" *) { in_wt_data83[2], in_wt_data83[3], in_wt_data83[4], in_wt_data83[5], in_wt_data83[6] };
  assign _08162_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2750" *) { in_wt_data81[2], in_wt_data81[3], in_wt_data81[4], in_wt_data81[5], in_wt_data81[6] };
  assign _08163_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2751" *) { in_wt_data79[2], in_wt_data79[3], in_wt_data79[4], in_wt_data79[5], in_wt_data79[6] };
  assign _08164_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2752" *) { in_wt_data77[2], in_wt_data77[3], in_wt_data77[4], in_wt_data77[5], in_wt_data77[6] };
  assign _08165_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2753" *) { in_wt_data75[2], in_wt_data75[3], in_wt_data75[4], in_wt_data75[5], in_wt_data75[6] };
  assign _08166_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2754" *) { in_wt_data73[2], in_wt_data73[3], in_wt_data73[4], in_wt_data73[5], in_wt_data73[6] };
  assign _08167_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2755" *) { in_wt_data71[2], in_wt_data71[3], in_wt_data71[4], in_wt_data71[5], in_wt_data71[6] };
  assign _08168_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2756" *) { in_wt_data69[2], in_wt_data69[3], in_wt_data69[4], in_wt_data69[5], in_wt_data69[6] };
  assign _08169_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2757" *) { in_wt_data67[2], in_wt_data67[3], in_wt_data67[4], in_wt_data67[5], in_wt_data67[6] };
  assign _08170_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2758" *) { in_wt_data65[2], in_wt_data65[3], in_wt_data65[4], in_wt_data65[5], in_wt_data65[6] };
  assign _08171_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2759" *) { in_wt_data63[2], in_wt_data63[3], in_wt_data63[4], in_wt_data63[5], in_wt_data63[6] };
  assign _08172_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2760" *) { in_wt_data61[2], in_wt_data61[3], in_wt_data61[4], in_wt_data61[5], in_wt_data61[6] };
  assign _08173_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2761" *) { in_wt_data59[2], in_wt_data59[3], in_wt_data59[4], in_wt_data59[5], in_wt_data59[6] };
  assign _08174_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2762" *) { in_wt_data57[2], in_wt_data57[3], in_wt_data57[4], in_wt_data57[5], in_wt_data57[6] };
  assign _08175_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2763" *) { in_wt_data55[2], in_wt_data55[3], in_wt_data55[4], in_wt_data55[5], in_wt_data55[6] };
  assign _08176_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2764" *) { in_wt_data53[2], in_wt_data53[3], in_wt_data53[4], in_wt_data53[5], in_wt_data53[6] };
  assign _08177_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2765" *) { in_wt_data51[2], in_wt_data51[3], in_wt_data51[4], in_wt_data51[5], in_wt_data51[6] };
  assign _08178_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2766" *) { in_wt_data49[2], in_wt_data49[3], in_wt_data49[4], in_wt_data49[5], in_wt_data49[6] };
  assign _08179_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27661" *) { in_dat_data126[0], in_dat_data126[1], in_dat_data126[2], in_dat_data126[3], in_dat_data126[4], in_dat_data126[5], in_dat_data126[6], in_dat_data126[7], in_dat_data127[0], in_dat_data127[1] };
  assign _08180_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27662" *) { in_dat_data124[0], in_dat_data124[1], in_dat_data124[2], in_dat_data124[3], in_dat_data124[4], in_dat_data124[5], in_dat_data124[6], in_dat_data124[7], in_dat_data125[0], in_dat_data125[1] };
  assign _08181_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27663" *) { in_dat_data122[0], in_dat_data122[1], in_dat_data122[2], in_dat_data122[3], in_dat_data122[4], in_dat_data122[5], in_dat_data122[6], in_dat_data122[7], in_dat_data123[0], in_dat_data123[1] };
  assign _08182_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27664" *) { in_dat_data120[0], in_dat_data120[1], in_dat_data120[2], in_dat_data120[3], in_dat_data120[4], in_dat_data120[5], in_dat_data120[6], in_dat_data120[7], in_dat_data121[0], in_dat_data121[1] };
  assign _08183_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27665" *) { in_dat_data118[0], in_dat_data118[1], in_dat_data118[2], in_dat_data118[3], in_dat_data118[4], in_dat_data118[5], in_dat_data118[6], in_dat_data118[7], in_dat_data119[0], in_dat_data119[1] };
  assign _08184_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27666" *) { in_dat_data116[0], in_dat_data116[1], in_dat_data116[2], in_dat_data116[3], in_dat_data116[4], in_dat_data116[5], in_dat_data116[6], in_dat_data116[7], in_dat_data117[0], in_dat_data117[1] };
  assign _08185_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27667" *) { in_dat_data114[0], in_dat_data114[1], in_dat_data114[2], in_dat_data114[3], in_dat_data114[4], in_dat_data114[5], in_dat_data114[6], in_dat_data114[7], in_dat_data115[0], in_dat_data115[1] };
  assign _08186_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27668" *) { in_dat_data112[0], in_dat_data112[1], in_dat_data112[2], in_dat_data112[3], in_dat_data112[4], in_dat_data112[5], in_dat_data112[6], in_dat_data112[7], in_dat_data113[0], in_dat_data113[1] };
  assign _08187_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27669" *) { in_dat_data110[0], in_dat_data110[1], in_dat_data110[2], in_dat_data110[3], in_dat_data110[4], in_dat_data110[5], in_dat_data110[6], in_dat_data110[7], in_dat_data111[0], in_dat_data111[1] };
  assign _08188_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2767" *) { in_wt_data47[2], in_wt_data47[3], in_wt_data47[4], in_wt_data47[5], in_wt_data47[6] };
  assign _08189_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27670" *) { in_dat_data108[0], in_dat_data108[1], in_dat_data108[2], in_dat_data108[3], in_dat_data108[4], in_dat_data108[5], in_dat_data108[6], in_dat_data108[7], in_dat_data109[0], in_dat_data109[1] };
  assign _08190_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27671" *) { in_dat_data106[0], in_dat_data106[1], in_dat_data106[2], in_dat_data106[3], in_dat_data106[4], in_dat_data106[5], in_dat_data106[6], in_dat_data106[7], in_dat_data107[0], in_dat_data107[1] };
  assign _08191_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27672" *) { in_dat_data104[0], in_dat_data104[1], in_dat_data104[2], in_dat_data104[3], in_dat_data104[4], in_dat_data104[5], in_dat_data104[6], in_dat_data104[7], in_dat_data105[0], in_dat_data105[1] };
  assign _08192_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27673" *) { in_dat_data102[0], in_dat_data102[1], in_dat_data102[2], in_dat_data102[3], in_dat_data102[4], in_dat_data102[5], in_dat_data102[6], in_dat_data102[7], in_dat_data103[0], in_dat_data103[1] };
  assign _08193_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27674" *) { in_dat_data100[0], in_dat_data100[1], in_dat_data100[2], in_dat_data100[3], in_dat_data100[4], in_dat_data100[5], in_dat_data100[6], in_dat_data100[7], in_dat_data101[0], in_dat_data101[1] };
  assign _08194_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27675" *) { in_dat_data98[0], in_dat_data98[1], in_dat_data98[2], in_dat_data98[3], in_dat_data98[4], in_dat_data98[5], in_dat_data98[6], in_dat_data98[7], in_dat_data99[0], in_dat_data99[1] };
  assign _08195_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27676" *) { in_dat_data96[0], in_dat_data96[1], in_dat_data96[2], in_dat_data96[3], in_dat_data96[4], in_dat_data96[5], in_dat_data96[6], in_dat_data96[7], in_dat_data97[0], in_dat_data97[1] };
  assign _08196_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27677" *) { in_dat_data94[0], in_dat_data94[1], in_dat_data94[2], in_dat_data94[3], in_dat_data94[4], in_dat_data94[5], in_dat_data94[6], in_dat_data94[7], in_dat_data95[0], in_dat_data95[1] };
  assign _08197_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27678" *) { in_dat_data92[0], in_dat_data92[1], in_dat_data92[2], in_dat_data92[3], in_dat_data92[4], in_dat_data92[5], in_dat_data92[6], in_dat_data92[7], in_dat_data93[0], in_dat_data93[1] };
  assign _08198_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27679" *) { in_dat_data90[0], in_dat_data90[1], in_dat_data90[2], in_dat_data90[3], in_dat_data90[4], in_dat_data90[5], in_dat_data90[6], in_dat_data90[7], in_dat_data91[0], in_dat_data91[1] };
  assign _08199_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2768" *) { in_wt_data45[2], in_wt_data45[3], in_wt_data45[4], in_wt_data45[5], in_wt_data45[6] };
  assign _08200_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27680" *) { in_dat_data88[0], in_dat_data88[1], in_dat_data88[2], in_dat_data88[3], in_dat_data88[4], in_dat_data88[5], in_dat_data88[6], in_dat_data88[7], in_dat_data89[0], in_dat_data89[1] };
  assign _08201_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27681" *) { in_dat_data86[0], in_dat_data86[1], in_dat_data86[2], in_dat_data86[3], in_dat_data86[4], in_dat_data86[5], in_dat_data86[6], in_dat_data86[7], in_dat_data87[0], in_dat_data87[1] };
  assign _08202_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27682" *) { in_dat_data84[0], in_dat_data84[1], in_dat_data84[2], in_dat_data84[3], in_dat_data84[4], in_dat_data84[5], in_dat_data84[6], in_dat_data84[7], in_dat_data85[0], in_dat_data85[1] };
  assign _08203_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27683" *) { in_dat_data82[0], in_dat_data82[1], in_dat_data82[2], in_dat_data82[3], in_dat_data82[4], in_dat_data82[5], in_dat_data82[6], in_dat_data82[7], in_dat_data83[0], in_dat_data83[1] };
  assign _08204_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27684" *) { in_dat_data80[0], in_dat_data80[1], in_dat_data80[2], in_dat_data80[3], in_dat_data80[4], in_dat_data80[5], in_dat_data80[6], in_dat_data80[7], in_dat_data81[0], in_dat_data81[1] };
  assign _08205_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27685" *) { in_dat_data78[0], in_dat_data78[1], in_dat_data78[2], in_dat_data78[3], in_dat_data78[4], in_dat_data78[5], in_dat_data78[6], in_dat_data78[7], in_dat_data79[0], in_dat_data79[1] };
  assign _08206_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27686" *) { in_dat_data76[0], in_dat_data76[1], in_dat_data76[2], in_dat_data76[3], in_dat_data76[4], in_dat_data76[5], in_dat_data76[6], in_dat_data76[7], in_dat_data77[0], in_dat_data77[1] };
  assign _08207_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27687" *) { in_dat_data74[0], in_dat_data74[1], in_dat_data74[2], in_dat_data74[3], in_dat_data74[4], in_dat_data74[5], in_dat_data74[6], in_dat_data74[7], in_dat_data75[0], in_dat_data75[1] };
  assign _08208_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27688" *) { in_dat_data72[0], in_dat_data72[1], in_dat_data72[2], in_dat_data72[3], in_dat_data72[4], in_dat_data72[5], in_dat_data72[6], in_dat_data72[7], in_dat_data73[0], in_dat_data73[1] };
  assign _08209_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27689" *) { in_dat_data70[0], in_dat_data70[1], in_dat_data70[2], in_dat_data70[3], in_dat_data70[4], in_dat_data70[5], in_dat_data70[6], in_dat_data70[7], in_dat_data71[0], in_dat_data71[1] };
  assign _08210_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2769" *) { in_wt_data43[2], in_wt_data43[3], in_wt_data43[4], in_wt_data43[5], in_wt_data43[6] };
  assign _08211_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27690" *) { in_dat_data68[0], in_dat_data68[1], in_dat_data68[2], in_dat_data68[3], in_dat_data68[4], in_dat_data68[5], in_dat_data68[6], in_dat_data68[7], in_dat_data69[0], in_dat_data69[1] };
  assign _08212_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27691" *) { in_dat_data66[0], in_dat_data66[1], in_dat_data66[2], in_dat_data66[3], in_dat_data66[4], in_dat_data66[5], in_dat_data66[6], in_dat_data66[7], in_dat_data67[0], in_dat_data67[1] };
  assign _08213_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27692" *) { in_dat_data64[0], in_dat_data64[1], in_dat_data64[2], in_dat_data64[3], in_dat_data64[4], in_dat_data64[5], in_dat_data64[6], in_dat_data64[7], in_dat_data65[0], in_dat_data65[1] };
  assign _08214_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27693" *) { in_dat_data62[0], in_dat_data62[1], in_dat_data62[2], in_dat_data62[3], in_dat_data62[4], in_dat_data62[5], in_dat_data62[6], in_dat_data62[7], in_dat_data63[0], in_dat_data63[1] };
  assign _08215_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27694" *) { in_dat_data60[0], in_dat_data60[1], in_dat_data60[2], in_dat_data60[3], in_dat_data60[4], in_dat_data60[5], in_dat_data60[6], in_dat_data60[7], in_dat_data61[0], in_dat_data61[1] };
  assign _08216_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27695" *) { in_dat_data58[0], in_dat_data58[1], in_dat_data58[2], in_dat_data58[3], in_dat_data58[4], in_dat_data58[5], in_dat_data58[6], in_dat_data58[7], in_dat_data59[0], in_dat_data59[1] };
  assign _08217_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27696" *) { in_dat_data56[0], in_dat_data56[1], in_dat_data56[2], in_dat_data56[3], in_dat_data56[4], in_dat_data56[5], in_dat_data56[6], in_dat_data56[7], in_dat_data57[0], in_dat_data57[1] };
  assign _08218_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27697" *) { in_dat_data54[0], in_dat_data54[1], in_dat_data54[2], in_dat_data54[3], in_dat_data54[4], in_dat_data54[5], in_dat_data54[6], in_dat_data54[7], in_dat_data55[0], in_dat_data55[1] };
  assign _08219_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27698" *) { in_dat_data52[0], in_dat_data52[1], in_dat_data52[2], in_dat_data52[3], in_dat_data52[4], in_dat_data52[5], in_dat_data52[6], in_dat_data52[7], in_dat_data53[0], in_dat_data53[1] };
  assign _08220_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27699" *) { in_dat_data50[0], in_dat_data50[1], in_dat_data50[2], in_dat_data50[3], in_dat_data50[4], in_dat_data50[5], in_dat_data50[6], in_dat_data50[7], in_dat_data51[0], in_dat_data51[1] };
  assign _08221_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2770" *) { in_wt_data41[2], in_wt_data41[3], in_wt_data41[4], in_wt_data41[5], in_wt_data41[6] };
  assign _08222_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27700" *) { in_dat_data48[0], in_dat_data48[1], in_dat_data48[2], in_dat_data48[3], in_dat_data48[4], in_dat_data48[5], in_dat_data48[6], in_dat_data48[7], in_dat_data49[0], in_dat_data49[1] };
  assign _08223_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27701" *) { in_dat_data46[0], in_dat_data46[1], in_dat_data46[2], in_dat_data46[3], in_dat_data46[4], in_dat_data46[5], in_dat_data46[6], in_dat_data46[7], in_dat_data47[0], in_dat_data47[1] };
  assign _08224_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27702" *) { in_dat_data44[0], in_dat_data44[1], in_dat_data44[2], in_dat_data44[3], in_dat_data44[4], in_dat_data44[5], in_dat_data44[6], in_dat_data44[7], in_dat_data45[0], in_dat_data45[1] };
  assign _08225_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27703" *) { in_dat_data42[0], in_dat_data42[1], in_dat_data42[2], in_dat_data42[3], in_dat_data42[4], in_dat_data42[5], in_dat_data42[6], in_dat_data42[7], in_dat_data43[0], in_dat_data43[1] };
  assign _08226_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27704" *) { in_dat_data40[0], in_dat_data40[1], in_dat_data40[2], in_dat_data40[3], in_dat_data40[4], in_dat_data40[5], in_dat_data40[6], in_dat_data40[7], in_dat_data41[0], in_dat_data41[1] };
  assign _08227_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27705" *) { in_dat_data38[0], in_dat_data38[1], in_dat_data38[2], in_dat_data38[3], in_dat_data38[4], in_dat_data38[5], in_dat_data38[6], in_dat_data38[7], in_dat_data39[0], in_dat_data39[1] };
  assign _08228_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27706" *) { in_dat_data36[0], in_dat_data36[1], in_dat_data36[2], in_dat_data36[3], in_dat_data36[4], in_dat_data36[5], in_dat_data36[6], in_dat_data36[7], in_dat_data37[0], in_dat_data37[1] };
  assign _08229_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27707" *) { in_dat_data34[0], in_dat_data34[1], in_dat_data34[2], in_dat_data34[3], in_dat_data34[4], in_dat_data34[5], in_dat_data34[6], in_dat_data34[7], in_dat_data35[0], in_dat_data35[1] };
  assign _08230_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27708" *) { in_dat_data32[0], in_dat_data32[1], in_dat_data32[2], in_dat_data32[3], in_dat_data32[4], in_dat_data32[5], in_dat_data32[6], in_dat_data32[7], in_dat_data33[0], in_dat_data33[1] };
  assign _08231_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27709" *) { in_dat_data30[0], in_dat_data30[1], in_dat_data30[2], in_dat_data30[3], in_dat_data30[4], in_dat_data30[5], in_dat_data30[6], in_dat_data30[7], in_dat_data31[0], in_dat_data31[1] };
  assign _08232_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2771" *) { in_wt_data39[2], in_wt_data39[3], in_wt_data39[4], in_wt_data39[5], in_wt_data39[6] };
  assign _08233_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27710" *) { in_dat_data28[0], in_dat_data28[1], in_dat_data28[2], in_dat_data28[3], in_dat_data28[4], in_dat_data28[5], in_dat_data28[6], in_dat_data28[7], in_dat_data29[0], in_dat_data29[1] };
  assign _08234_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27711" *) { in_dat_data26[0], in_dat_data26[1], in_dat_data26[2], in_dat_data26[3], in_dat_data26[4], in_dat_data26[5], in_dat_data26[6], in_dat_data26[7], in_dat_data27[0], in_dat_data27[1] };
  assign _08235_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27712" *) { in_dat_data24[0], in_dat_data24[1], in_dat_data24[2], in_dat_data24[3], in_dat_data24[4], in_dat_data24[5], in_dat_data24[6], in_dat_data24[7], in_dat_data25[0], in_dat_data25[1] };
  assign _08236_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27713" *) { in_dat_data22[0], in_dat_data22[1], in_dat_data22[2], in_dat_data22[3], in_dat_data22[4], in_dat_data22[5], in_dat_data22[6], in_dat_data22[7], in_dat_data23[0], in_dat_data23[1] };
  assign _08237_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27714" *) { in_dat_data20[0], in_dat_data20[1], in_dat_data20[2], in_dat_data20[3], in_dat_data20[4], in_dat_data20[5], in_dat_data20[6], in_dat_data20[7], in_dat_data21[0], in_dat_data21[1] };
  assign _08238_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27715" *) { in_dat_data18[0], in_dat_data18[1], in_dat_data18[2], in_dat_data18[3], in_dat_data18[4], in_dat_data18[5], in_dat_data18[6], in_dat_data18[7], in_dat_data19[0], in_dat_data19[1] };
  assign _08239_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27716" *) { in_dat_data16[0], in_dat_data16[1], in_dat_data16[2], in_dat_data16[3], in_dat_data16[4], in_dat_data16[5], in_dat_data16[6], in_dat_data16[7], in_dat_data17[0], in_dat_data17[1] };
  assign _08240_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27717" *) { in_dat_data14[0], in_dat_data14[1], in_dat_data14[2], in_dat_data14[3], in_dat_data14[4], in_dat_data14[5], in_dat_data14[6], in_dat_data14[7], in_dat_data15[0], in_dat_data15[1] };
  assign _08241_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27718" *) { in_dat_data12[0], in_dat_data12[1], in_dat_data12[2], in_dat_data12[3], in_dat_data12[4], in_dat_data12[5], in_dat_data12[6], in_dat_data12[7], in_dat_data13[0], in_dat_data13[1] };
  assign _08242_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27719" *) { in_dat_data10[0], in_dat_data10[1], in_dat_data10[2], in_dat_data10[3], in_dat_data10[4], in_dat_data10[5], in_dat_data10[6], in_dat_data10[7], in_dat_data11[0], in_dat_data11[1] };
  assign _08243_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2772" *) { in_wt_data37[2], in_wt_data37[3], in_wt_data37[4], in_wt_data37[5], in_wt_data37[6] };
  assign _08244_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27720" *) { in_dat_data8[0], in_dat_data8[1], in_dat_data8[2], in_dat_data8[3], in_dat_data8[4], in_dat_data8[5], in_dat_data8[6], in_dat_data8[7], in_dat_data9[0], in_dat_data9[1] };
  assign _08245_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27721" *) { in_dat_data6[0], in_dat_data6[1], in_dat_data6[2], in_dat_data6[3], in_dat_data6[4], in_dat_data6[5], in_dat_data6[6], in_dat_data6[7], in_dat_data7[0], in_dat_data7[1] };
  assign _08246_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27722" *) { in_dat_data4[0], in_dat_data4[1], in_dat_data4[2], in_dat_data4[3], in_dat_data4[4], in_dat_data4[5], in_dat_data4[6], in_dat_data4[7], in_dat_data5[0], in_dat_data5[1] };
  assign _08247_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27723" *) { in_dat_data2[0], in_dat_data2[1], in_dat_data2[2], in_dat_data2[3], in_dat_data2[4], in_dat_data2[5], in_dat_data2[6], in_dat_data2[7], in_dat_data3[0], in_dat_data3[1] };
  assign _08248_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27724" *) { in_dat_data0[0], in_dat_data0[1], in_dat_data0[2], in_dat_data0[3], in_dat_data0[4], in_dat_data0[5], in_dat_data0[6], in_dat_data0[7], in_dat_data1[0], in_dat_data1[1] };
  assign _08249_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2773" *) { in_wt_data35[2], in_wt_data35[3], in_wt_data35[4], in_wt_data35[5], in_wt_data35[6] };
  assign _08250_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2774" *) { in_wt_data33[2], in_wt_data33[3], in_wt_data33[4], in_wt_data33[5], in_wt_data33[6] };
  assign _08251_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2775" *) { in_wt_data31[2], in_wt_data31[3], in_wt_data31[4], in_wt_data31[5], in_wt_data31[6] };
  assign _08252_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2776" *) { in_wt_data29[2], in_wt_data29[3], in_wt_data29[4], in_wt_data29[5], in_wt_data29[6] };
  assign _08253_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2777" *) { in_wt_data27[2], in_wt_data27[3], in_wt_data27[4], in_wt_data27[5], in_wt_data27[6] };
  assign _08254_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2778" *) { in_wt_data25[2], in_wt_data25[3], in_wt_data25[4], in_wt_data25[5], in_wt_data25[6] };
  assign _08255_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2779" *) { in_wt_data23[2], in_wt_data23[3], in_wt_data23[4], in_wt_data23[5], in_wt_data23[6] };
  assign _08256_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2780" *) { in_wt_data21[2], in_wt_data21[3], in_wt_data21[4], in_wt_data21[5], in_wt_data21[6] };
  assign _08257_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27800" *) { in_dat_data127[2], in_dat_data127[3], in_dat_data127[4], in_dat_data127[5], in_dat_data127[6] };
  assign _08258_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27801" *) { in_dat_data125[2], in_dat_data125[3], in_dat_data125[4], in_dat_data125[5], in_dat_data125[6] };
  assign _08259_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27802" *) { in_dat_data123[2], in_dat_data123[3], in_dat_data123[4], in_dat_data123[5], in_dat_data123[6] };
  assign _08260_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27803" *) { in_dat_data121[2], in_dat_data121[3], in_dat_data121[4], in_dat_data121[5], in_dat_data121[6] };
  assign _08261_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27804" *) { in_dat_data119[2], in_dat_data119[3], in_dat_data119[4], in_dat_data119[5], in_dat_data119[6] };
  assign _08262_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27805" *) { in_dat_data117[2], in_dat_data117[3], in_dat_data117[4], in_dat_data117[5], in_dat_data117[6] };
  assign _08263_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27806" *) { in_dat_data115[2], in_dat_data115[3], in_dat_data115[4], in_dat_data115[5], in_dat_data115[6] };
  assign _08264_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27807" *) { in_dat_data113[2], in_dat_data113[3], in_dat_data113[4], in_dat_data113[5], in_dat_data113[6] };
  assign _08265_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27808" *) { in_dat_data111[2], in_dat_data111[3], in_dat_data111[4], in_dat_data111[5], in_dat_data111[6] };
  assign _08266_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27809" *) { in_dat_data109[2], in_dat_data109[3], in_dat_data109[4], in_dat_data109[5], in_dat_data109[6] };
  assign _08267_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2781" *) { in_wt_data19[2], in_wt_data19[3], in_wt_data19[4], in_wt_data19[5], in_wt_data19[6] };
  assign _08268_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27810" *) { in_dat_data107[2], in_dat_data107[3], in_dat_data107[4], in_dat_data107[5], in_dat_data107[6] };
  assign _08269_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27811" *) { in_dat_data105[2], in_dat_data105[3], in_dat_data105[4], in_dat_data105[5], in_dat_data105[6] };
  assign _08270_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27812" *) { in_dat_data103[2], in_dat_data103[3], in_dat_data103[4], in_dat_data103[5], in_dat_data103[6] };
  assign _08271_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27813" *) { in_dat_data101[2], in_dat_data101[3], in_dat_data101[4], in_dat_data101[5], in_dat_data101[6] };
  assign _08272_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27814" *) { in_dat_data99[2], in_dat_data99[3], in_dat_data99[4], in_dat_data99[5], in_dat_data99[6] };
  assign _08273_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27815" *) { in_dat_data97[2], in_dat_data97[3], in_dat_data97[4], in_dat_data97[5], in_dat_data97[6] };
  assign _08274_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27816" *) { in_dat_data95[2], in_dat_data95[3], in_dat_data95[4], in_dat_data95[5], in_dat_data95[6] };
  assign _08275_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27817" *) { in_dat_data93[2], in_dat_data93[3], in_dat_data93[4], in_dat_data93[5], in_dat_data93[6] };
  assign _08276_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27818" *) { in_dat_data91[2], in_dat_data91[3], in_dat_data91[4], in_dat_data91[5], in_dat_data91[6] };
  assign _08277_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27819" *) { in_dat_data89[2], in_dat_data89[3], in_dat_data89[4], in_dat_data89[5], in_dat_data89[6] };
  assign _08278_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2782" *) { in_wt_data17[2], in_wt_data17[3], in_wt_data17[4], in_wt_data17[5], in_wt_data17[6] };
  assign _08279_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27820" *) { in_dat_data87[2], in_dat_data87[3], in_dat_data87[4], in_dat_data87[5], in_dat_data87[6] };
  assign _08280_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27821" *) { in_dat_data85[2], in_dat_data85[3], in_dat_data85[4], in_dat_data85[5], in_dat_data85[6] };
  assign _08281_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27822" *) { in_dat_data83[2], in_dat_data83[3], in_dat_data83[4], in_dat_data83[5], in_dat_data83[6] };
  assign _08282_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27823" *) { in_dat_data81[2], in_dat_data81[3], in_dat_data81[4], in_dat_data81[5], in_dat_data81[6] };
  assign _08283_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27824" *) { in_dat_data79[2], in_dat_data79[3], in_dat_data79[4], in_dat_data79[5], in_dat_data79[6] };
  assign _08284_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27825" *) { in_dat_data77[2], in_dat_data77[3], in_dat_data77[4], in_dat_data77[5], in_dat_data77[6] };
  assign _08285_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27826" *) { in_dat_data75[2], in_dat_data75[3], in_dat_data75[4], in_dat_data75[5], in_dat_data75[6] };
  assign _08286_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27827" *) { in_dat_data73[2], in_dat_data73[3], in_dat_data73[4], in_dat_data73[5], in_dat_data73[6] };
  assign _08287_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27828" *) { in_dat_data71[2], in_dat_data71[3], in_dat_data71[4], in_dat_data71[5], in_dat_data71[6] };
  assign _08288_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27829" *) { in_dat_data69[2], in_dat_data69[3], in_dat_data69[4], in_dat_data69[5], in_dat_data69[6] };
  assign _08289_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2783" *) { in_wt_data15[2], in_wt_data15[3], in_wt_data15[4], in_wt_data15[5], in_wt_data15[6] };
  assign _08290_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27830" *) { in_dat_data67[2], in_dat_data67[3], in_dat_data67[4], in_dat_data67[5], in_dat_data67[6] };
  assign _08291_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27831" *) { in_dat_data65[2], in_dat_data65[3], in_dat_data65[4], in_dat_data65[5], in_dat_data65[6] };
  assign _08292_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27832" *) { in_dat_data63[2], in_dat_data63[3], in_dat_data63[4], in_dat_data63[5], in_dat_data63[6] };
  assign _08293_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27833" *) { in_dat_data61[2], in_dat_data61[3], in_dat_data61[4], in_dat_data61[5], in_dat_data61[6] };
  assign _08294_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27834" *) { in_dat_data59[2], in_dat_data59[3], in_dat_data59[4], in_dat_data59[5], in_dat_data59[6] };
  assign _08295_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27835" *) { in_dat_data57[2], in_dat_data57[3], in_dat_data57[4], in_dat_data57[5], in_dat_data57[6] };
  assign _08296_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27836" *) { in_dat_data55[2], in_dat_data55[3], in_dat_data55[4], in_dat_data55[5], in_dat_data55[6] };
  assign _08297_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27837" *) { in_dat_data53[2], in_dat_data53[3], in_dat_data53[4], in_dat_data53[5], in_dat_data53[6] };
  assign _08298_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27838" *) { in_dat_data51[2], in_dat_data51[3], in_dat_data51[4], in_dat_data51[5], in_dat_data51[6] };
  assign _08299_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27839" *) { in_dat_data49[2], in_dat_data49[3], in_dat_data49[4], in_dat_data49[5], in_dat_data49[6] };
  assign _08300_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2784" *) { in_wt_data13[2], in_wt_data13[3], in_wt_data13[4], in_wt_data13[5], in_wt_data13[6] };
  assign _08301_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27840" *) { in_dat_data47[2], in_dat_data47[3], in_dat_data47[4], in_dat_data47[5], in_dat_data47[6] };
  assign _08302_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27841" *) { in_dat_data45[2], in_dat_data45[3], in_dat_data45[4], in_dat_data45[5], in_dat_data45[6] };
  assign _08303_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27842" *) { in_dat_data43[2], in_dat_data43[3], in_dat_data43[4], in_dat_data43[5], in_dat_data43[6] };
  assign _08304_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27843" *) { in_dat_data41[2], in_dat_data41[3], in_dat_data41[4], in_dat_data41[5], in_dat_data41[6] };
  assign _08305_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27844" *) { in_dat_data39[2], in_dat_data39[3], in_dat_data39[4], in_dat_data39[5], in_dat_data39[6] };
  assign _08306_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27845" *) { in_dat_data37[2], in_dat_data37[3], in_dat_data37[4], in_dat_data37[5], in_dat_data37[6] };
  assign _08307_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27846" *) { in_dat_data35[2], in_dat_data35[3], in_dat_data35[4], in_dat_data35[5], in_dat_data35[6] };
  assign _08308_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27847" *) { in_dat_data33[2], in_dat_data33[3], in_dat_data33[4], in_dat_data33[5], in_dat_data33[6] };
  assign _08309_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27848" *) { in_dat_data31[2], in_dat_data31[3], in_dat_data31[4], in_dat_data31[5], in_dat_data31[6] };
  assign _08310_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27849" *) { in_dat_data29[2], in_dat_data29[3], in_dat_data29[4], in_dat_data29[5], in_dat_data29[6] };
  assign _08311_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2785" *) { in_wt_data11[2], in_wt_data11[3], in_wt_data11[4], in_wt_data11[5], in_wt_data11[6] };
  assign _08312_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27850" *) { in_dat_data27[2], in_dat_data27[3], in_dat_data27[4], in_dat_data27[5], in_dat_data27[6] };
  assign _08313_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27851" *) { in_dat_data25[2], in_dat_data25[3], in_dat_data25[4], in_dat_data25[5], in_dat_data25[6] };
  assign _08314_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27852" *) { in_dat_data23[2], in_dat_data23[3], in_dat_data23[4], in_dat_data23[5], in_dat_data23[6] };
  assign _08315_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27853" *) { in_dat_data21[2], in_dat_data21[3], in_dat_data21[4], in_dat_data21[5], in_dat_data21[6] };
  assign _08316_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27854" *) { in_dat_data19[2], in_dat_data19[3], in_dat_data19[4], in_dat_data19[5], in_dat_data19[6] };
  assign _08317_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27855" *) { in_dat_data17[2], in_dat_data17[3], in_dat_data17[4], in_dat_data17[5], in_dat_data17[6] };
  assign _08318_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27856" *) { in_dat_data15[2], in_dat_data15[3], in_dat_data15[4], in_dat_data15[5], in_dat_data15[6] };
  assign _08319_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27857" *) { in_dat_data13[2], in_dat_data13[3], in_dat_data13[4], in_dat_data13[5], in_dat_data13[6] };
  assign _08320_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27858" *) { in_dat_data11[2], in_dat_data11[3], in_dat_data11[4], in_dat_data11[5], in_dat_data11[6] };
  assign _08321_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27859" *) { in_dat_data9[2], in_dat_data9[3], in_dat_data9[4], in_dat_data9[5], in_dat_data9[6] };
  assign _08322_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2786" *) { in_wt_data9[2], in_wt_data9[3], in_wt_data9[4], in_wt_data9[5], in_wt_data9[6] };
  assign _08323_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27860" *) { in_dat_data7[2], in_dat_data7[3], in_dat_data7[4], in_dat_data7[5], in_dat_data7[6] };
  assign _08324_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27861" *) { in_dat_data5[2], in_dat_data5[3], in_dat_data5[4], in_dat_data5[5], in_dat_data5[6] };
  assign _08325_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27862" *) { in_dat_data3[2], in_dat_data3[3], in_dat_data3[4], in_dat_data3[5], in_dat_data3[6] };
  assign _08326_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27863" *) { in_dat_data1[2], in_dat_data1[3], in_dat_data1[4], in_dat_data1[5], in_dat_data1[6] };
  assign _08327_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2787" *) { in_wt_data7[2], in_wt_data7[3], in_wt_data7[4], in_wt_data7[5], in_wt_data7[6] };
  assign _08328_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2788" *) { in_wt_data5[2], in_wt_data5[3], in_wt_data5[4], in_wt_data5[5], in_wt_data5[6] };
  assign _08329_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2789" *) { in_wt_data3[2], in_wt_data3[3], in_wt_data3[4], in_wt_data3[5], in_wt_data3[6] };
  assign _08330_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2790" *) { in_wt_data1[2], in_wt_data1[3], in_wt_data1[4], in_wt_data1[5], in_wt_data1[6] };
  assign dat_has_nan = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28956" *) { in_dat_nan[0], in_dat_nan[1], in_dat_nan[2], in_dat_nan[3], in_dat_nan[4], in_dat_nan[5], in_dat_nan[6], in_dat_nan[7], in_dat_nan[8], in_dat_nan[9], in_dat_nan[10], in_dat_nan[11], in_dat_nan[12], in_dat_nan[13], in_dat_nan[14], in_dat_nan[15], in_dat_nan[16], in_dat_nan[17], in_dat_nan[18], in_dat_nan[19], in_dat_nan[20], in_dat_nan[21], in_dat_nan[22], in_dat_nan[23], in_dat_nan[24], in_dat_nan[25], in_dat_nan[26], in_dat_nan[27], in_dat_nan[28], in_dat_nan[29], in_dat_nan[30], in_dat_nan[31], in_dat_nan[32], in_dat_nan[33], in_dat_nan[34], in_dat_nan[35], in_dat_nan[36], in_dat_nan[37], in_dat_nan[38], in_dat_nan[39], in_dat_nan[40], in_dat_nan[41], in_dat_nan[42], in_dat_nan[43], in_dat_nan[44], in_dat_nan[45], in_dat_nan[46], in_dat_nan[47], in_dat_nan[48], in_dat_nan[49], in_dat_nan[50], in_dat_nan[51], in_dat_nan[52], in_dat_nan[53], in_dat_nan[54], in_dat_nan[55], in_dat_nan[56], in_dat_nan[57], in_dat_nan[58], in_dat_nan[59], in_dat_nan[60], in_dat_nan[61], in_dat_nan[62], in_dat_nan[63] };
  assign wt_has_nan = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3883" *) { in_wt_nan[0], in_wt_nan[1], in_wt_nan[2], in_wt_nan[3], in_wt_nan[4], in_wt_nan[5], in_wt_nan[6], in_wt_nan[7], in_wt_nan[8], in_wt_nan[9], in_wt_nan[10], in_wt_nan[11], in_wt_nan[12], in_wt_nan[13], in_wt_nan[14], in_wt_nan[15], in_wt_nan[16], in_wt_nan[17], in_wt_nan[18], in_wt_nan[19], in_wt_nan[20], in_wt_nan[21], in_wt_nan[22], in_wt_nan[23], in_wt_nan[24], in_wt_nan[25], in_wt_nan[26], in_wt_nan[27], in_wt_nan[28], in_wt_nan[29], in_wt_nan[30], in_wt_nan[31], in_wt_nan[32], in_wt_nan[33], in_wt_nan[34], in_wt_nan[35], in_wt_nan[36], in_wt_nan[37], in_wt_nan[38], in_wt_nan[39], in_wt_nan[40], in_wt_nan[41], in_wt_nan[42], in_wt_nan[43], in_wt_nan[44], in_wt_nan[45], in_wt_nan[46], in_wt_nan[47], in_wt_nan[48], in_wt_nan[49], in_wt_nan[50], in_wt_nan[51], in_wt_nan[52], in_wt_nan[53], in_wt_nan[54], in_wt_nan[55], in_wt_nan[56], in_wt_nan[57], in_wt_nan[58], in_wt_nan[59], in_wt_nan[60], in_wt_nan[61], in_wt_nan[62], in_wt_nan[63] };
  assign in_dat_data_fp16_mts_sft63 = in_dat_data_fp16_mts_ori63 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28446" *) in_dat_data127[3:2];
  assign in_dat_data_fp16_mts_sft62 = in_dat_data_fp16_mts_ori62 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28454" *) in_dat_data125[3:2];
  assign in_dat_data_fp16_mts_sft61 = in_dat_data_fp16_mts_ori61 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28462" *) in_dat_data123[3:2];
  assign in_dat_data_fp16_mts_sft60 = in_dat_data_fp16_mts_ori60 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28470" *) in_dat_data121[3:2];
  assign in_dat_data_fp16_mts_sft59 = in_dat_data_fp16_mts_ori59 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28478" *) in_dat_data119[3:2];
  assign in_dat_data_fp16_mts_sft58 = in_dat_data_fp16_mts_ori58 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28486" *) in_dat_data117[3:2];
  assign in_dat_data_fp16_mts_sft57 = in_dat_data_fp16_mts_ori57 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28494" *) in_dat_data115[3:2];
  assign in_dat_data_fp16_mts_sft56 = in_dat_data_fp16_mts_ori56 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28502" *) in_dat_data113[3:2];
  assign in_dat_data_fp16_mts_sft55 = in_dat_data_fp16_mts_ori55 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28510" *) in_dat_data111[3:2];
  assign in_dat_data_fp16_mts_sft54 = in_dat_data_fp16_mts_ori54 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28518" *) in_dat_data109[3:2];
  assign in_dat_data_fp16_mts_sft53 = in_dat_data_fp16_mts_ori53 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28526" *) in_dat_data107[3:2];
  assign in_dat_data_fp16_mts_sft52 = in_dat_data_fp16_mts_ori52 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28534" *) in_dat_data105[3:2];
  assign in_dat_data_fp16_mts_sft51 = in_dat_data_fp16_mts_ori51 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28542" *) in_dat_data103[3:2];
  assign in_dat_data_fp16_mts_sft50 = in_dat_data_fp16_mts_ori50 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28550" *) in_dat_data101[3:2];
  assign in_dat_data_fp16_mts_sft49 = in_dat_data_fp16_mts_ori49 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28558" *) in_dat_data99[3:2];
  assign in_dat_data_fp16_mts_sft48 = in_dat_data_fp16_mts_ori48 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28566" *) in_dat_data97[3:2];
  assign in_dat_data_fp16_mts_sft47 = in_dat_data_fp16_mts_ori47 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28574" *) in_dat_data95[3:2];
  assign in_dat_data_fp16_mts_sft46 = in_dat_data_fp16_mts_ori46 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28582" *) in_dat_data93[3:2];
  assign in_dat_data_fp16_mts_sft45 = in_dat_data_fp16_mts_ori45 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28590" *) in_dat_data91[3:2];
  assign in_dat_data_fp16_mts_sft44 = in_dat_data_fp16_mts_ori44 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28598" *) in_dat_data89[3:2];
  assign in_dat_data_fp16_mts_sft43 = in_dat_data_fp16_mts_ori43 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28606" *) in_dat_data87[3:2];
  assign in_dat_data_fp16_mts_sft42 = in_dat_data_fp16_mts_ori42 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28614" *) in_dat_data85[3:2];
  assign in_dat_data_fp16_mts_sft41 = in_dat_data_fp16_mts_ori41 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28622" *) in_dat_data83[3:2];
  assign in_dat_data_fp16_mts_sft40 = in_dat_data_fp16_mts_ori40 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28630" *) in_dat_data81[3:2];
  assign in_dat_data_fp16_mts_sft39 = in_dat_data_fp16_mts_ori39 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28638" *) in_dat_data79[3:2];
  assign in_dat_data_fp16_mts_sft38 = in_dat_data_fp16_mts_ori38 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28646" *) in_dat_data77[3:2];
  assign in_dat_data_fp16_mts_sft37 = in_dat_data_fp16_mts_ori37 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28654" *) in_dat_data75[3:2];
  assign in_dat_data_fp16_mts_sft36 = in_dat_data_fp16_mts_ori36 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28662" *) in_dat_data73[3:2];
  assign in_dat_data_fp16_mts_sft35 = in_dat_data_fp16_mts_ori35 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28670" *) in_dat_data71[3:2];
  assign in_dat_data_fp16_mts_sft34 = in_dat_data_fp16_mts_ori34 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28678" *) in_dat_data69[3:2];
  assign in_dat_data_fp16_mts_sft33 = in_dat_data_fp16_mts_ori33 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28686" *) in_dat_data67[3:2];
  assign in_dat_data_fp16_mts_sft32 = in_dat_data_fp16_mts_ori32 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28694" *) in_dat_data65[3:2];
  assign in_dat_data_fp16_mts_sft31 = in_dat_data_fp16_mts_ori31 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28702" *) in_dat_data63[3:2];
  assign in_dat_data_fp16_mts_sft30 = in_dat_data_fp16_mts_ori30 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28710" *) in_dat_data61[3:2];
  assign in_dat_data_fp16_mts_sft29 = in_dat_data_fp16_mts_ori29 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28718" *) in_dat_data59[3:2];
  assign in_dat_data_fp16_mts_sft28 = in_dat_data_fp16_mts_ori28 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28726" *) in_dat_data57[3:2];
  assign in_dat_data_fp16_mts_sft27 = in_dat_data_fp16_mts_ori27 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28734" *) in_dat_data55[3:2];
  assign in_dat_data_fp16_mts_sft26 = in_dat_data_fp16_mts_ori26 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28742" *) in_dat_data53[3:2];
  assign in_dat_data_fp16_mts_sft25 = in_dat_data_fp16_mts_ori25 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28750" *) in_dat_data51[3:2];
  assign in_dat_data_fp16_mts_sft24 = in_dat_data_fp16_mts_ori24 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28758" *) in_dat_data49[3:2];
  assign in_dat_data_fp16_mts_sft23 = in_dat_data_fp16_mts_ori23 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28766" *) in_dat_data47[3:2];
  assign in_dat_data_fp16_mts_sft22 = in_dat_data_fp16_mts_ori22 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28774" *) in_dat_data45[3:2];
  assign in_dat_data_fp16_mts_sft21 = in_dat_data_fp16_mts_ori21 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28782" *) in_dat_data43[3:2];
  assign in_dat_data_fp16_mts_sft20 = in_dat_data_fp16_mts_ori20 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28790" *) in_dat_data41[3:2];
  assign in_dat_data_fp16_mts_sft19 = in_dat_data_fp16_mts_ori19 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28798" *) in_dat_data39[3:2];
  assign in_dat_data_fp16_mts_sft18 = in_dat_data_fp16_mts_ori18 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28806" *) in_dat_data37[3:2];
  assign in_dat_data_fp16_mts_sft17 = in_dat_data_fp16_mts_ori17 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28814" *) in_dat_data35[3:2];
  assign in_dat_data_fp16_mts_sft16 = in_dat_data_fp16_mts_ori16 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28822" *) in_dat_data33[3:2];
  assign in_dat_data_fp16_mts_sft15 = in_dat_data_fp16_mts_ori15 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28830" *) in_dat_data31[3:2];
  assign in_dat_data_fp16_mts_sft14 = in_dat_data_fp16_mts_ori14 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28838" *) in_dat_data29[3:2];
  assign in_dat_data_fp16_mts_sft13 = in_dat_data_fp16_mts_ori13 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28846" *) in_dat_data27[3:2];
  assign in_dat_data_fp16_mts_sft12 = in_dat_data_fp16_mts_ori12 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28854" *) in_dat_data25[3:2];
  assign in_dat_data_fp16_mts_sft11 = in_dat_data_fp16_mts_ori11 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28862" *) in_dat_data23[3:2];
  assign in_dat_data_fp16_mts_sft10 = in_dat_data_fp16_mts_ori10 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28870" *) in_dat_data21[3:2];
  assign in_dat_data_fp16_mts_sft9 = in_dat_data_fp16_mts_ori9 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28878" *) in_dat_data19[3:2];
  assign in_dat_data_fp16_mts_sft8 = in_dat_data_fp16_mts_ori8 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28886" *) in_dat_data17[3:2];
  assign in_dat_data_fp16_mts_sft7 = in_dat_data_fp16_mts_ori7 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28894" *) in_dat_data15[3:2];
  assign in_dat_data_fp16_mts_sft6 = in_dat_data_fp16_mts_ori6 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28902" *) in_dat_data13[3:2];
  assign in_dat_data_fp16_mts_sft5 = in_dat_data_fp16_mts_ori5 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28910" *) in_dat_data11[3:2];
  assign in_dat_data_fp16_mts_sft4 = in_dat_data_fp16_mts_ori4 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28918" *) in_dat_data9[3:2];
  assign in_dat_data_fp16_mts_sft3 = in_dat_data_fp16_mts_ori3 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28926" *) in_dat_data7[3:2];
  assign in_dat_data_fp16_mts_sft2 = in_dat_data_fp16_mts_ori2 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28934" *) in_dat_data5[3:2];
  assign in_dat_data_fp16_mts_sft1 = in_dat_data_fp16_mts_ori1 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28942" *) in_dat_data3[3:2];
  assign in_dat_data_fp16_mts_sft0 = in_dat_data_fp16_mts_ori0 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28950" *) in_dat_data1[3:2];
  assign in_wt_data_fp16_mts_sft63 = in_wt_data_fp16_mts_ori63 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3373" *) in_wt_data127[3:2];
  assign in_wt_data_fp16_mts_sft62 = in_wt_data_fp16_mts_ori62 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3381" *) in_wt_data125[3:2];
  assign in_wt_data_fp16_mts_sft61 = in_wt_data_fp16_mts_ori61 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3389" *) in_wt_data123[3:2];
  assign in_wt_data_fp16_mts_sft60 = in_wt_data_fp16_mts_ori60 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3397" *) in_wt_data121[3:2];
  assign in_wt_data_fp16_mts_sft59 = in_wt_data_fp16_mts_ori59 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3405" *) in_wt_data119[3:2];
  assign in_wt_data_fp16_mts_sft58 = in_wt_data_fp16_mts_ori58 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3413" *) in_wt_data117[3:2];
  assign in_wt_data_fp16_mts_sft57 = in_wt_data_fp16_mts_ori57 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3421" *) in_wt_data115[3:2];
  assign in_wt_data_fp16_mts_sft56 = in_wt_data_fp16_mts_ori56 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3429" *) in_wt_data113[3:2];
  assign in_wt_data_fp16_mts_sft55 = in_wt_data_fp16_mts_ori55 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3437" *) in_wt_data111[3:2];
  assign in_wt_data_fp16_mts_sft54 = in_wt_data_fp16_mts_ori54 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3445" *) in_wt_data109[3:2];
  assign in_wt_data_fp16_mts_sft53 = in_wt_data_fp16_mts_ori53 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3453" *) in_wt_data107[3:2];
  assign in_wt_data_fp16_mts_sft52 = in_wt_data_fp16_mts_ori52 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3461" *) in_wt_data105[3:2];
  assign in_wt_data_fp16_mts_sft51 = in_wt_data_fp16_mts_ori51 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3469" *) in_wt_data103[3:2];
  assign in_wt_data_fp16_mts_sft50 = in_wt_data_fp16_mts_ori50 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3477" *) in_wt_data101[3:2];
  assign in_wt_data_fp16_mts_sft49 = in_wt_data_fp16_mts_ori49 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3485" *) in_wt_data99[3:2];
  assign in_wt_data_fp16_mts_sft48 = in_wt_data_fp16_mts_ori48 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3493" *) in_wt_data97[3:2];
  assign in_wt_data_fp16_mts_sft47 = in_wt_data_fp16_mts_ori47 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3501" *) in_wt_data95[3:2];
  assign in_wt_data_fp16_mts_sft46 = in_wt_data_fp16_mts_ori46 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3509" *) in_wt_data93[3:2];
  assign in_wt_data_fp16_mts_sft45 = in_wt_data_fp16_mts_ori45 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3517" *) in_wt_data91[3:2];
  assign in_wt_data_fp16_mts_sft44 = in_wt_data_fp16_mts_ori44 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3525" *) in_wt_data89[3:2];
  assign in_wt_data_fp16_mts_sft43 = in_wt_data_fp16_mts_ori43 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3533" *) in_wt_data87[3:2];
  assign in_wt_data_fp16_mts_sft42 = in_wt_data_fp16_mts_ori42 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3541" *) in_wt_data85[3:2];
  assign in_wt_data_fp16_mts_sft41 = in_wt_data_fp16_mts_ori41 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3549" *) in_wt_data83[3:2];
  assign in_wt_data_fp16_mts_sft40 = in_wt_data_fp16_mts_ori40 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3557" *) in_wt_data81[3:2];
  assign in_wt_data_fp16_mts_sft39 = in_wt_data_fp16_mts_ori39 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3565" *) in_wt_data79[3:2];
  assign in_wt_data_fp16_mts_sft38 = in_wt_data_fp16_mts_ori38 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3573" *) in_wt_data77[3:2];
  assign in_wt_data_fp16_mts_sft37 = in_wt_data_fp16_mts_ori37 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3581" *) in_wt_data75[3:2];
  assign in_wt_data_fp16_mts_sft36 = in_wt_data_fp16_mts_ori36 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3589" *) in_wt_data73[3:2];
  assign in_wt_data_fp16_mts_sft35 = in_wt_data_fp16_mts_ori35 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3597" *) in_wt_data71[3:2];
  assign in_wt_data_fp16_mts_sft34 = in_wt_data_fp16_mts_ori34 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3605" *) in_wt_data69[3:2];
  assign in_wt_data_fp16_mts_sft33 = in_wt_data_fp16_mts_ori33 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3613" *) in_wt_data67[3:2];
  assign in_wt_data_fp16_mts_sft32 = in_wt_data_fp16_mts_ori32 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3621" *) in_wt_data65[3:2];
  assign in_wt_data_fp16_mts_sft31 = in_wt_data_fp16_mts_ori31 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3629" *) in_wt_data63[3:2];
  assign in_wt_data_fp16_mts_sft30 = in_wt_data_fp16_mts_ori30 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3637" *) in_wt_data61[3:2];
  assign in_wt_data_fp16_mts_sft29 = in_wt_data_fp16_mts_ori29 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3645" *) in_wt_data59[3:2];
  assign in_wt_data_fp16_mts_sft28 = in_wt_data_fp16_mts_ori28 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3653" *) in_wt_data57[3:2];
  assign in_wt_data_fp16_mts_sft27 = in_wt_data_fp16_mts_ori27 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3661" *) in_wt_data55[3:2];
  assign in_wt_data_fp16_mts_sft26 = in_wt_data_fp16_mts_ori26 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3669" *) in_wt_data53[3:2];
  assign in_wt_data_fp16_mts_sft25 = in_wt_data_fp16_mts_ori25 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3677" *) in_wt_data51[3:2];
  assign in_wt_data_fp16_mts_sft24 = in_wt_data_fp16_mts_ori24 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3685" *) in_wt_data49[3:2];
  assign in_wt_data_fp16_mts_sft23 = in_wt_data_fp16_mts_ori23 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3693" *) in_wt_data47[3:2];
  assign in_wt_data_fp16_mts_sft22 = in_wt_data_fp16_mts_ori22 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3701" *) in_wt_data45[3:2];
  assign in_wt_data_fp16_mts_sft21 = in_wt_data_fp16_mts_ori21 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3709" *) in_wt_data43[3:2];
  assign in_wt_data_fp16_mts_sft20 = in_wt_data_fp16_mts_ori20 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3717" *) in_wt_data41[3:2];
  assign in_wt_data_fp16_mts_sft19 = in_wt_data_fp16_mts_ori19 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3725" *) in_wt_data39[3:2];
  assign in_wt_data_fp16_mts_sft18 = in_wt_data_fp16_mts_ori18 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3733" *) in_wt_data37[3:2];
  assign in_wt_data_fp16_mts_sft17 = in_wt_data_fp16_mts_ori17 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3741" *) in_wt_data35[3:2];
  assign in_wt_data_fp16_mts_sft16 = in_wt_data_fp16_mts_ori16 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3749" *) in_wt_data33[3:2];
  assign in_wt_data_fp16_mts_sft15 = in_wt_data_fp16_mts_ori15 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3757" *) in_wt_data31[3:2];
  assign in_wt_data_fp16_mts_sft14 = in_wt_data_fp16_mts_ori14 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3765" *) in_wt_data29[3:2];
  assign in_wt_data_fp16_mts_sft13 = in_wt_data_fp16_mts_ori13 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3773" *) in_wt_data27[3:2];
  assign in_wt_data_fp16_mts_sft12 = in_wt_data_fp16_mts_ori12 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3781" *) in_wt_data25[3:2];
  assign in_wt_data_fp16_mts_sft11 = in_wt_data_fp16_mts_ori11 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3789" *) in_wt_data23[3:2];
  assign in_wt_data_fp16_mts_sft10 = in_wt_data_fp16_mts_ori10 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3797" *) in_wt_data21[3:2];
  assign in_wt_data_fp16_mts_sft9 = in_wt_data_fp16_mts_ori9 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3805" *) in_wt_data19[3:2];
  assign in_wt_data_fp16_mts_sft8 = in_wt_data_fp16_mts_ori8 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3813" *) in_wt_data17[3:2];
  assign in_wt_data_fp16_mts_sft7 = in_wt_data_fp16_mts_ori7 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3821" *) in_wt_data15[3:2];
  assign in_wt_data_fp16_mts_sft6 = in_wt_data_fp16_mts_ori6 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3829" *) in_wt_data13[3:2];
  assign in_wt_data_fp16_mts_sft5 = in_wt_data_fp16_mts_ori5 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3837" *) in_wt_data11[3:2];
  assign in_wt_data_fp16_mts_sft4 = in_wt_data_fp16_mts_ori4 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3845" *) in_wt_data9[3:2];
  assign in_wt_data_fp16_mts_sft3 = in_wt_data_fp16_mts_ori3 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3853" *) in_wt_data7[3:2];
  assign in_wt_data_fp16_mts_sft2 = in_wt_data_fp16_mts_ori2 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3861" *) in_wt_data5[3:2];
  assign in_wt_data_fp16_mts_sft1 = in_wt_data_fp16_mts_ori1 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3869" *) in_wt_data3[3:2];
  assign in_wt_data_fp16_mts_sft0 = in_wt_data_fp16_mts_ori0 << (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3877" *) in_wt_data1[3:2];
  assign _08331_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10666" *) 1'b0 : wt4_sd_pvld;
  assign wt4_sd_pvld_w = wt_pre_sel[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:10666" *) 1'b1 : _08331_;
  assign _08332_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12002" *) 1'b0 : wt5_sd_pvld;
  assign wt5_sd_pvld_w = wt_pre_sel[5] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:12002" *) 1'b1 : _08332_;
  assign _08333_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13338" *) 1'b0 : wt6_sd_pvld;
  assign wt6_sd_pvld_w = wt_pre_sel[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:13338" *) 1'b1 : _08333_;
  assign _08334_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14674" *) 1'b0 : wt7_sd_pvld;
  assign wt7_sd_pvld_w = wt_pre_sel[7] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:14674" *) 1'b1 : _08334_;
  assign _08335_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16011" *) 1'b0 : wt0_actv_pvld[0];
  assign wt0_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:16011" *) wt0_sd_pvld : _08335_;
  assign _08336_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17335" *) 1'b0 : wt1_actv_pvld[0];
  assign wt1_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:17335" *) wt1_sd_pvld : _08336_;
  assign _08337_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18659" *) 1'b0 : wt2_actv_pvld[0];
  assign wt2_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:18659" *) wt2_sd_pvld : _08337_;
  assign _08338_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19983" *) 1'b0 : wt3_actv_pvld[0];
  assign wt3_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:19983" *) wt3_sd_pvld : _08338_;
  assign _08339_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21307" *) 1'b0 : wt4_actv_pvld[0];
  assign wt4_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:21307" *) wt4_sd_pvld : _08339_;
  assign _08340_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22631" *) 1'b0 : wt5_actv_pvld[0];
  assign wt5_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:22631" *) wt5_sd_pvld : _08340_;
  assign _08341_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23955" *) 1'b0 : wt6_actv_pvld[0];
  assign wt6_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:23955" *) wt6_sd_pvld : _08341_;
  assign _08342_ = dat_actv_stripe_end ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25279" *) 1'b0 : wt7_actv_pvld[0];
  assign wt7_actv_pvld_w = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:25279" *) wt7_sd_pvld : _08342_;
  assign _06279_[10:0] = in_dat_norm[63] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27872" *) { 1'b1, in_dat_data127[1:0], in_dat_data126 } : { in_dat_data127[1:0], in_dat_data126, 1'b0 };
  assign in_dat_data_fp16_mts_ori63 = cfg_is_fp16_d1[63] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27872" *) _06279_[10:0] : 11'b00000000000;
  assign _06280_[10:0] = in_dat_norm[62] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27881" *) { 1'b1, in_dat_data125[1:0], in_dat_data124 } : { in_dat_data125[1:0], in_dat_data124, 1'b0 };
  assign in_dat_data_fp16_mts_ori62 = cfg_is_fp16_d1[62] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27881" *) _06280_[10:0] : 11'b00000000000;
  assign _06281_[10:0] = in_dat_norm[61] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27890" *) { 1'b1, in_dat_data123[1:0], in_dat_data122 } : { in_dat_data123[1:0], in_dat_data122, 1'b0 };
  assign in_dat_data_fp16_mts_ori61 = cfg_is_fp16_d1[61] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27890" *) _06281_[10:0] : 11'b00000000000;
  assign _06282_[10:0] = in_dat_norm[60] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27899" *) { 1'b1, in_dat_data121[1:0], in_dat_data120 } : { in_dat_data121[1:0], in_dat_data120, 1'b0 };
  assign in_dat_data_fp16_mts_ori60 = cfg_is_fp16_d1[60] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27899" *) _06282_[10:0] : 11'b00000000000;
  assign _06283_[10:0] = in_dat_norm[59] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27908" *) { 1'b1, in_dat_data119[1:0], in_dat_data118 } : { in_dat_data119[1:0], in_dat_data118, 1'b0 };
  assign in_dat_data_fp16_mts_ori59 = cfg_is_fp16_d1[59] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27908" *) _06283_[10:0] : 11'b00000000000;
  assign _06284_[10:0] = in_dat_norm[58] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27917" *) { 1'b1, in_dat_data117[1:0], in_dat_data116 } : { in_dat_data117[1:0], in_dat_data116, 1'b0 };
  assign in_dat_data_fp16_mts_ori58 = cfg_is_fp16_d1[58] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27917" *) _06284_[10:0] : 11'b00000000000;
  assign _06285_[10:0] = in_dat_norm[57] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27926" *) { 1'b1, in_dat_data115[1:0], in_dat_data114 } : { in_dat_data115[1:0], in_dat_data114, 1'b0 };
  assign in_dat_data_fp16_mts_ori57 = cfg_is_fp16_d1[57] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27926" *) _06285_[10:0] : 11'b00000000000;
  assign _06286_[10:0] = in_dat_norm[56] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27935" *) { 1'b1, in_dat_data113[1:0], in_dat_data112 } : { in_dat_data113[1:0], in_dat_data112, 1'b0 };
  assign in_dat_data_fp16_mts_ori56 = cfg_is_fp16_d1[56] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27935" *) _06286_[10:0] : 11'b00000000000;
  assign _06287_[10:0] = in_dat_norm[55] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27944" *) { 1'b1, in_dat_data111[1:0], in_dat_data110 } : { in_dat_data111[1:0], in_dat_data110, 1'b0 };
  assign in_dat_data_fp16_mts_ori55 = cfg_is_fp16_d1[55] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27944" *) _06287_[10:0] : 11'b00000000000;
  assign _06288_[10:0] = in_dat_norm[54] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27953" *) { 1'b1, in_dat_data109[1:0], in_dat_data108 } : { in_dat_data109[1:0], in_dat_data108, 1'b0 };
  assign in_dat_data_fp16_mts_ori54 = cfg_is_fp16_d1[54] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27953" *) _06288_[10:0] : 11'b00000000000;
  assign _06289_[10:0] = in_dat_norm[53] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27962" *) { 1'b1, in_dat_data107[1:0], in_dat_data106 } : { in_dat_data107[1:0], in_dat_data106, 1'b0 };
  assign in_dat_data_fp16_mts_ori53 = cfg_is_fp16_d1[53] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27962" *) _06289_[10:0] : 11'b00000000000;
  assign _06290_[10:0] = in_dat_norm[52] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27971" *) { 1'b1, in_dat_data105[1:0], in_dat_data104 } : { in_dat_data105[1:0], in_dat_data104, 1'b0 };
  assign in_dat_data_fp16_mts_ori52 = cfg_is_fp16_d1[52] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27971" *) _06290_[10:0] : 11'b00000000000;
  assign _06291_[10:0] = in_dat_norm[51] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27980" *) { 1'b1, in_dat_data103[1:0], in_dat_data102 } : { in_dat_data103[1:0], in_dat_data102, 1'b0 };
  assign in_dat_data_fp16_mts_ori51 = cfg_is_fp16_d1[51] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27980" *) _06291_[10:0] : 11'b00000000000;
  assign _06292_[10:0] = in_dat_norm[50] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27989" *) { 1'b1, in_dat_data101[1:0], in_dat_data100 } : { in_dat_data101[1:0], in_dat_data100, 1'b0 };
  assign in_dat_data_fp16_mts_ori50 = cfg_is_fp16_d1[50] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27989" *) _06292_[10:0] : 11'b00000000000;
  assign _06293_[10:0] = in_wt_norm[63] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2799" *) { 1'b1, in_wt_data127[1:0], in_wt_data126 } : { in_wt_data127[1:0], in_wt_data126, 1'b0 };
  assign in_wt_data_fp16_mts_ori63 = cfg_is_fp16_d1[63] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2799" *) _06293_[10:0] : 11'b00000000000;
  assign _06294_[10:0] = in_dat_norm[49] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27998" *) { 1'b1, in_dat_data99[1:0], in_dat_data98 } : { in_dat_data99[1:0], in_dat_data98, 1'b0 };
  assign in_dat_data_fp16_mts_ori49 = cfg_is_fp16_d1[49] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:27998" *) _06294_[10:0] : 11'b00000000000;
  assign _06295_[10:0] = in_dat_norm[48] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28007" *) { 1'b1, in_dat_data97[1:0], in_dat_data96 } : { in_dat_data97[1:0], in_dat_data96, 1'b0 };
  assign in_dat_data_fp16_mts_ori48 = cfg_is_fp16_d1[48] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28007" *) _06295_[10:0] : 11'b00000000000;
  assign _06296_[10:0] = in_dat_norm[47] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28016" *) { 1'b1, in_dat_data95[1:0], in_dat_data94 } : { in_dat_data95[1:0], in_dat_data94, 1'b0 };
  assign in_dat_data_fp16_mts_ori47 = cfg_is_fp16_d1[47] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28016" *) _06296_[10:0] : 11'b00000000000;
  assign _06297_[10:0] = in_dat_norm[46] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28025" *) { 1'b1, in_dat_data93[1:0], in_dat_data92 } : { in_dat_data93[1:0], in_dat_data92, 1'b0 };
  assign in_dat_data_fp16_mts_ori46 = cfg_is_fp16_d1[46] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28025" *) _06297_[10:0] : 11'b00000000000;
  assign _06298_[10:0] = in_dat_norm[45] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28034" *) { 1'b1, in_dat_data91[1:0], in_dat_data90 } : { in_dat_data91[1:0], in_dat_data90, 1'b0 };
  assign in_dat_data_fp16_mts_ori45 = cfg_is_fp16_d1[45] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28034" *) _06298_[10:0] : 11'b00000000000;
  assign _06299_[10:0] = in_dat_norm[44] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28043" *) { 1'b1, in_dat_data89[1:0], in_dat_data88 } : { in_dat_data89[1:0], in_dat_data88, 1'b0 };
  assign in_dat_data_fp16_mts_ori44 = cfg_is_fp16_d1[44] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28043" *) _06299_[10:0] : 11'b00000000000;
  assign _06300_[10:0] = in_dat_norm[43] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28052" *) { 1'b1, in_dat_data87[1:0], in_dat_data86 } : { in_dat_data87[1:0], in_dat_data86, 1'b0 };
  assign in_dat_data_fp16_mts_ori43 = cfg_is_fp16_d1[43] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28052" *) _06300_[10:0] : 11'b00000000000;
  assign _06301_[10:0] = in_dat_norm[42] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28061" *) { 1'b1, in_dat_data85[1:0], in_dat_data84 } : { in_dat_data85[1:0], in_dat_data84, 1'b0 };
  assign in_dat_data_fp16_mts_ori42 = cfg_is_fp16_d1[42] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28061" *) _06301_[10:0] : 11'b00000000000;
  assign _06302_[10:0] = in_dat_norm[41] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28070" *) { 1'b1, in_dat_data83[1:0], in_dat_data82 } : { in_dat_data83[1:0], in_dat_data82, 1'b0 };
  assign in_dat_data_fp16_mts_ori41 = cfg_is_fp16_d1[41] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28070" *) _06302_[10:0] : 11'b00000000000;
  assign _06303_[10:0] = in_dat_norm[40] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28079" *) { 1'b1, in_dat_data81[1:0], in_dat_data80 } : { in_dat_data81[1:0], in_dat_data80, 1'b0 };
  assign in_dat_data_fp16_mts_ori40 = cfg_is_fp16_d1[40] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28079" *) _06303_[10:0] : 11'b00000000000;
  assign _06304_[10:0] = in_wt_norm[62] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2808" *) { 1'b1, in_wt_data125[1:0], in_wt_data124 } : { in_wt_data125[1:0], in_wt_data124, 1'b0 };
  assign in_wt_data_fp16_mts_ori62 = cfg_is_fp16_d1[62] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2808" *) _06304_[10:0] : 11'b00000000000;
  assign _06305_[10:0] = in_dat_norm[39] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28088" *) { 1'b1, in_dat_data79[1:0], in_dat_data78 } : { in_dat_data79[1:0], in_dat_data78, 1'b0 };
  assign in_dat_data_fp16_mts_ori39 = cfg_is_fp16_d1[39] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28088" *) _06305_[10:0] : 11'b00000000000;
  assign _06306_[10:0] = in_dat_norm[38] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28097" *) { 1'b1, in_dat_data77[1:0], in_dat_data76 } : { in_dat_data77[1:0], in_dat_data76, 1'b0 };
  assign in_dat_data_fp16_mts_ori38 = cfg_is_fp16_d1[38] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28097" *) _06306_[10:0] : 11'b00000000000;
  assign _06307_[10:0] = in_dat_norm[37] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28106" *) { 1'b1, in_dat_data75[1:0], in_dat_data74 } : { in_dat_data75[1:0], in_dat_data74, 1'b0 };
  assign in_dat_data_fp16_mts_ori37 = cfg_is_fp16_d1[37] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28106" *) _06307_[10:0] : 11'b00000000000;
  assign _06308_[10:0] = in_dat_norm[36] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28115" *) { 1'b1, in_dat_data73[1:0], in_dat_data72 } : { in_dat_data73[1:0], in_dat_data72, 1'b0 };
  assign in_dat_data_fp16_mts_ori36 = cfg_is_fp16_d1[36] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28115" *) _06308_[10:0] : 11'b00000000000;
  assign _06309_[10:0] = in_dat_norm[35] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28124" *) { 1'b1, in_dat_data71[1:0], in_dat_data70 } : { in_dat_data71[1:0], in_dat_data70, 1'b0 };
  assign in_dat_data_fp16_mts_ori35 = cfg_is_fp16_d1[35] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28124" *) _06309_[10:0] : 11'b00000000000;
  assign _06310_[10:0] = in_dat_norm[34] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28133" *) { 1'b1, in_dat_data69[1:0], in_dat_data68 } : { in_dat_data69[1:0], in_dat_data68, 1'b0 };
  assign in_dat_data_fp16_mts_ori34 = cfg_is_fp16_d1[34] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28133" *) _06310_[10:0] : 11'b00000000000;
  assign _06311_[10:0] = in_dat_norm[33] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28142" *) { 1'b1, in_dat_data67[1:0], in_dat_data66 } : { in_dat_data67[1:0], in_dat_data66, 1'b0 };
  assign in_dat_data_fp16_mts_ori33 = cfg_is_fp16_d1[33] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28142" *) _06311_[10:0] : 11'b00000000000;
  assign _06312_[10:0] = in_dat_norm[32] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28151" *) { 1'b1, in_dat_data65[1:0], in_dat_data64 } : { in_dat_data65[1:0], in_dat_data64, 1'b0 };
  assign in_dat_data_fp16_mts_ori32 = cfg_is_fp16_d1[32] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28151" *) _06312_[10:0] : 11'b00000000000;
  assign _06313_[10:0] = in_dat_norm[31] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28160" *) { 1'b1, in_dat_data63[1:0], in_dat_data62 } : { in_dat_data63[1:0], in_dat_data62, 1'b0 };
  assign in_dat_data_fp16_mts_ori31 = cfg_is_fp16_d1[31] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28160" *) _06313_[10:0] : 11'b00000000000;
  assign _06314_[10:0] = in_dat_norm[30] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28169" *) { 1'b1, in_dat_data61[1:0], in_dat_data60 } : { in_dat_data61[1:0], in_dat_data60, 1'b0 };
  assign in_dat_data_fp16_mts_ori30 = cfg_is_fp16_d1[30] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28169" *) _06314_[10:0] : 11'b00000000000;
  assign _06315_[10:0] = in_wt_norm[61] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2817" *) { 1'b1, in_wt_data123[1:0], in_wt_data122 } : { in_wt_data123[1:0], in_wt_data122, 1'b0 };
  assign in_wt_data_fp16_mts_ori61 = cfg_is_fp16_d1[61] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2817" *) _06315_[10:0] : 11'b00000000000;
  assign _06316_[10:0] = in_dat_norm[29] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28178" *) { 1'b1, in_dat_data59[1:0], in_dat_data58 } : { in_dat_data59[1:0], in_dat_data58, 1'b0 };
  assign in_dat_data_fp16_mts_ori29 = cfg_is_fp16_d1[29] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28178" *) _06316_[10:0] : 11'b00000000000;
  assign _06317_[10:0] = in_dat_norm[28] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28187" *) { 1'b1, in_dat_data57[1:0], in_dat_data56 } : { in_dat_data57[1:0], in_dat_data56, 1'b0 };
  assign in_dat_data_fp16_mts_ori28 = cfg_is_fp16_d1[28] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28187" *) _06317_[10:0] : 11'b00000000000;
  assign _06318_[10:0] = in_dat_norm[27] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28196" *) { 1'b1, in_dat_data55[1:0], in_dat_data54 } : { in_dat_data55[1:0], in_dat_data54, 1'b0 };
  assign in_dat_data_fp16_mts_ori27 = cfg_is_fp16_d1[27] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28196" *) _06318_[10:0] : 11'b00000000000;
  assign _06319_[10:0] = in_dat_norm[26] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28205" *) { 1'b1, in_dat_data53[1:0], in_dat_data52 } : { in_dat_data53[1:0], in_dat_data52, 1'b0 };
  assign in_dat_data_fp16_mts_ori26 = cfg_is_fp16_d1[26] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28205" *) _06319_[10:0] : 11'b00000000000;
  assign _06320_[10:0] = in_dat_norm[25] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28214" *) { 1'b1, in_dat_data51[1:0], in_dat_data50 } : { in_dat_data51[1:0], in_dat_data50, 1'b0 };
  assign in_dat_data_fp16_mts_ori25 = cfg_is_fp16_d1[25] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28214" *) _06320_[10:0] : 11'b00000000000;
  assign _06321_[10:0] = in_dat_norm[24] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28223" *) { 1'b1, in_dat_data49[1:0], in_dat_data48 } : { in_dat_data49[1:0], in_dat_data48, 1'b0 };
  assign in_dat_data_fp16_mts_ori24 = cfg_is_fp16_d1[24] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28223" *) _06321_[10:0] : 11'b00000000000;
  assign _06322_[10:0] = in_dat_norm[23] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28232" *) { 1'b1, in_dat_data47[1:0], in_dat_data46 } : { in_dat_data47[1:0], in_dat_data46, 1'b0 };
  assign in_dat_data_fp16_mts_ori23 = cfg_is_fp16_d1[23] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28232" *) _06322_[10:0] : 11'b00000000000;
  assign _06323_[10:0] = in_dat_norm[22] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28241" *) { 1'b1, in_dat_data45[1:0], in_dat_data44 } : { in_dat_data45[1:0], in_dat_data44, 1'b0 };
  assign in_dat_data_fp16_mts_ori22 = cfg_is_fp16_d1[22] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28241" *) _06323_[10:0] : 11'b00000000000;
  assign _06324_[10:0] = in_dat_norm[21] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28250" *) { 1'b1, in_dat_data43[1:0], in_dat_data42 } : { in_dat_data43[1:0], in_dat_data42, 1'b0 };
  assign in_dat_data_fp16_mts_ori21 = cfg_is_fp16_d1[21] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28250" *) _06324_[10:0] : 11'b00000000000;
  assign _06325_[10:0] = in_dat_norm[20] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28259" *) { 1'b1, in_dat_data41[1:0], in_dat_data40 } : { in_dat_data41[1:0], in_dat_data40, 1'b0 };
  assign in_dat_data_fp16_mts_ori20 = cfg_is_fp16_d1[20] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28259" *) _06325_[10:0] : 11'b00000000000;
  assign _06326_[10:0] = in_wt_norm[60] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2826" *) { 1'b1, in_wt_data121[1:0], in_wt_data120 } : { in_wt_data121[1:0], in_wt_data120, 1'b0 };
  assign in_wt_data_fp16_mts_ori60 = cfg_is_fp16_d1[60] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2826" *) _06326_[10:0] : 11'b00000000000;
  assign _06327_[10:0] = in_dat_norm[19] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28268" *) { 1'b1, in_dat_data39[1:0], in_dat_data38 } : { in_dat_data39[1:0], in_dat_data38, 1'b0 };
  assign in_dat_data_fp16_mts_ori19 = cfg_is_fp16_d1[19] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28268" *) _06327_[10:0] : 11'b00000000000;
  assign _06328_[10:0] = in_dat_norm[18] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28277" *) { 1'b1, in_dat_data37[1:0], in_dat_data36 } : { in_dat_data37[1:0], in_dat_data36, 1'b0 };
  assign in_dat_data_fp16_mts_ori18 = cfg_is_fp16_d1[18] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28277" *) _06328_[10:0] : 11'b00000000000;
  assign _06329_[10:0] = in_dat_norm[17] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28286" *) { 1'b1, in_dat_data35[1:0], in_dat_data34 } : { in_dat_data35[1:0], in_dat_data34, 1'b0 };
  assign in_dat_data_fp16_mts_ori17 = cfg_is_fp16_d1[17] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28286" *) _06329_[10:0] : 11'b00000000000;
  assign _06330_[10:0] = in_dat_norm[16] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28295" *) { 1'b1, in_dat_data33[1:0], in_dat_data32 } : { in_dat_data33[1:0], in_dat_data32, 1'b0 };
  assign in_dat_data_fp16_mts_ori16 = cfg_is_fp16_d1[16] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28295" *) _06330_[10:0] : 11'b00000000000;
  assign _06331_[10:0] = in_dat_norm[15] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28304" *) { 1'b1, in_dat_data31[1:0], in_dat_data30 } : { in_dat_data31[1:0], in_dat_data30, 1'b0 };
  assign in_dat_data_fp16_mts_ori15 = cfg_is_fp16_d1[15] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28304" *) _06331_[10:0] : 11'b00000000000;
  assign _06332_[10:0] = in_dat_norm[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28313" *) { 1'b1, in_dat_data29[1:0], in_dat_data28 } : { in_dat_data29[1:0], in_dat_data28, 1'b0 };
  assign in_dat_data_fp16_mts_ori14 = cfg_is_fp16_d1[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28313" *) _06332_[10:0] : 11'b00000000000;
  assign _06333_[10:0] = in_dat_norm[13] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28322" *) { 1'b1, in_dat_data27[1:0], in_dat_data26 } : { in_dat_data27[1:0], in_dat_data26, 1'b0 };
  assign in_dat_data_fp16_mts_ori13 = cfg_is_fp16_d1[13] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28322" *) _06333_[10:0] : 11'b00000000000;
  assign _06334_[10:0] = in_dat_norm[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28331" *) { 1'b1, in_dat_data25[1:0], in_dat_data24 } : { in_dat_data25[1:0], in_dat_data24, 1'b0 };
  assign in_dat_data_fp16_mts_ori12 = cfg_is_fp16_d1[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28331" *) _06334_[10:0] : 11'b00000000000;
  assign _06335_[10:0] = in_dat_norm[11] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28340" *) { 1'b1, in_dat_data23[1:0], in_dat_data22 } : { in_dat_data23[1:0], in_dat_data22, 1'b0 };
  assign in_dat_data_fp16_mts_ori11 = cfg_is_fp16_d1[11] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28340" *) _06335_[10:0] : 11'b00000000000;
  assign _06336_[10:0] = in_dat_norm[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28349" *) { 1'b1, in_dat_data21[1:0], in_dat_data20 } : { in_dat_data21[1:0], in_dat_data20, 1'b0 };
  assign in_dat_data_fp16_mts_ori10 = cfg_is_fp16_d1[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28349" *) _06336_[10:0] : 11'b00000000000;
  assign _06337_[10:0] = in_wt_norm[59] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2835" *) { 1'b1, in_wt_data119[1:0], in_wt_data118 } : { in_wt_data119[1:0], in_wt_data118, 1'b0 };
  assign in_wt_data_fp16_mts_ori59 = cfg_is_fp16_d1[59] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2835" *) _06337_[10:0] : 11'b00000000000;
  assign _06338_[10:0] = in_dat_norm[9] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28358" *) { 1'b1, in_dat_data19[1:0], in_dat_data18 } : { in_dat_data19[1:0], in_dat_data18, 1'b0 };
  assign in_dat_data_fp16_mts_ori9 = cfg_is_fp16_d1[9] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28358" *) _06338_[10:0] : 11'b00000000000;
  assign _06339_[10:0] = in_dat_norm[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28367" *) { 1'b1, in_dat_data17[1:0], in_dat_data16 } : { in_dat_data17[1:0], in_dat_data16, 1'b0 };
  assign in_dat_data_fp16_mts_ori8 = cfg_is_fp16_d1[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28367" *) _06339_[10:0] : 11'b00000000000;
  assign _06340_[10:0] = in_dat_norm[7] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28376" *) { 1'b1, in_dat_data15[1:0], in_dat_data14 } : { in_dat_data15[1:0], in_dat_data14, 1'b0 };
  assign in_dat_data_fp16_mts_ori7 = cfg_is_fp16_d1[7] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28376" *) _06340_[10:0] : 11'b00000000000;
  assign _06341_[10:0] = in_dat_norm[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28385" *) { 1'b1, in_dat_data13[1:0], in_dat_data12 } : { in_dat_data13[1:0], in_dat_data12, 1'b0 };
  assign in_dat_data_fp16_mts_ori6 = cfg_is_fp16_d1[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28385" *) _06341_[10:0] : 11'b00000000000;
  assign _06342_[10:0] = in_dat_norm[5] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28394" *) { 1'b1, in_dat_data11[1:0], in_dat_data10 } : { in_dat_data11[1:0], in_dat_data10, 1'b0 };
  assign in_dat_data_fp16_mts_ori5 = cfg_is_fp16_d1[5] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28394" *) _06342_[10:0] : 11'b00000000000;
  assign _06343_[10:0] = in_dat_norm[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28403" *) { 1'b1, in_dat_data9[1:0], in_dat_data8 } : { in_dat_data9[1:0], in_dat_data8, 1'b0 };
  assign in_dat_data_fp16_mts_ori4 = cfg_is_fp16_d1[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28403" *) _06343_[10:0] : 11'b00000000000;
  assign _06344_[10:0] = in_dat_norm[3] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28412" *) { 1'b1, in_dat_data7[1:0], in_dat_data6 } : { in_dat_data7[1:0], in_dat_data6, 1'b0 };
  assign in_dat_data_fp16_mts_ori3 = cfg_is_fp16_d1[3] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28412" *) _06344_[10:0] : 11'b00000000000;
  assign _06345_[10:0] = in_dat_norm[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28421" *) { 1'b1, in_dat_data5[1:0], in_dat_data4 } : { in_dat_data5[1:0], in_dat_data4, 1'b0 };
  assign in_dat_data_fp16_mts_ori2 = cfg_is_fp16_d1[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28421" *) _06345_[10:0] : 11'b00000000000;
  assign _06346_[10:0] = in_dat_norm[1] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28430" *) { 1'b1, in_dat_data3[1:0], in_dat_data2 } : { in_dat_data3[1:0], in_dat_data2, 1'b0 };
  assign in_dat_data_fp16_mts_ori1 = cfg_is_fp16_d1[1] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28430" *) _06346_[10:0] : 11'b00000000000;
  assign _06347_[10:0] = in_dat_norm[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28439" *) { 1'b1, in_dat_data1[1:0], in_dat_data0 } : { in_dat_data1[1:0], in_dat_data0, 1'b0 };
  assign in_dat_data_fp16_mts_ori0 = cfg_is_fp16_d1[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:28439" *) _06347_[10:0] : 11'b00000000000;
  assign _06348_[10:0] = in_wt_norm[58] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2844" *) { 1'b1, in_wt_data117[1:0], in_wt_data116 } : { in_wt_data117[1:0], in_wt_data116, 1'b0 };
  assign in_wt_data_fp16_mts_ori58 = cfg_is_fp16_d1[58] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2844" *) _06348_[10:0] : 11'b00000000000;
  assign _06349_[10:0] = in_wt_norm[57] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2853" *) { 1'b1, in_wt_data115[1:0], in_wt_data114 } : { in_wt_data115[1:0], in_wt_data114, 1'b0 };
  assign in_wt_data_fp16_mts_ori57 = cfg_is_fp16_d1[57] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2853" *) _06349_[10:0] : 11'b00000000000;
  assign _06350_[10:0] = in_wt_norm[56] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2862" *) { 1'b1, in_wt_data113[1:0], in_wt_data112 } : { in_wt_data113[1:0], in_wt_data112, 1'b0 };
  assign in_wt_data_fp16_mts_ori56 = cfg_is_fp16_d1[56] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2862" *) _06350_[10:0] : 11'b00000000000;
  assign _06351_[10:0] = in_wt_norm[55] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2871" *) { 1'b1, in_wt_data111[1:0], in_wt_data110 } : { in_wt_data111[1:0], in_wt_data110, 1'b0 };
  assign in_wt_data_fp16_mts_ori55 = cfg_is_fp16_d1[55] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2871" *) _06351_[10:0] : 11'b00000000000;
  assign _06352_[10:0] = in_wt_norm[54] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2880" *) { 1'b1, in_wt_data109[1:0], in_wt_data108 } : { in_wt_data109[1:0], in_wt_data108, 1'b0 };
  assign in_wt_data_fp16_mts_ori54 = cfg_is_fp16_d1[54] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2880" *) _06352_[10:0] : 11'b00000000000;
  assign _06353_[10:0] = in_wt_norm[53] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2889" *) { 1'b1, in_wt_data107[1:0], in_wt_data106 } : { in_wt_data107[1:0], in_wt_data106, 1'b0 };
  assign in_wt_data_fp16_mts_ori53 = cfg_is_fp16_d1[53] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2889" *) _06353_[10:0] : 11'b00000000000;
  assign _06354_[10:0] = in_wt_norm[52] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2898" *) { 1'b1, in_wt_data105[1:0], in_wt_data104 } : { in_wt_data105[1:0], in_wt_data104, 1'b0 };
  assign in_wt_data_fp16_mts_ori52 = cfg_is_fp16_d1[52] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2898" *) _06354_[10:0] : 11'b00000000000;
  assign _08343_[126:0] = cfg_is_int8_d1[64] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29043" *) { in_dat_mask[63], in_dat_mask[126], in_dat_mask[62], in_dat_mask[125], in_dat_mask[61], in_dat_mask[124], in_dat_mask[60], in_dat_mask[123], in_dat_mask[59], in_dat_mask[122], in_dat_mask[58], in_dat_mask[121], in_dat_mask[57], in_dat_mask[120], in_dat_mask[56], in_dat_mask[119], in_dat_mask[55], in_dat_mask[118], in_dat_mask[54], in_dat_mask[117], in_dat_mask[53], in_dat_mask[116], in_dat_mask[52], in_dat_mask[115], in_dat_mask[51], in_dat_mask[114], in_dat_mask[50], in_dat_mask[113], in_dat_mask[49], in_dat_mask[112], in_dat_mask[48], in_dat_mask[111], in_dat_mask[47], in_dat_mask[110], in_dat_mask[46], in_dat_mask[109], in_dat_mask[45], in_dat_mask[108], in_dat_mask[44], in_dat_mask[107], in_dat_mask[43], in_dat_mask[106], in_dat_mask[42], in_dat_mask[105], in_dat_mask[41], in_dat_mask[104], in_dat_mask[40], in_dat_mask[103], in_dat_mask[39], in_dat_mask[102], in_dat_mask[38], in_dat_mask[101], in_dat_mask[37], in_dat_mask[100], in_dat_mask[36], in_dat_mask[99], in_dat_mask[35], in_dat_mask[98], in_dat_mask[34], in_dat_mask[97], in_dat_mask[33], in_dat_mask[96], in_dat_mask[32], in_dat_mask[95], in_dat_mask[31], in_dat_mask[94], in_dat_mask[30], in_dat_mask[93], in_dat_mask[29], in_dat_mask[92], in_dat_mask[28], in_dat_mask[91], in_dat_mask[27], in_dat_mask[90], in_dat_mask[26], in_dat_mask[89], in_dat_mask[25], in_dat_mask[88], in_dat_mask[24], in_dat_mask[87], in_dat_mask[23], in_dat_mask[86], in_dat_mask[22], in_dat_mask[85], in_dat_mask[21], in_dat_mask[84], in_dat_mask[20], in_dat_mask[83], in_dat_mask[19], in_dat_mask[82], in_dat_mask[18], in_dat_mask[81], in_dat_mask[17], in_dat_mask[80], in_dat_mask[16], in_dat_mask[79], in_dat_mask[15], in_dat_mask[78], in_dat_mask[14], in_dat_mask[77], in_dat_mask[13], in_dat_mask[76], in_dat_mask[12], in_dat_mask[75], in_dat_mask[11], in_dat_mask[74], in_dat_mask[10], in_dat_mask[73], in_dat_mask[9], in_dat_mask[72], in_dat_mask[8], in_dat_mask[71], in_dat_mask[7], in_dat_mask[70], in_dat_mask[6], in_dat_mask[69], in_dat_mask[5], in_dat_mask[68], in_dat_mask[4], in_dat_mask[67], in_dat_mask[3], in_dat_mask[66], in_dat_mask[2], in_dat_mask[65], in_dat_mask[1], in_dat_mask[64], in_dat_mask[0] } : in_dat_mask[126:0];
  assign dat_pre_nz_w = cfg_is_fp16_d1[64] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:29043" *) _05425_ : { in_dat_mask[127], _08343_[126:0] };
  assign _06355_[10:0] = in_wt_norm[51] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2907" *) { 1'b1, in_wt_data103[1:0], in_wt_data102 } : { in_wt_data103[1:0], in_wt_data102, 1'b0 };
  assign in_wt_data_fp16_mts_ori51 = cfg_is_fp16_d1[51] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2907" *) _06355_[10:0] : 11'b00000000000;
  assign _06356_[10:0] = in_wt_norm[50] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2916" *) { 1'b1, in_wt_data101[1:0], in_wt_data100 } : { in_wt_data101[1:0], in_wt_data100, 1'b0 };
  assign in_wt_data_fp16_mts_ori50 = cfg_is_fp16_d1[50] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2916" *) _06356_[10:0] : 11'b00000000000;
  assign _06357_[10:0] = in_wt_norm[49] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2925" *) { 1'b1, in_wt_data99[1:0], in_wt_data98 } : { in_wt_data99[1:0], in_wt_data98, 1'b0 };
  assign in_wt_data_fp16_mts_ori49 = cfg_is_fp16_d1[49] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2925" *) _06357_[10:0] : 11'b00000000000;
  assign _06358_[10:0] = in_wt_norm[48] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2934" *) { 1'b1, in_wt_data97[1:0], in_wt_data96 } : { in_wt_data97[1:0], in_wt_data96, 1'b0 };
  assign in_wt_data_fp16_mts_ori48 = cfg_is_fp16_d1[48] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2934" *) _06358_[10:0] : 11'b00000000000;
  assign _06359_[10:0] = in_wt_norm[47] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2943" *) { 1'b1, in_wt_data95[1:0], in_wt_data94 } : { in_wt_data95[1:0], in_wt_data94, 1'b0 };
  assign in_wt_data_fp16_mts_ori47 = cfg_is_fp16_d1[47] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2943" *) _06359_[10:0] : 11'b00000000000;
  assign _06360_[10:0] = in_wt_norm[46] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2952" *) { 1'b1, in_wt_data93[1:0], in_wt_data92 } : { in_wt_data93[1:0], in_wt_data92, 1'b0 };
  assign in_wt_data_fp16_mts_ori46 = cfg_is_fp16_d1[46] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2952" *) _06360_[10:0] : 11'b00000000000;
  assign _06361_[10:0] = in_wt_norm[45] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2961" *) { 1'b1, in_wt_data91[1:0], in_wt_data90 } : { in_wt_data91[1:0], in_wt_data90, 1'b0 };
  assign in_wt_data_fp16_mts_ori45 = cfg_is_fp16_d1[45] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2961" *) _06361_[10:0] : 11'b00000000000;
  assign _06362_[10:0] = in_wt_norm[44] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2970" *) { 1'b1, in_wt_data89[1:0], in_wt_data88 } : { in_wt_data89[1:0], in_wt_data88, 1'b0 };
  assign in_wt_data_fp16_mts_ori44 = cfg_is_fp16_d1[44] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2970" *) _06362_[10:0] : 11'b00000000000;
  assign _06363_[10:0] = in_wt_norm[43] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2979" *) { 1'b1, in_wt_data87[1:0], in_wt_data86 } : { in_wt_data87[1:0], in_wt_data86, 1'b0 };
  assign in_wt_data_fp16_mts_ori43 = cfg_is_fp16_d1[43] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2979" *) _06363_[10:0] : 11'b00000000000;
  assign _06364_[10:0] = in_wt_norm[42] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2988" *) { 1'b1, in_wt_data85[1:0], in_wt_data84 } : { in_wt_data85[1:0], in_wt_data84, 1'b0 };
  assign in_wt_data_fp16_mts_ori42 = cfg_is_fp16_d1[42] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2988" *) _06364_[10:0] : 11'b00000000000;
  assign _06365_[10:0] = in_wt_norm[41] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2997" *) { 1'b1, in_wt_data83[1:0], in_wt_data82 } : { in_wt_data83[1:0], in_wt_data82, 1'b0 };
  assign in_wt_data_fp16_mts_ori41 = cfg_is_fp16_d1[41] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:2997" *) _06365_[10:0] : 11'b00000000000;
  assign _06366_[10:0] = in_wt_norm[40] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3006" *) { 1'b1, in_wt_data81[1:0], in_wt_data80 } : { in_wt_data81[1:0], in_wt_data80, 1'b0 };
  assign in_wt_data_fp16_mts_ori40 = cfg_is_fp16_d1[40] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3006" *) _06366_[10:0] : 11'b00000000000;
  assign _06367_[10:0] = in_wt_norm[39] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3015" *) { 1'b1, in_wt_data79[1:0], in_wt_data78 } : { in_wt_data79[1:0], in_wt_data78, 1'b0 };
  assign in_wt_data_fp16_mts_ori39 = cfg_is_fp16_d1[39] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3015" *) _06367_[10:0] : 11'b00000000000;
  assign _06368_[10:0] = in_wt_norm[38] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3024" *) { 1'b1, in_wt_data77[1:0], in_wt_data76 } : { in_wt_data77[1:0], in_wt_data76, 1'b0 };
  assign in_wt_data_fp16_mts_ori38 = cfg_is_fp16_d1[38] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3024" *) _06368_[10:0] : 11'b00000000000;
  assign _06369_[10:0] = in_wt_norm[37] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3033" *) { 1'b1, in_wt_data75[1:0], in_wt_data74 } : { in_wt_data75[1:0], in_wt_data74, 1'b0 };
  assign in_wt_data_fp16_mts_ori37 = cfg_is_fp16_d1[37] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3033" *) _06369_[10:0] : 11'b00000000000;
  assign _06370_[10:0] = in_wt_norm[36] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3042" *) { 1'b1, in_wt_data73[1:0], in_wt_data72 } : { in_wt_data73[1:0], in_wt_data72, 1'b0 };
  assign in_wt_data_fp16_mts_ori36 = cfg_is_fp16_d1[36] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3042" *) _06370_[10:0] : 11'b00000000000;
  assign _06371_[10:0] = in_wt_norm[35] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3051" *) { 1'b1, in_wt_data71[1:0], in_wt_data70 } : { in_wt_data71[1:0], in_wt_data70, 1'b0 };
  assign in_wt_data_fp16_mts_ori35 = cfg_is_fp16_d1[35] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3051" *) _06371_[10:0] : 11'b00000000000;
  assign _06372_[10:0] = in_wt_norm[34] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3060" *) { 1'b1, in_wt_data69[1:0], in_wt_data68 } : { in_wt_data69[1:0], in_wt_data68, 1'b0 };
  assign in_wt_data_fp16_mts_ori34 = cfg_is_fp16_d1[34] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3060" *) _06372_[10:0] : 11'b00000000000;
  assign _06373_[10:0] = in_wt_norm[33] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3069" *) { 1'b1, in_wt_data67[1:0], in_wt_data66 } : { in_wt_data67[1:0], in_wt_data66, 1'b0 };
  assign in_wt_data_fp16_mts_ori33 = cfg_is_fp16_d1[33] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3069" *) _06373_[10:0] : 11'b00000000000;
  assign _06374_[10:0] = in_wt_norm[32] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3078" *) { 1'b1, in_wt_data65[1:0], in_wt_data64 } : { in_wt_data65[1:0], in_wt_data64, 1'b0 };
  assign in_wt_data_fp16_mts_ori32 = cfg_is_fp16_d1[32] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3078" *) _06374_[10:0] : 11'b00000000000;
  assign _06375_[10:0] = in_wt_norm[31] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3087" *) { 1'b1, in_wt_data63[1:0], in_wt_data62 } : { in_wt_data63[1:0], in_wt_data62, 1'b0 };
  assign in_wt_data_fp16_mts_ori31 = cfg_is_fp16_d1[31] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3087" *) _06375_[10:0] : 11'b00000000000;
  assign _06376_[10:0] = in_wt_norm[30] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3096" *) { 1'b1, in_wt_data61[1:0], in_wt_data60 } : { in_wt_data61[1:0], in_wt_data60, 1'b0 };
  assign in_wt_data_fp16_mts_ori30 = cfg_is_fp16_d1[30] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3096" *) _06376_[10:0] : 11'b00000000000;
  assign _06377_[10:0] = in_wt_norm[29] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3105" *) { 1'b1, in_wt_data59[1:0], in_wt_data58 } : { in_wt_data59[1:0], in_wt_data58, 1'b0 };
  assign in_wt_data_fp16_mts_ori29 = cfg_is_fp16_d1[29] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3105" *) _06377_[10:0] : 11'b00000000000;
  assign _06378_[10:0] = in_wt_norm[28] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3114" *) { 1'b1, in_wt_data57[1:0], in_wt_data56 } : { in_wt_data57[1:0], in_wt_data56, 1'b0 };
  assign in_wt_data_fp16_mts_ori28 = cfg_is_fp16_d1[28] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3114" *) _06378_[10:0] : 11'b00000000000;
  assign _06379_[10:0] = in_wt_norm[27] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3123" *) { 1'b1, in_wt_data55[1:0], in_wt_data54 } : { in_wt_data55[1:0], in_wt_data54, 1'b0 };
  assign in_wt_data_fp16_mts_ori27 = cfg_is_fp16_d1[27] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3123" *) _06379_[10:0] : 11'b00000000000;
  assign _06380_[10:0] = in_wt_norm[26] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3132" *) { 1'b1, in_wt_data53[1:0], in_wt_data52 } : { in_wt_data53[1:0], in_wt_data52, 1'b0 };
  assign in_wt_data_fp16_mts_ori26 = cfg_is_fp16_d1[26] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3132" *) _06380_[10:0] : 11'b00000000000;
  assign _06381_[10:0] = in_wt_norm[25] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3141" *) { 1'b1, in_wt_data51[1:0], in_wt_data50 } : { in_wt_data51[1:0], in_wt_data50, 1'b0 };
  assign in_wt_data_fp16_mts_ori25 = cfg_is_fp16_d1[25] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3141" *) _06381_[10:0] : 11'b00000000000;
  assign _06382_[10:0] = in_wt_norm[24] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3150" *) { 1'b1, in_wt_data49[1:0], in_wt_data48 } : { in_wt_data49[1:0], in_wt_data48, 1'b0 };
  assign in_wt_data_fp16_mts_ori24 = cfg_is_fp16_d1[24] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3150" *) _06382_[10:0] : 11'b00000000000;
  assign _06383_[10:0] = in_wt_norm[23] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3159" *) { 1'b1, in_wt_data47[1:0], in_wt_data46 } : { in_wt_data47[1:0], in_wt_data46, 1'b0 };
  assign in_wt_data_fp16_mts_ori23 = cfg_is_fp16_d1[23] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3159" *) _06383_[10:0] : 11'b00000000000;
  assign _06384_[10:0] = in_wt_norm[22] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3168" *) { 1'b1, in_wt_data45[1:0], in_wt_data44 } : { in_wt_data45[1:0], in_wt_data44, 1'b0 };
  assign in_wt_data_fp16_mts_ori22 = cfg_is_fp16_d1[22] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3168" *) _06384_[10:0] : 11'b00000000000;
  assign _06385_[10:0] = in_wt_norm[21] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3177" *) { 1'b1, in_wt_data43[1:0], in_wt_data42 } : { in_wt_data43[1:0], in_wt_data42, 1'b0 };
  assign in_wt_data_fp16_mts_ori21 = cfg_is_fp16_d1[21] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3177" *) _06385_[10:0] : 11'b00000000000;
  assign _06386_[10:0] = in_wt_norm[20] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3186" *) { 1'b1, in_wt_data41[1:0], in_wt_data40 } : { in_wt_data41[1:0], in_wt_data40, 1'b0 };
  assign in_wt_data_fp16_mts_ori20 = cfg_is_fp16_d1[20] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3186" *) _06386_[10:0] : 11'b00000000000;
  assign _06387_[10:0] = in_wt_norm[19] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3195" *) { 1'b1, in_wt_data39[1:0], in_wt_data38 } : { in_wt_data39[1:0], in_wt_data38, 1'b0 };
  assign in_wt_data_fp16_mts_ori19 = cfg_is_fp16_d1[19] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3195" *) _06387_[10:0] : 11'b00000000000;
  assign _06388_[10:0] = in_wt_norm[18] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3204" *) { 1'b1, in_wt_data37[1:0], in_wt_data36 } : { in_wt_data37[1:0], in_wt_data36, 1'b0 };
  assign in_wt_data_fp16_mts_ori18 = cfg_is_fp16_d1[18] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3204" *) _06388_[10:0] : 11'b00000000000;
  assign _06389_[10:0] = in_wt_norm[17] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3213" *) { 1'b1, in_wt_data35[1:0], in_wt_data34 } : { in_wt_data35[1:0], in_wt_data34, 1'b0 };
  assign in_wt_data_fp16_mts_ori17 = cfg_is_fp16_d1[17] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3213" *) _06389_[10:0] : 11'b00000000000;
  assign _06390_[10:0] = in_wt_norm[16] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3222" *) { 1'b1, in_wt_data33[1:0], in_wt_data32 } : { in_wt_data33[1:0], in_wt_data32, 1'b0 };
  assign in_wt_data_fp16_mts_ori16 = cfg_is_fp16_d1[16] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3222" *) _06390_[10:0] : 11'b00000000000;
  assign _06391_[10:0] = in_wt_norm[15] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3231" *) { 1'b1, in_wt_data31[1:0], in_wt_data30 } : { in_wt_data31[1:0], in_wt_data30, 1'b0 };
  assign in_wt_data_fp16_mts_ori15 = cfg_is_fp16_d1[15] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3231" *) _06391_[10:0] : 11'b00000000000;
  assign _06392_[10:0] = in_wt_norm[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3240" *) { 1'b1, in_wt_data29[1:0], in_wt_data28 } : { in_wt_data29[1:0], in_wt_data28, 1'b0 };
  assign in_wt_data_fp16_mts_ori14 = cfg_is_fp16_d1[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3240" *) _06392_[10:0] : 11'b00000000000;
  assign _06393_[10:0] = in_wt_norm[13] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3249" *) { 1'b1, in_wt_data27[1:0], in_wt_data26 } : { in_wt_data27[1:0], in_wt_data26, 1'b0 };
  assign in_wt_data_fp16_mts_ori13 = cfg_is_fp16_d1[13] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3249" *) _06393_[10:0] : 11'b00000000000;
  assign _06394_[10:0] = in_wt_norm[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3258" *) { 1'b1, in_wt_data25[1:0], in_wt_data24 } : { in_wt_data25[1:0], in_wt_data24, 1'b0 };
  assign in_wt_data_fp16_mts_ori12 = cfg_is_fp16_d1[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3258" *) _06394_[10:0] : 11'b00000000000;
  assign _06395_[10:0] = in_wt_norm[11] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3267" *) { 1'b1, in_wt_data23[1:0], in_wt_data22 } : { in_wt_data23[1:0], in_wt_data22, 1'b0 };
  assign in_wt_data_fp16_mts_ori11 = cfg_is_fp16_d1[11] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3267" *) _06395_[10:0] : 11'b00000000000;
  assign _06396_[10:0] = in_wt_norm[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3276" *) { 1'b1, in_wt_data21[1:0], in_wt_data20 } : { in_wt_data21[1:0], in_wt_data20, 1'b0 };
  assign in_wt_data_fp16_mts_ori10 = cfg_is_fp16_d1[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3276" *) _06396_[10:0] : 11'b00000000000;
  assign _06397_[10:0] = in_wt_norm[9] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3285" *) { 1'b1, in_wt_data19[1:0], in_wt_data18 } : { in_wt_data19[1:0], in_wt_data18, 1'b0 };
  assign in_wt_data_fp16_mts_ori9 = cfg_is_fp16_d1[9] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3285" *) _06397_[10:0] : 11'b00000000000;
  assign _06398_[10:0] = in_wt_norm[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3294" *) { 1'b1, in_wt_data17[1:0], in_wt_data16 } : { in_wt_data17[1:0], in_wt_data16, 1'b0 };
  assign in_wt_data_fp16_mts_ori8 = cfg_is_fp16_d1[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3294" *) _06398_[10:0] : 11'b00000000000;
  assign _06399_[10:0] = in_wt_norm[7] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3303" *) { 1'b1, in_wt_data15[1:0], in_wt_data14 } : { in_wt_data15[1:0], in_wt_data14, 1'b0 };
  assign in_wt_data_fp16_mts_ori7 = cfg_is_fp16_d1[7] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3303" *) _06399_[10:0] : 11'b00000000000;
  assign _06400_[10:0] = in_wt_norm[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3312" *) { 1'b1, in_wt_data13[1:0], in_wt_data12 } : { in_wt_data13[1:0], in_wt_data12, 1'b0 };
  assign in_wt_data_fp16_mts_ori6 = cfg_is_fp16_d1[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3312" *) _06400_[10:0] : 11'b00000000000;
  assign _06401_[10:0] = in_wt_norm[5] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3321" *) { 1'b1, in_wt_data11[1:0], in_wt_data10 } : { in_wt_data11[1:0], in_wt_data10, 1'b0 };
  assign in_wt_data_fp16_mts_ori5 = cfg_is_fp16_d1[5] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3321" *) _06401_[10:0] : 11'b00000000000;
  assign _06402_[10:0] = in_wt_norm[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3330" *) { 1'b1, in_wt_data9[1:0], in_wt_data8 } : { in_wt_data9[1:0], in_wt_data8, 1'b0 };
  assign in_wt_data_fp16_mts_ori4 = cfg_is_fp16_d1[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3330" *) _06402_[10:0] : 11'b00000000000;
  assign _06403_[10:0] = in_wt_norm[3] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3339" *) { 1'b1, in_wt_data7[1:0], in_wt_data6 } : { in_wt_data7[1:0], in_wt_data6, 1'b0 };
  assign in_wt_data_fp16_mts_ori3 = cfg_is_fp16_d1[3] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3339" *) _06403_[10:0] : 11'b00000000000;
  assign _06404_[10:0] = in_wt_norm[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3348" *) { 1'b1, in_wt_data5[1:0], in_wt_data4 } : { in_wt_data5[1:0], in_wt_data4, 1'b0 };
  assign in_wt_data_fp16_mts_ori2 = cfg_is_fp16_d1[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3348" *) _06404_[10:0] : 11'b00000000000;
  assign _06405_[10:0] = in_wt_norm[1] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3357" *) { 1'b1, in_wt_data3[1:0], in_wt_data2 } : { in_wt_data3[1:0], in_wt_data2, 1'b0 };
  assign in_wt_data_fp16_mts_ori1 = cfg_is_fp16_d1[1] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3357" *) _06405_[10:0] : 11'b00000000000;
  assign _06406_[10:0] = in_wt_norm[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3366" *) { 1'b1, in_wt_data1[1:0], in_wt_data0 } : { in_wt_data1[1:0], in_wt_data0, 1'b0 };
  assign in_wt_data_fp16_mts_ori0 = cfg_is_fp16_d1[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3366" *) _06406_[10:0] : 11'b00000000000;
  assign _08344_[126:0] = cfg_is_int8_d1[64] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3970" *) { in_wt_mask[63], in_wt_mask[126], in_wt_mask[62], in_wt_mask[125], in_wt_mask[61], in_wt_mask[124], in_wt_mask[60], in_wt_mask[123], in_wt_mask[59], in_wt_mask[122], in_wt_mask[58], in_wt_mask[121], in_wt_mask[57], in_wt_mask[120], in_wt_mask[56], in_wt_mask[119], in_wt_mask[55], in_wt_mask[118], in_wt_mask[54], in_wt_mask[117], in_wt_mask[53], in_wt_mask[116], in_wt_mask[52], in_wt_mask[115], in_wt_mask[51], in_wt_mask[114], in_wt_mask[50], in_wt_mask[113], in_wt_mask[49], in_wt_mask[112], in_wt_mask[48], in_wt_mask[111], in_wt_mask[47], in_wt_mask[110], in_wt_mask[46], in_wt_mask[109], in_wt_mask[45], in_wt_mask[108], in_wt_mask[44], in_wt_mask[107], in_wt_mask[43], in_wt_mask[106], in_wt_mask[42], in_wt_mask[105], in_wt_mask[41], in_wt_mask[104], in_wt_mask[40], in_wt_mask[103], in_wt_mask[39], in_wt_mask[102], in_wt_mask[38], in_wt_mask[101], in_wt_mask[37], in_wt_mask[100], in_wt_mask[36], in_wt_mask[99], in_wt_mask[35], in_wt_mask[98], in_wt_mask[34], in_wt_mask[97], in_wt_mask[33], in_wt_mask[96], in_wt_mask[32], in_wt_mask[95], in_wt_mask[31], in_wt_mask[94], in_wt_mask[30], in_wt_mask[93], in_wt_mask[29], in_wt_mask[92], in_wt_mask[28], in_wt_mask[91], in_wt_mask[27], in_wt_mask[90], in_wt_mask[26], in_wt_mask[89], in_wt_mask[25], in_wt_mask[88], in_wt_mask[24], in_wt_mask[87], in_wt_mask[23], in_wt_mask[86], in_wt_mask[22], in_wt_mask[85], in_wt_mask[21], in_wt_mask[84], in_wt_mask[20], in_wt_mask[83], in_wt_mask[19], in_wt_mask[82], in_wt_mask[18], in_wt_mask[81], in_wt_mask[17], in_wt_mask[80], in_wt_mask[16], in_wt_mask[79], in_wt_mask[15], in_wt_mask[78], in_wt_mask[14], in_wt_mask[77], in_wt_mask[13], in_wt_mask[76], in_wt_mask[12], in_wt_mask[75], in_wt_mask[11], in_wt_mask[74], in_wt_mask[10], in_wt_mask[73], in_wt_mask[9], in_wt_mask[72], in_wt_mask[8], in_wt_mask[71], in_wt_mask[7], in_wt_mask[70], in_wt_mask[6], in_wt_mask[69], in_wt_mask[5], in_wt_mask[68], in_wt_mask[4], in_wt_mask[67], in_wt_mask[3], in_wt_mask[66], in_wt_mask[2], in_wt_mask[65], in_wt_mask[1], in_wt_mask[64], in_wt_mask[0] } : in_wt_mask[126:0];
  assign wt_pre_nz_w = cfg_is_fp16_d1[64] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:3970" *) _05698_ : { in_wt_mask[127], _08344_[126:0] };
  assign _08345_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5322" *) 1'b0 : wt0_sd_pvld;
  assign wt0_sd_pvld_w = wt_pre_sel[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:5322" *) 1'b1 : _08345_;
  assign _08346_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6658" *) 1'b0 : wt1_sd_pvld;
  assign wt1_sd_pvld_w = wt_pre_sel[1] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:6658" *) 1'b1 : _08346_;
  assign _08347_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7994" *) 1'b0 : wt2_sd_pvld;
  assign wt2_sd_pvld_w = wt_pre_sel[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:7994" *) 1'b1 : _08347_;
  assign _08348_ = dat_pre_stripe_st[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9330" *) 1'b0 : wt3_sd_pvld;
  assign wt3_sd_pvld_w = wt_pre_sel[3] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_active.v:9330" *) 1'b1 : _08348_;
  assign _01189_[7:0] = { _01189_[8], _01189_[8], _01189_[8], _01189_[8], _01189_[8], _01189_[8], _01189_[8], _01189_[8] };
  assign _01190_[14:0] = { _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15], _01190_[15] };
  assign _06279_[11] = 1'b0;
  assign _06280_[11] = 1'b0;
  assign _06281_[11] = 1'b0;
  assign _06282_[11] = 1'b0;
  assign _06283_[11] = 1'b0;
  assign _06284_[11] = 1'b0;
  assign _06285_[11] = 1'b0;
  assign _06286_[11] = 1'b0;
  assign _06287_[11] = 1'b0;
  assign _06288_[11] = 1'b0;
  assign _06289_[11] = 1'b0;
  assign _06290_[11] = 1'b0;
  assign _06291_[11] = 1'b0;
  assign _06292_[11] = 1'b0;
  assign _06293_[11] = 1'b0;
  assign _06294_[11] = 1'b0;
  assign _06295_[11] = 1'b0;
  assign _06296_[11] = 1'b0;
  assign _06297_[11] = 1'b0;
  assign _06298_[11] = 1'b0;
  assign _06299_[11] = 1'b0;
  assign _06300_[11] = 1'b0;
  assign _06301_[11] = 1'b0;
  assign _06302_[11] = 1'b0;
  assign _06303_[11] = 1'b0;
  assign _06304_[11] = 1'b0;
  assign _06305_[11] = 1'b0;
  assign _06306_[11] = 1'b0;
  assign _06307_[11] = 1'b0;
  assign _06308_[11] = 1'b0;
  assign _06309_[11] = 1'b0;
  assign _06310_[11] = 1'b0;
  assign _06311_[11] = 1'b0;
  assign _06312_[11] = 1'b0;
  assign _06313_[11] = 1'b0;
  assign _06314_[11] = 1'b0;
  assign _06315_[11] = 1'b0;
  assign _06316_[11] = 1'b0;
  assign _06317_[11] = 1'b0;
  assign _06318_[11] = 1'b0;
  assign _06319_[11] = 1'b0;
  assign _06320_[11] = 1'b0;
  assign _06321_[11] = 1'b0;
  assign _06322_[11] = 1'b0;
  assign _06323_[11] = 1'b0;
  assign _06324_[11] = 1'b0;
  assign _06325_[11] = 1'b0;
  assign _06326_[11] = 1'b0;
  assign _06327_[11] = 1'b0;
  assign _06328_[11] = 1'b0;
  assign _06329_[11] = 1'b0;
  assign _06330_[11] = 1'b0;
  assign _06331_[11] = 1'b0;
  assign _06332_[11] = 1'b0;
  assign _06333_[11] = 1'b0;
  assign _06334_[11] = 1'b0;
  assign _06335_[11] = 1'b0;
  assign _06336_[11] = 1'b0;
  assign _06337_[11] = 1'b0;
  assign _06338_[11] = 1'b0;
  assign _06339_[11] = 1'b0;
  assign _06340_[11] = 1'b0;
  assign _06341_[11] = 1'b0;
  assign _06342_[11] = 1'b0;
  assign _06343_[11] = 1'b0;
  assign _06344_[11] = 1'b0;
  assign _06345_[11] = 1'b0;
  assign _06346_[11] = 1'b0;
  assign _06347_[11] = 1'b0;
  assign _06348_[11] = 1'b0;
  assign _06349_[11] = 1'b0;
  assign _06350_[11] = 1'b0;
  assign _06351_[11] = 1'b0;
  assign _06352_[11] = 1'b0;
  assign _06353_[11] = 1'b0;
  assign _06354_[11] = 1'b0;
  assign _06355_[11] = 1'b0;
  assign _06356_[11] = 1'b0;
  assign _06357_[11] = 1'b0;
  assign _06358_[11] = 1'b0;
  assign _06359_[11] = 1'b0;
  assign _06360_[11] = 1'b0;
  assign _06361_[11] = 1'b0;
  assign _06362_[11] = 1'b0;
  assign _06363_[11] = 1'b0;
  assign _06364_[11] = 1'b0;
  assign _06365_[11] = 1'b0;
  assign _06366_[11] = 1'b0;
  assign _06367_[11] = 1'b0;
  assign _06368_[11] = 1'b0;
  assign _06369_[11] = 1'b0;
  assign _06370_[11] = 1'b0;
  assign _06371_[11] = 1'b0;
  assign _06372_[11] = 1'b0;
  assign _06373_[11] = 1'b0;
  assign _06374_[11] = 1'b0;
  assign _06375_[11] = 1'b0;
  assign _06376_[11] = 1'b0;
  assign _06377_[11] = 1'b0;
  assign _06378_[11] = 1'b0;
  assign _06379_[11] = 1'b0;
  assign _06380_[11] = 1'b0;
  assign _06381_[11] = 1'b0;
  assign _06382_[11] = 1'b0;
  assign _06383_[11] = 1'b0;
  assign _06384_[11] = 1'b0;
  assign _06385_[11] = 1'b0;
  assign _06386_[11] = 1'b0;
  assign _06387_[11] = 1'b0;
  assign _06388_[11] = 1'b0;
  assign _06389_[11] = 1'b0;
  assign _06390_[11] = 1'b0;
  assign _06391_[11] = 1'b0;
  assign _06392_[11] = 1'b0;
  assign _06393_[11] = 1'b0;
  assign _06394_[11] = 1'b0;
  assign _06395_[11] = 1'b0;
  assign _06396_[11] = 1'b0;
  assign _06397_[11] = 1'b0;
  assign _06398_[11] = 1'b0;
  assign _06399_[11] = 1'b0;
  assign _06400_[11] = 1'b0;
  assign _06401_[11] = 1'b0;
  assign _06402_[11] = 1'b0;
  assign _06403_[11] = 1'b0;
  assign _06404_[11] = 1'b0;
  assign _06405_[11] = 1'b0;
  assign _06406_[11] = 1'b0;
  assign _08343_[127] = in_dat_mask[127];
  assign _08344_[127] = in_wt_mask[127];
  assign dat0_actv_data = dat_actv_data_reg0;
  assign dat0_actv_nan = dat_actv_nan_reg0;
  assign dat0_actv_nz = dat_actv_nz_reg0;
  assign dat0_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat0_pre_exp = dat_pre_exp_reg0;
  assign dat0_pre_mask = dat_pre_mask0;
  assign dat0_pre_pvld = dat_pre_pvld[0];
  assign dat0_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat0_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat1_actv_data = dat_actv_data_reg1;
  assign dat1_actv_nan = dat_actv_nan_reg1;
  assign dat1_actv_nz = dat_actv_nz_reg1;
  assign dat1_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat1_pre_exp = dat_pre_exp_reg1;
  assign dat1_pre_mask = dat_pre_mask1;
  assign dat1_pre_pvld = dat_pre_pvld[0];
  assign dat1_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat1_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat2_actv_data = dat_actv_data_reg2;
  assign dat2_actv_nan = dat_actv_nan_reg2;
  assign dat2_actv_nz = dat_actv_nz_reg2;
  assign dat2_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat2_pre_exp = dat_pre_exp_reg2;
  assign dat2_pre_mask = dat_pre_mask2;
  assign dat2_pre_pvld = dat_pre_pvld[0];
  assign dat2_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat2_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat3_actv_data = dat_actv_data_reg3;
  assign dat3_actv_nan = dat_actv_nan_reg3;
  assign dat3_actv_nz = dat_actv_nz_reg3;
  assign dat3_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat3_pre_exp = dat_pre_exp_reg3;
  assign dat3_pre_mask = dat_pre_mask3;
  assign dat3_pre_pvld = dat_pre_pvld[0];
  assign dat3_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat3_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat4_actv_data = dat_actv_data_reg4;
  assign dat4_actv_nan = dat_actv_nan_reg4;
  assign dat4_actv_nz = dat_actv_nz_reg4;
  assign dat4_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat4_pre_exp = dat_pre_exp_reg4;
  assign dat4_pre_mask = dat_pre_mask4;
  assign dat4_pre_pvld = dat_pre_pvld[0];
  assign dat4_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat4_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat5_actv_data = dat_actv_data_reg5;
  assign dat5_actv_nan = dat_actv_nan_reg5;
  assign dat5_actv_nz = dat_actv_nz_reg5;
  assign dat5_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat5_pre_exp = dat_pre_exp_reg5;
  assign dat5_pre_mask = dat_pre_mask5;
  assign dat5_pre_pvld = dat_pre_pvld[0];
  assign dat5_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat5_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat6_actv_data = dat_actv_data_reg6;
  assign dat6_actv_nan = dat_actv_nan_reg6;
  assign dat6_actv_nz = dat_actv_nz_reg6;
  assign dat6_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat6_pre_exp = dat_pre_exp_reg6;
  assign dat6_pre_mask = dat_pre_mask6;
  assign dat6_pre_pvld = dat_pre_pvld[0];
  assign dat6_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat6_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat7_actv_data = dat_actv_data_reg7;
  assign dat7_actv_nan = dat_actv_nan_reg7;
  assign dat7_actv_nz = dat_actv_nz_reg7;
  assign dat7_actv_pvld = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat7_pre_exp = dat_pre_exp_reg7;
  assign dat7_pre_mask = dat_pre_mask7;
  assign dat7_pre_pvld = dat_pre_pvld[0];
  assign dat7_pre_stripe_end = dat_pre_stripe_end[0];
  assign dat7_pre_stripe_st = dat_pre_stripe_st[0];
  assign dat_actv_pvld_reg0 = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_actv_pvld_reg1 = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_actv_pvld_reg2 = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_actv_pvld_reg3 = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_actv_pvld_reg4 = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_actv_pvld_reg5 = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_actv_pvld_reg6 = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_actv_pvld_reg7[103:1] = { dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0], dat_actv_pvld_reg7[0] };
  assign dat_pre_mask_w = { dat_pre_nz_w[126], dat_pre_nz_w[124], dat_pre_nz_w[122], dat_pre_nz_w[120], dat_pre_nz_w[118], dat_pre_nz_w[116], dat_pre_nz_w[114], dat_pre_nz_w[112], dat_pre_nz_w[110], dat_pre_nz_w[108], dat_pre_nz_w[106], dat_pre_nz_w[104], dat_pre_nz_w[102], dat_pre_nz_w[100], dat_pre_nz_w[98], dat_pre_nz_w[96], dat_pre_nz_w[94], dat_pre_nz_w[92], dat_pre_nz_w[90], dat_pre_nz_w[88], dat_pre_nz_w[86], dat_pre_nz_w[84], dat_pre_nz_w[82], dat_pre_nz_w[80], dat_pre_nz_w[78], dat_pre_nz_w[76], dat_pre_nz_w[74], dat_pre_nz_w[72], dat_pre_nz_w[70], dat_pre_nz_w[68], dat_pre_nz_w[66], dat_pre_nz_w[64], dat_pre_nz_w[62], dat_pre_nz_w[60], dat_pre_nz_w[58], dat_pre_nz_w[56], dat_pre_nz_w[54], dat_pre_nz_w[52], dat_pre_nz_w[50], dat_pre_nz_w[48], dat_pre_nz_w[46], dat_pre_nz_w[44], dat_pre_nz_w[42], dat_pre_nz_w[40], dat_pre_nz_w[38], dat_pre_nz_w[36], dat_pre_nz_w[34], dat_pre_nz_w[32], dat_pre_nz_w[30], dat_pre_nz_w[28], dat_pre_nz_w[26], dat_pre_nz_w[24], dat_pre_nz_w[22], dat_pre_nz_w[20], dat_pre_nz_w[18], dat_pre_nz_w[16], dat_pre_nz_w[14], dat_pre_nz_w[12], dat_pre_nz_w[10], dat_pre_nz_w[8], dat_pre_nz_w[6], dat_pre_nz_w[4], dat_pre_nz_w[2], dat_pre_nz_w[0] };
  assign dat_pre_pvld[15:1] = { dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0], dat_pre_pvld[0] };
  assign dat_pre_stripe_end[8:1] = { dat_pre_stripe_end[0], dat_pre_stripe_end[0], dat_pre_stripe_end[0], dat_pre_stripe_end[0], dat_pre_stripe_end[0], dat_pre_stripe_end[0], dat_pre_stripe_end[0], dat_pre_stripe_end[0] };
  assign dat_pre_stripe_st[15:1] = { dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0], dat_pre_stripe_st[0] };
  assign in_dat_data_fp16 = { in_dat_data_fp16_63, in_dat_data_fp16_62, in_dat_data_fp16_61, in_dat_data_fp16_60, in_dat_data_fp16_59, in_dat_data_fp16_58, in_dat_data_fp16_57, in_dat_data_fp16_56, in_dat_data_fp16_55, in_dat_data_fp16_54, in_dat_data_fp16_53, in_dat_data_fp16_52, in_dat_data_fp16_51, in_dat_data_fp16_50, in_dat_data_fp16_49, in_dat_data_fp16_48, in_dat_data_fp16_47, in_dat_data_fp16_46, in_dat_data_fp16_45, in_dat_data_fp16_44, in_dat_data_fp16_43, in_dat_data_fp16_42, in_dat_data_fp16_41, in_dat_data_fp16_40, in_dat_data_fp16_39, in_dat_data_fp16_38, in_dat_data_fp16_37, in_dat_data_fp16_36, in_dat_data_fp16_35, in_dat_data_fp16_34, in_dat_data_fp16_33, in_dat_data_fp16_32, in_dat_data_fp16_31, in_dat_data_fp16_30, in_dat_data_fp16_29, in_dat_data_fp16_28, in_dat_data_fp16_27, in_dat_data_fp16_26, in_dat_data_fp16_25, in_dat_data_fp16_24, in_dat_data_fp16_23, in_dat_data_fp16_22, in_dat_data_fp16_21, in_dat_data_fp16_20, in_dat_data_fp16_19, in_dat_data_fp16_18, in_dat_data_fp16_17, in_dat_data_fp16_16, in_dat_data_fp16_15, in_dat_data_fp16_14, in_dat_data_fp16_13, in_dat_data_fp16_12, in_dat_data_fp16_11, in_dat_data_fp16_10, in_dat_data_fp16_9, in_dat_data_fp16_8, in_dat_data_fp16_7, in_dat_data_fp16_6, in_dat_data_fp16_5, in_dat_data_fp16_4, in_dat_data_fp16_3, in_dat_data_fp16_2, in_dat_data_fp16_1, in_dat_data_fp16_0 };
  assign in_dat_data_int16 = { in_dat_data_int16_63, in_dat_data_int16_62, in_dat_data_int16_61, in_dat_data_int16_60, in_dat_data_int16_59, in_dat_data_int16_58, in_dat_data_int16_57, in_dat_data_int16_56, in_dat_data_int16_55, in_dat_data_int16_54, in_dat_data_int16_53, in_dat_data_int16_52, in_dat_data_int16_51, in_dat_data_int16_50, in_dat_data_int16_49, in_dat_data_int16_48, in_dat_data_int16_47, in_dat_data_int16_46, in_dat_data_int16_45, in_dat_data_int16_44, in_dat_data_int16_43, in_dat_data_int16_42, in_dat_data_int16_41, in_dat_data_int16_40, in_dat_data_int16_39, in_dat_data_int16_38, in_dat_data_int16_37, in_dat_data_int16_36, in_dat_data_int16_35, in_dat_data_int16_34, in_dat_data_int16_33, in_dat_data_int16_32, in_dat_data_int16_31, in_dat_data_int16_30, in_dat_data_int16_29, in_dat_data_int16_28, in_dat_data_int16_27, in_dat_data_int16_26, in_dat_data_int16_25, in_dat_data_int16_24, in_dat_data_int16_23, in_dat_data_int16_22, in_dat_data_int16_21, in_dat_data_int16_20, in_dat_data_int16_19, in_dat_data_int16_18, in_dat_data_int16_17, in_dat_data_int16_16, in_dat_data_int16_15, in_dat_data_int16_14, in_dat_data_int16_13, in_dat_data_int16_12, in_dat_data_int16_11, in_dat_data_int16_10, in_dat_data_int16_9, in_dat_data_int16_8, in_dat_data_int16_7, in_dat_data_int16_6, in_dat_data_int16_5, in_dat_data_int16_4, in_dat_data_int16_3, in_dat_data_int16_2, in_dat_data_int16_1, in_dat_data_int16_0 };
  assign in_dat_data_int8 = { in_dat_data_int8_63, in_dat_data_int8_62, in_dat_data_int8_61, in_dat_data_int8_60, in_dat_data_int8_59, in_dat_data_int8_58, in_dat_data_int8_57, in_dat_data_int8_56, in_dat_data_int8_55, in_dat_data_int8_54, in_dat_data_int8_53, in_dat_data_int8_52, in_dat_data_int8_51, in_dat_data_int8_50, in_dat_data_int8_49, in_dat_data_int8_48, in_dat_data_int8_47, in_dat_data_int8_46, in_dat_data_int8_45, in_dat_data_int8_44, in_dat_data_int8_43, in_dat_data_int8_42, in_dat_data_int8_41, in_dat_data_int8_40, in_dat_data_int8_39, in_dat_data_int8_38, in_dat_data_int8_37, in_dat_data_int8_36, in_dat_data_int8_35, in_dat_data_int8_34, in_dat_data_int8_33, in_dat_data_int8_32, in_dat_data_int8_31, in_dat_data_int8_30, in_dat_data_int8_29, in_dat_data_int8_28, in_dat_data_int8_27, in_dat_data_int8_26, in_dat_data_int8_25, in_dat_data_int8_24, in_dat_data_int8_23, in_dat_data_int8_22, in_dat_data_int8_21, in_dat_data_int8_20, in_dat_data_int8_19, in_dat_data_int8_18, in_dat_data_int8_17, in_dat_data_int8_16, in_dat_data_int8_15, in_dat_data_int8_14, in_dat_data_int8_13, in_dat_data_int8_12, in_dat_data_int8_11, in_dat_data_int8_10, in_dat_data_int8_9, in_dat_data_int8_8, in_dat_data_int8_7, in_dat_data_int8_6, in_dat_data_int8_5, in_dat_data_int8_4, in_dat_data_int8_3, in_dat_data_int8_2, in_dat_data_int8_1, in_dat_data_int8_0 };
  assign in_dat_data_pack = { in_dat_data127, in_dat_data126, in_dat_data125, in_dat_data124, in_dat_data123, in_dat_data122, in_dat_data121, in_dat_data120, in_dat_data119, in_dat_data118, in_dat_data117, in_dat_data116, in_dat_data115, in_dat_data114, in_dat_data113, in_dat_data112, in_dat_data111, in_dat_data110, in_dat_data109, in_dat_data108, in_dat_data107, in_dat_data106, in_dat_data105, in_dat_data104, in_dat_data103, in_dat_data102, in_dat_data101, in_dat_data100, in_dat_data99, in_dat_data98, in_dat_data97, in_dat_data96, in_dat_data95, in_dat_data94, in_dat_data93, in_dat_data92, in_dat_data91, in_dat_data90, in_dat_data89, in_dat_data88, in_dat_data87, in_dat_data86, in_dat_data85, in_dat_data84, in_dat_data83, in_dat_data82, in_dat_data81, in_dat_data80, in_dat_data79, in_dat_data78, in_dat_data77, in_dat_data76, in_dat_data75, in_dat_data74, in_dat_data73, in_dat_data72, in_dat_data71, in_dat_data70, in_dat_data69, in_dat_data68, in_dat_data67, in_dat_data66, in_dat_data65, in_dat_data64, in_dat_data63, in_dat_data62, in_dat_data61, in_dat_data60, in_dat_data59, in_dat_data58, in_dat_data57, in_dat_data56, in_dat_data55, in_dat_data54, in_dat_data53, in_dat_data52, in_dat_data51, in_dat_data50, in_dat_data49, in_dat_data48, in_dat_data47, in_dat_data46, in_dat_data45, in_dat_data44, in_dat_data43, in_dat_data42, in_dat_data41, in_dat_data40, in_dat_data39, in_dat_data38, in_dat_data37, in_dat_data36, in_dat_data35, in_dat_data34, in_dat_data33, in_dat_data32, in_dat_data31, in_dat_data30, in_dat_data29, in_dat_data28, in_dat_data27, in_dat_data26, in_dat_data25, in_dat_data24, in_dat_data23, in_dat_data22, in_dat_data21, in_dat_data20, in_dat_data19, in_dat_data18, in_dat_data17, in_dat_data16, in_dat_data15, in_dat_data14, in_dat_data13, in_dat_data12, in_dat_data11, in_dat_data10, in_dat_data9, in_dat_data8, in_dat_data7, in_dat_data6, in_dat_data5, in_dat_data4, in_dat_data3, in_dat_data2, in_dat_data1, in_dat_data0 };
  assign in_dat_exp = dat_pre_exp_w;
  assign in_dat_mask_int8 = { in_dat_mask[127], in_dat_mask[63], in_dat_mask[126], in_dat_mask[62], in_dat_mask[125], in_dat_mask[61], in_dat_mask[124], in_dat_mask[60], in_dat_mask[123], in_dat_mask[59], in_dat_mask[122], in_dat_mask[58], in_dat_mask[121], in_dat_mask[57], in_dat_mask[120], in_dat_mask[56], in_dat_mask[119], in_dat_mask[55], in_dat_mask[118], in_dat_mask[54], in_dat_mask[117], in_dat_mask[53], in_dat_mask[116], in_dat_mask[52], in_dat_mask[115], in_dat_mask[51], in_dat_mask[114], in_dat_mask[50], in_dat_mask[113], in_dat_mask[49], in_dat_mask[112], in_dat_mask[48], in_dat_mask[111], in_dat_mask[47], in_dat_mask[110], in_dat_mask[46], in_dat_mask[109], in_dat_mask[45], in_dat_mask[108], in_dat_mask[44], in_dat_mask[107], in_dat_mask[43], in_dat_mask[106], in_dat_mask[42], in_dat_mask[105], in_dat_mask[41], in_dat_mask[104], in_dat_mask[40], in_dat_mask[103], in_dat_mask[39], in_dat_mask[102], in_dat_mask[38], in_dat_mask[101], in_dat_mask[37], in_dat_mask[100], in_dat_mask[36], in_dat_mask[99], in_dat_mask[35], in_dat_mask[98], in_dat_mask[34], in_dat_mask[97], in_dat_mask[33], in_dat_mask[96], in_dat_mask[32], in_dat_mask[95], in_dat_mask[31], in_dat_mask[94], in_dat_mask[30], in_dat_mask[93], in_dat_mask[29], in_dat_mask[92], in_dat_mask[28], in_dat_mask[91], in_dat_mask[27], in_dat_mask[90], in_dat_mask[26], in_dat_mask[89], in_dat_mask[25], in_dat_mask[88], in_dat_mask[24], in_dat_mask[87], in_dat_mask[23], in_dat_mask[86], in_dat_mask[22], in_dat_mask[85], in_dat_mask[21], in_dat_mask[84], in_dat_mask[20], in_dat_mask[83], in_dat_mask[19], in_dat_mask[82], in_dat_mask[18], in_dat_mask[81], in_dat_mask[17], in_dat_mask[80], in_dat_mask[16], in_dat_mask[79], in_dat_mask[15], in_dat_mask[78], in_dat_mask[14], in_dat_mask[77], in_dat_mask[13], in_dat_mask[76], in_dat_mask[12], in_dat_mask[75], in_dat_mask[11], in_dat_mask[74], in_dat_mask[10], in_dat_mask[73], in_dat_mask[9], in_dat_mask[72], in_dat_mask[8], in_dat_mask[71], in_dat_mask[7], in_dat_mask[70], in_dat_mask[6], in_dat_mask[69], in_dat_mask[5], in_dat_mask[68], in_dat_mask[4], in_dat_mask[67], in_dat_mask[3], in_dat_mask[66], in_dat_mask[2], in_dat_mask[65], in_dat_mask[1], in_dat_mask[64], in_dat_mask[0] };
  assign in_wt_data_fp16 = { in_wt_data_fp16_63, in_wt_data_fp16_62, in_wt_data_fp16_61, in_wt_data_fp16_60, in_wt_data_fp16_59, in_wt_data_fp16_58, in_wt_data_fp16_57, in_wt_data_fp16_56, in_wt_data_fp16_55, in_wt_data_fp16_54, in_wt_data_fp16_53, in_wt_data_fp16_52, in_wt_data_fp16_51, in_wt_data_fp16_50, in_wt_data_fp16_49, in_wt_data_fp16_48, in_wt_data_fp16_47, in_wt_data_fp16_46, in_wt_data_fp16_45, in_wt_data_fp16_44, in_wt_data_fp16_43, in_wt_data_fp16_42, in_wt_data_fp16_41, in_wt_data_fp16_40, in_wt_data_fp16_39, in_wt_data_fp16_38, in_wt_data_fp16_37, in_wt_data_fp16_36, in_wt_data_fp16_35, in_wt_data_fp16_34, in_wt_data_fp16_33, in_wt_data_fp16_32, in_wt_data_fp16_31, in_wt_data_fp16_30, in_wt_data_fp16_29, in_wt_data_fp16_28, in_wt_data_fp16_27, in_wt_data_fp16_26, in_wt_data_fp16_25, in_wt_data_fp16_24, in_wt_data_fp16_23, in_wt_data_fp16_22, in_wt_data_fp16_21, in_wt_data_fp16_20, in_wt_data_fp16_19, in_wt_data_fp16_18, in_wt_data_fp16_17, in_wt_data_fp16_16, in_wt_data_fp16_15, in_wt_data_fp16_14, in_wt_data_fp16_13, in_wt_data_fp16_12, in_wt_data_fp16_11, in_wt_data_fp16_10, in_wt_data_fp16_9, in_wt_data_fp16_8, in_wt_data_fp16_7, in_wt_data_fp16_6, in_wt_data_fp16_5, in_wt_data_fp16_4, in_wt_data_fp16_3, in_wt_data_fp16_2, in_wt_data_fp16_1, in_wt_data_fp16_0 };
  assign in_wt_data_int16 = { in_wt_data_int16_63, in_wt_data_int16_62, in_wt_data_int16_61, in_wt_data_int16_60, in_wt_data_int16_59, in_wt_data_int16_58, in_wt_data_int16_57, in_wt_data_int16_56, in_wt_data_int16_55, in_wt_data_int16_54, in_wt_data_int16_53, in_wt_data_int16_52, in_wt_data_int16_51, in_wt_data_int16_50, in_wt_data_int16_49, in_wt_data_int16_48, in_wt_data_int16_47, in_wt_data_int16_46, in_wt_data_int16_45, in_wt_data_int16_44, in_wt_data_int16_43, in_wt_data_int16_42, in_wt_data_int16_41, in_wt_data_int16_40, in_wt_data_int16_39, in_wt_data_int16_38, in_wt_data_int16_37, in_wt_data_int16_36, in_wt_data_int16_35, in_wt_data_int16_34, in_wt_data_int16_33, in_wt_data_int16_32, in_wt_data_int16_31, in_wt_data_int16_30, in_wt_data_int16_29, in_wt_data_int16_28, in_wt_data_int16_27, in_wt_data_int16_26, in_wt_data_int16_25, in_wt_data_int16_24, in_wt_data_int16_23, in_wt_data_int16_22, in_wt_data_int16_21, in_wt_data_int16_20, in_wt_data_int16_19, in_wt_data_int16_18, in_wt_data_int16_17, in_wt_data_int16_16, in_wt_data_int16_15, in_wt_data_int16_14, in_wt_data_int16_13, in_wt_data_int16_12, in_wt_data_int16_11, in_wt_data_int16_10, in_wt_data_int16_9, in_wt_data_int16_8, in_wt_data_int16_7, in_wt_data_int16_6, in_wt_data_int16_5, in_wt_data_int16_4, in_wt_data_int16_3, in_wt_data_int16_2, in_wt_data_int16_1, in_wt_data_int16_0 };
  assign in_wt_data_int8 = { in_wt_data_int8_63, in_wt_data_int8_62, in_wt_data_int8_61, in_wt_data_int8_60, in_wt_data_int8_59, in_wt_data_int8_58, in_wt_data_int8_57, in_wt_data_int8_56, in_wt_data_int8_55, in_wt_data_int8_54, in_wt_data_int8_53, in_wt_data_int8_52, in_wt_data_int8_51, in_wt_data_int8_50, in_wt_data_int8_49, in_wt_data_int8_48, in_wt_data_int8_47, in_wt_data_int8_46, in_wt_data_int8_45, in_wt_data_int8_44, in_wt_data_int8_43, in_wt_data_int8_42, in_wt_data_int8_41, in_wt_data_int8_40, in_wt_data_int8_39, in_wt_data_int8_38, in_wt_data_int8_37, in_wt_data_int8_36, in_wt_data_int8_35, in_wt_data_int8_34, in_wt_data_int8_33, in_wt_data_int8_32, in_wt_data_int8_31, in_wt_data_int8_30, in_wt_data_int8_29, in_wt_data_int8_28, in_wt_data_int8_27, in_wt_data_int8_26, in_wt_data_int8_25, in_wt_data_int8_24, in_wt_data_int8_23, in_wt_data_int8_22, in_wt_data_int8_21, in_wt_data_int8_20, in_wt_data_int8_19, in_wt_data_int8_18, in_wt_data_int8_17, in_wt_data_int8_16, in_wt_data_int8_15, in_wt_data_int8_14, in_wt_data_int8_13, in_wt_data_int8_12, in_wt_data_int8_11, in_wt_data_int8_10, in_wt_data_int8_9, in_wt_data_int8_8, in_wt_data_int8_7, in_wt_data_int8_6, in_wt_data_int8_5, in_wt_data_int8_4, in_wt_data_int8_3, in_wt_data_int8_2, in_wt_data_int8_1, in_wt_data_int8_0 };
  assign in_wt_data_pack = { in_wt_data127, in_wt_data126, in_wt_data125, in_wt_data124, in_wt_data123, in_wt_data122, in_wt_data121, in_wt_data120, in_wt_data119, in_wt_data118, in_wt_data117, in_wt_data116, in_wt_data115, in_wt_data114, in_wt_data113, in_wt_data112, in_wt_data111, in_wt_data110, in_wt_data109, in_wt_data108, in_wt_data107, in_wt_data106, in_wt_data105, in_wt_data104, in_wt_data103, in_wt_data102, in_wt_data101, in_wt_data100, in_wt_data99, in_wt_data98, in_wt_data97, in_wt_data96, in_wt_data95, in_wt_data94, in_wt_data93, in_wt_data92, in_wt_data91, in_wt_data90, in_wt_data89, in_wt_data88, in_wt_data87, in_wt_data86, in_wt_data85, in_wt_data84, in_wt_data83, in_wt_data82, in_wt_data81, in_wt_data80, in_wt_data79, in_wt_data78, in_wt_data77, in_wt_data76, in_wt_data75, in_wt_data74, in_wt_data73, in_wt_data72, in_wt_data71, in_wt_data70, in_wt_data69, in_wt_data68, in_wt_data67, in_wt_data66, in_wt_data65, in_wt_data64, in_wt_data63, in_wt_data62, in_wt_data61, in_wt_data60, in_wt_data59, in_wt_data58, in_wt_data57, in_wt_data56, in_wt_data55, in_wt_data54, in_wt_data53, in_wt_data52, in_wt_data51, in_wt_data50, in_wt_data49, in_wt_data48, in_wt_data47, in_wt_data46, in_wt_data45, in_wt_data44, in_wt_data43, in_wt_data42, in_wt_data41, in_wt_data40, in_wt_data39, in_wt_data38, in_wt_data37, in_wt_data36, in_wt_data35, in_wt_data34, in_wt_data33, in_wt_data32, in_wt_data31, in_wt_data30, in_wt_data29, in_wt_data28, in_wt_data27, in_wt_data26, in_wt_data25, in_wt_data24, in_wt_data23, in_wt_data22, in_wt_data21, in_wt_data20, in_wt_data19, in_wt_data18, in_wt_data17, in_wt_data16, in_wt_data15, in_wt_data14, in_wt_data13, in_wt_data12, in_wt_data11, in_wt_data10, in_wt_data9, in_wt_data8, in_wt_data7, in_wt_data6, in_wt_data5, in_wt_data4, in_wt_data3, in_wt_data2, in_wt_data1, in_wt_data0 };
  assign in_wt_exp = wt_pre_exp_w;
  assign in_wt_mask_int8 = { in_wt_mask[127], in_wt_mask[63], in_wt_mask[126], in_wt_mask[62], in_wt_mask[125], in_wt_mask[61], in_wt_mask[124], in_wt_mask[60], in_wt_mask[123], in_wt_mask[59], in_wt_mask[122], in_wt_mask[58], in_wt_mask[121], in_wt_mask[57], in_wt_mask[120], in_wt_mask[56], in_wt_mask[119], in_wt_mask[55], in_wt_mask[118], in_wt_mask[54], in_wt_mask[117], in_wt_mask[53], in_wt_mask[116], in_wt_mask[52], in_wt_mask[115], in_wt_mask[51], in_wt_mask[114], in_wt_mask[50], in_wt_mask[113], in_wt_mask[49], in_wt_mask[112], in_wt_mask[48], in_wt_mask[111], in_wt_mask[47], in_wt_mask[110], in_wt_mask[46], in_wt_mask[109], in_wt_mask[45], in_wt_mask[108], in_wt_mask[44], in_wt_mask[107], in_wt_mask[43], in_wt_mask[106], in_wt_mask[42], in_wt_mask[105], in_wt_mask[41], in_wt_mask[104], in_wt_mask[40], in_wt_mask[103], in_wt_mask[39], in_wt_mask[102], in_wt_mask[38], in_wt_mask[101], in_wt_mask[37], in_wt_mask[100], in_wt_mask[36], in_wt_mask[99], in_wt_mask[35], in_wt_mask[98], in_wt_mask[34], in_wt_mask[97], in_wt_mask[33], in_wt_mask[96], in_wt_mask[32], in_wt_mask[95], in_wt_mask[31], in_wt_mask[94], in_wt_mask[30], in_wt_mask[93], in_wt_mask[29], in_wt_mask[92], in_wt_mask[28], in_wt_mask[91], in_wt_mask[27], in_wt_mask[90], in_wt_mask[26], in_wt_mask[89], in_wt_mask[25], in_wt_mask[88], in_wt_mask[24], in_wt_mask[87], in_wt_mask[23], in_wt_mask[86], in_wt_mask[22], in_wt_mask[85], in_wt_mask[21], in_wt_mask[84], in_wt_mask[20], in_wt_mask[83], in_wt_mask[19], in_wt_mask[82], in_wt_mask[18], in_wt_mask[81], in_wt_mask[17], in_wt_mask[80], in_wt_mask[16], in_wt_mask[79], in_wt_mask[15], in_wt_mask[78], in_wt_mask[14], in_wt_mask[77], in_wt_mask[13], in_wt_mask[76], in_wt_mask[12], in_wt_mask[75], in_wt_mask[11], in_wt_mask[74], in_wt_mask[10], in_wt_mask[73], in_wt_mask[9], in_wt_mask[72], in_wt_mask[8], in_wt_mask[71], in_wt_mask[7], in_wt_mask[70], in_wt_mask[6], in_wt_mask[69], in_wt_mask[5], in_wt_mask[68], in_wt_mask[4], in_wt_mask[67], in_wt_mask[3], in_wt_mask[66], in_wt_mask[2], in_wt_mask[65], in_wt_mask[1], in_wt_mask[64], in_wt_mask[0] };
  assign wt0_actv_pvld[103:1] = { wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0], wt0_actv_pvld[0] };
  assign wt0_actv_vld = wt0_actv_pvld[0];
  assign wt1_actv_pvld[103:1] = { wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0], wt1_actv_pvld[0] };
  assign wt1_actv_vld = wt1_actv_pvld[0];
  assign wt2_actv_pvld[103:1] = { wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0], wt2_actv_pvld[0] };
  assign wt2_actv_vld = wt2_actv_pvld[0];
  assign wt3_actv_pvld[103:1] = { wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0], wt3_actv_pvld[0] };
  assign wt3_actv_vld = wt3_actv_pvld[0];
  assign wt4_actv_pvld[103:1] = { wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0], wt4_actv_pvld[0] };
  assign wt4_actv_vld = wt4_actv_pvld[0];
  assign wt5_actv_pvld[103:1] = { wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0], wt5_actv_pvld[0] };
  assign wt5_actv_vld = wt5_actv_pvld[0];
  assign wt6_actv_pvld[103:1] = { wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0], wt6_actv_pvld[0] };
  assign wt6_actv_vld = wt6_actv_pvld[0];
  assign wt7_actv_pvld[103:1] = { wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0], wt7_actv_pvld[0] };
  assign wt7_actv_vld = wt7_actv_pvld[0];
  assign wt_pre_mask_w = { wt_pre_nz_w[126], wt_pre_nz_w[124], wt_pre_nz_w[122], wt_pre_nz_w[120], wt_pre_nz_w[118], wt_pre_nz_w[116], wt_pre_nz_w[114], wt_pre_nz_w[112], wt_pre_nz_w[110], wt_pre_nz_w[108], wt_pre_nz_w[106], wt_pre_nz_w[104], wt_pre_nz_w[102], wt_pre_nz_w[100], wt_pre_nz_w[98], wt_pre_nz_w[96], wt_pre_nz_w[94], wt_pre_nz_w[92], wt_pre_nz_w[90], wt_pre_nz_w[88], wt_pre_nz_w[86], wt_pre_nz_w[84], wt_pre_nz_w[82], wt_pre_nz_w[80], wt_pre_nz_w[78], wt_pre_nz_w[76], wt_pre_nz_w[74], wt_pre_nz_w[72], wt_pre_nz_w[70], wt_pre_nz_w[68], wt_pre_nz_w[66], wt_pre_nz_w[64], wt_pre_nz_w[62], wt_pre_nz_w[60], wt_pre_nz_w[58], wt_pre_nz_w[56], wt_pre_nz_w[54], wt_pre_nz_w[52], wt_pre_nz_w[50], wt_pre_nz_w[48], wt_pre_nz_w[46], wt_pre_nz_w[44], wt_pre_nz_w[42], wt_pre_nz_w[40], wt_pre_nz_w[38], wt_pre_nz_w[36], wt_pre_nz_w[34], wt_pre_nz_w[32], wt_pre_nz_w[30], wt_pre_nz_w[28], wt_pre_nz_w[26], wt_pre_nz_w[24], wt_pre_nz_w[22], wt_pre_nz_w[20], wt_pre_nz_w[18], wt_pre_nz_w[16], wt_pre_nz_w[14], wt_pre_nz_w[12], wt_pre_nz_w[10], wt_pre_nz_w[8], wt_pre_nz_w[6], wt_pre_nz_w[4], wt_pre_nz_w[2], wt_pre_nz_w[0] };
endmodule
