module \$paramod\SDP_C_mgc_in_wire_v1\rscid=7\width=1 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:78" *)
  output d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:79" *)
  input z;
  assign d = z;
endmodule
