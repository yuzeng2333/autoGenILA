module sha_top(clk, rst, wr, addr, data_in, data_out, ack, stb, in_addr_range, xram_addr, xram_data_out, xram_data_in, xram_ack, xram_stb, xram_wr);
  wire [15:0] _000_;
  wire [5:0] _001_;
  wire [15:0] _002_;
  wire [511:0] _003_;
  wire _004_;
  wire [159:0] _005_;
  wire [2:0] _006_;
  wire [5:0] _007_;
  wire [15:0] _008_;
  wire [15:0] _009_;
  wire [15:0] _010_;
  wire [15:0] _011_;
  wire [15:0] _012_;
  wire [31:0] _013_;
  wire [159:0] _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire [2:0] _095_;
  wire [2:0] _096_;
  wire [2:0] _097_;
  wire [2:0] _098_;
  wire [2:0] _099_;
  wire [5:0] _100_;
  wire [5:0] _101_;
  wire [31:0] _102_;
  wire [511:0] _103_;
  wire [7:0] _104_;
  wire [7:0] _105_;
  wire [7:0] _106_;
  wire [15:0] _107_;
  wire [7:0] _108_;
  wire [7:0] _109_;
  wire [7:0] _110_;
  wire [7:0] _111_;
  wire [7:0] _112_;
  wire [7:0] _113_;
  wire [7:0] _114_;
  wire [7:0] _115_;
  wire [7:0] _116_;
  wire [7:0] _117_;
  wire [7:0] _118_;
  wire [7:0] _119_;
  wire [7:0] _120_;
  wire [7:0] _121_;
  wire [7:0] _122_;
  wire [7:0] _123_;
  wire [7:0] _124_;
  wire [7:0] _125_;
  wire [7:0] _126_;
  output ack;
  input [15:0] addr;
  reg [15:0] block_counter;
  wire [15:0] block_counter_next;
  reg [5:0] byte_counter;
  wire [5:0] byte_counter_next;
  wire [5:0] byte_counter_next_rw;
  wire [15:0] bytes_read_next;
  input clk;
  input [7:0] data_in;
  output [7:0] data_out;
  wire [7:0] data_out_len;
  wire [7:0] data_out_rd_addr;
  wire [7:0] data_out_state;
  wire [7:0] data_out_wr_addr;
  output in_addr_range;
  wire read_last_byte_acked;
  wire reading_last_byte;
  reg [15:0] reg_bytes_read;
  input rst;
  wire sel_reg_len;
  wire sel_reg_rd_addr;
  wire sel_reg_start;
  wire sel_reg_state;
  wire sel_reg_wr_addr;
  reg [511:0] sha_core_block;
  wire [511:0] sha_core_block_next;
  wire [511:0] sha_core_block_read_data_next;
  wire [159:0] sha_core_digest;
  wire sha_core_digest_valid;
  wire sha_core_init;
  wire sha_core_next;
  wire sha_core_ready;
  reg sha_core_ready_r;
  wire sha_core_rst_n;
  wire sha_finished;
  wire [15:0] sha_len;
  wire sha_more_blocks;
  wire [15:0] sha_rdaddr;
  reg [159:0] sha_reg_digest;
  wire [67:0] sha_reg_digest_next;
  wire [15:0] sha_reg_len;
  wire [15:0] sha_reg_rd_addr;
  reg [2:0] sha_reg_state;
  wire [15:0] sha_reg_wr_addr;
  wire [2:0] sha_state;
  wire sha_state_idle;
  wire [2:0] sha_state_next;
  wire sha_state_next_idle;
  wire [2:0] sha_state_next_op2;
  wire [1:0] sha_state_next_read_data;
  wire [2:0] sha_state_next_write_data;
  wire sha_state_op1;
  wire sha_state_op2;
  wire sha_state_read_data;
  wire sha_state_write_data;
  wire [15:0] sha_wraddr;
  wire start_op;
  input stb;
  input wr;
  wire wren;
  wire write_last_byte_acked;
  wire writing_last_byte;
  input xram_ack;
  output [15:0] xram_addr;
  input [7:0] xram_data_in;
  output [7:0] xram_data_out;
  output xram_stb;
  output xram_wr;
  assign _007_ = byte_counter + 1'b1;
  assign _008_ = reg_bytes_read + 1'b1;
  assign _009_ = block_counter + 7'b1000000;
  assign _010_ = sha_reg_rd_addr + byte_counter;
  assign _011_ = _010_ + block_counter;
  assign _012_ = sha_reg_wr_addr + byte_counter;
  assign _015_ = byte_counter == 6'b111111;
  assign _016_ = bytes_read_next == sha_reg_len;
  assign _017_ = byte_counter == 6'b111110;
  assign _018_ = byte_counter == 6'b111101;
  assign _019_ = byte_counter == 6'b111100;
  assign _020_ = byte_counter == 6'b111011;
  assign _021_ = byte_counter == 6'b111010;
  assign _022_ = byte_counter == 6'b111001;
  assign _023_ = byte_counter == 6'b111000;
  assign _024_ = byte_counter == 6'b110111;
  assign _025_ = byte_counter == 6'b110110;
  assign _026_ = byte_counter == 6'b110101;
  assign _027_ = byte_counter == 6'b110100;
  assign _028_ = byte_counter == 6'b110011;
  assign _029_ = byte_counter == 6'b110010;
  assign _030_ = byte_counter == 6'b110001;
  assign _031_ = byte_counter == 6'b110000;
  assign _032_ = byte_counter == 6'b101111;
  assign _033_ = byte_counter == 6'b101110;
  assign _034_ = byte_counter == 6'b101101;
  assign _035_ = byte_counter == 6'b101100;
  assign _036_ = byte_counter == 6'b101011;
  assign _037_ = byte_counter == 6'b101010;
  assign _038_ = byte_counter == 6'b101001;
  assign _039_ = byte_counter == 6'b101000;
  assign _040_ = byte_counter == 6'b100111;
  assign _041_ = byte_counter == 6'b100110;
  assign _042_ = byte_counter == 6'b100101;
  assign _043_ = byte_counter == 6'b100100;
  assign _044_ = byte_counter == 6'b100011;
  assign _045_ = byte_counter == 6'b100010;
  assign _046_ = byte_counter == 6'b100001;
  assign _047_ = byte_counter == 6'b100000;
  assign _048_ = byte_counter == 5'b11111;
  assign _049_ = byte_counter == 5'b11110;
  assign _050_ = byte_counter == 5'b11101;
  assign _051_ = byte_counter == 5'b11100;
  assign _052_ = byte_counter == 5'b11011;
  assign _053_ = byte_counter == 5'b11010;
  assign _054_ = byte_counter == 5'b11001;
  assign _055_ = byte_counter == 5'b11000;
  assign _056_ = byte_counter == 5'b10111;
  assign _057_ = byte_counter == 5'b10110;
  assign _058_ = byte_counter == 5'b10101;
  assign _059_ = byte_counter == 5'b10100;
  assign writing_last_byte = byte_counter == 5'b10011;
  assign _060_ = byte_counter == 5'b10010;
  assign _061_ = byte_counter == 5'b10001;
  assign _062_ = byte_counter == 5'b10000;
  assign _063_ = byte_counter == 4'b1111;
  assign _064_ = byte_counter == 4'b1110;
  assign _065_ = byte_counter == 4'b1101;
  assign _066_ = byte_counter == 4'b1100;
  assign _067_ = byte_counter == 4'b1011;
  assign _068_ = byte_counter == 4'b1010;
  assign _069_ = byte_counter == 4'b1001;
  assign _070_ = byte_counter == 4'b1000;
  assign _071_ = byte_counter == 3'b111;
  assign _072_ = byte_counter == 3'b110;
  assign _073_ = byte_counter == 3'b101;
  assign _074_ = byte_counter == 3'b100;
  assign _075_ = byte_counter == 2'b11;
  assign _076_ = byte_counter == 2'b10;
  assign _077_ = byte_counter == 1'b1;
  assign _078_ = ! byte_counter;
  assign _079_ = ! block_counter;
  assign sha_state_idle = ! sha_reg_state;
  assign sha_state_read_data = sha_reg_state == 1'b1;
  assign sha_state_op1 = sha_reg_state == 2'b10;
  assign sha_state_op2 = sha_reg_state == 2'b11;
  assign sha_state_write_data = sha_reg_state == 3'b100;
  assign sel_reg_start = addr == 16'b1111111000000000;
  assign sel_reg_state = addr == 16'b1111111000000001;
  assign sel_reg_rd_addr = addr[15:1] == 15'b111111100000001;
  assign sel_reg_wr_addr = addr[15:1] == 15'b111111100000010;
  assign sel_reg_len = addr[15:1] == 15'b111111100000011;
  assign _080_ = reg_bytes_read >= sha_reg_len;
  assign _081_ = addr >= 16'b1111111000000000;
  assign _082_ = sel_reg_start && data_in[0];
  assign _083_ = _082_ && stb;
  assign start_op = _083_ && wren;
  assign _084_ = sha_state_read_data && xram_ack;
  assign _085_ = sha_state_op2 && sha_more_blocks;
  assign read_last_byte_acked = reading_last_byte && xram_ack;
  assign sha_more_blocks = sha_core_digest_valid && _092_;
  assign sha_finished = sha_core_digest_valid && _080_;
  assign write_last_byte_acked = writing_last_byte && xram_ack;
  assign _086_ = sel_reg_rd_addr && wren;
  assign _087_ = sel_reg_wr_addr && wren;
  assign _088_ = sel_reg_len && wren;
  assign _089_ = sha_state_op1 && sha_core_ready_r;
  assign sha_core_init = _089_ && _079_;
  assign sha_core_next = _089_ && _094_;
  assign in_addr_range = _081_ && _093_;
  assign ack = stb && in_addr_range;
  assign wren = wr && sha_state_idle;
  assign sha_core_rst_n = ! rst;
  assign _090_ = sha_state_idle || sha_state_op1;
  assign _091_ = _090_ || sha_state_op2;
  assign reading_last_byte = _015_ || _016_;
  assign xram_stb = sha_state_read_data || sha_state_write_data;
  assign _092_ = reg_bytes_read < sha_reg_len;
  assign _093_ = addr < 16'b1111111000010000;
  assign _094_ = | block_counter;
  always @(posedge clk)
      sha_reg_state <= _006_;
  always @(posedge clk)
      byte_counter <= _001_;
  always @(posedge clk)
      reg_bytes_read <= _002_;
  always @(posedge clk)
      block_counter <= _000_;
  always @(posedge clk)
      sha_core_ready_r <= _004_;
  always @(posedge clk)
      sha_core_block <= _003_;
  always @(posedge clk)
      sha_reg_digest <= _005_;
  assign _005_ = rst ? 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : { _014_[159:68], sha_reg_digest_next };
  assign _003_ = rst ? 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : sha_core_block_next;
  assign _004_ = rst ? 1'b0 : sha_core_ready;
  assign _000_ = rst ? 16'b0000000000000000 : block_counter_next;
  assign _002_ = rst ? 16'b0000000000000000 : bytes_read_next;
  assign _001_ = rst ? 6'b000000 : byte_counter_next;
  assign _006_ = rst ? 3'b000 : sha_state_next;
  assign _095_ = sha_state_write_data ? sha_state_next_write_data : 3'b000;
  assign _096_ = sha_state_op2 ? sha_state_next_op2 : _095_;
  assign _097_ = sha_state_op1 ? 3'b011 : _096_;
  assign _098_ = sha_state_read_data ? { 1'b0, sha_state_next_read_data } : _097_;
  assign sha_state_next = sha_state_idle ? { 2'b00, start_op } : _098_;
  assign sha_state_next_read_data = read_last_byte_acked ? 2'b10 : 2'b01;
  assign _099_[1:0] = sha_more_blocks ? 2'b01 : 2'b11;
  assign sha_state_next_op2 = sha_finished ? 3'b100 : { 1'b0, _099_[1:0] };
  assign sha_state_next_write_data = write_last_byte_acked ? 3'b000 : 3'b100;
  assign byte_counter_next_rw = xram_ack ? _007_ : byte_counter;
  assign _100_ = sha_state_write_data ? byte_counter_next_rw : byte_counter;
  assign _101_ = sha_state_read_data ? byte_counter_next_rw : _100_;
  assign byte_counter_next = _091_ ? 6'b000000 : _101_;
  assign _102_[15:0] = _084_ ? _008_ : reg_bytes_read;
  assign bytes_read_next = sha_state_idle ? 16'b0000000000000000 : _102_[15:0];
  assign _013_[15:0] = _085_ ? _009_ : block_counter;
  assign block_counter_next = sha_state_idle ? 16'b0000000000000000 : _013_[15:0];
  assign sha_core_block_read_data_next[7:0] = _015_ ? xram_data_in : sha_core_block[7:0];
  assign sha_core_block_read_data_next[15:8] = _017_ ? xram_data_in : sha_core_block[15:8];
  assign sha_core_block_read_data_next[23:16] = _018_ ? xram_data_in : sha_core_block[23:16];
  assign sha_core_block_read_data_next[31:24] = _019_ ? xram_data_in : sha_core_block[31:24];
  assign sha_core_block_read_data_next[39:32] = _020_ ? xram_data_in : sha_core_block[39:32];
  assign sha_core_block_read_data_next[47:40] = _021_ ? xram_data_in : sha_core_block[47:40];
  assign sha_core_block_read_data_next[55:48] = _022_ ? xram_data_in : sha_core_block[55:48];
  assign sha_core_block_read_data_next[63:56] = _023_ ? xram_data_in : sha_core_block[63:56];
  assign sha_core_block_read_data_next[71:64] = _024_ ? xram_data_in : sha_core_block[71:64];
  assign sha_core_block_read_data_next[79:72] = _025_ ? xram_data_in : sha_core_block[79:72];
  assign sha_core_block_read_data_next[87:80] = _026_ ? xram_data_in : sha_core_block[87:80];
  assign sha_core_block_read_data_next[95:88] = _027_ ? xram_data_in : sha_core_block[95:88];
  assign sha_core_block_read_data_next[103:96] = _028_ ? xram_data_in : sha_core_block[103:96];
  assign sha_core_block_read_data_next[111:104] = _029_ ? xram_data_in : sha_core_block[111:104];
  assign sha_core_block_read_data_next[119:112] = _030_ ? xram_data_in : sha_core_block[119:112];
  assign sha_core_block_read_data_next[127:120] = _031_ ? xram_data_in : sha_core_block[127:120];
  assign sha_core_block_read_data_next[135:128] = _032_ ? xram_data_in : sha_core_block[135:128];
  assign sha_core_block_read_data_next[143:136] = _033_ ? xram_data_in : sha_core_block[143:136];
  assign sha_core_block_read_data_next[151:144] = _034_ ? xram_data_in : sha_core_block[151:144];
  assign sha_core_block_read_data_next[159:152] = _035_ ? xram_data_in : sha_core_block[159:152];
  assign sha_core_block_read_data_next[167:160] = _036_ ? xram_data_in : sha_core_block[167:160];
  assign sha_core_block_read_data_next[175:168] = _037_ ? xram_data_in : sha_core_block[175:168];
  assign sha_core_block_read_data_next[183:176] = _038_ ? xram_data_in : sha_core_block[183:176];
  assign sha_core_block_read_data_next[191:184] = _039_ ? xram_data_in : sha_core_block[191:184];
  assign sha_core_block_read_data_next[199:192] = _040_ ? xram_data_in : sha_core_block[199:192];
  assign sha_core_block_read_data_next[207:200] = _041_ ? xram_data_in : sha_core_block[207:200];
  assign sha_core_block_read_data_next[215:208] = _042_ ? xram_data_in : sha_core_block[215:208];
  assign sha_core_block_read_data_next[223:216] = _043_ ? xram_data_in : sha_core_block[223:216];
  assign sha_core_block_read_data_next[231:224] = _044_ ? xram_data_in : sha_core_block[231:224];
  assign sha_core_block_read_data_next[239:232] = _045_ ? xram_data_in : sha_core_block[239:232];
  assign sha_core_block_read_data_next[247:240] = _046_ ? xram_data_in : sha_core_block[247:240];
  assign sha_core_block_read_data_next[255:248] = _047_ ? xram_data_in : sha_core_block[255:248];
  assign sha_core_block_read_data_next[263:256] = _048_ ? xram_data_in : sha_core_block[263:256];
  assign sha_core_block_read_data_next[271:264] = _049_ ? xram_data_in : sha_core_block[271:264];
  assign sha_core_block_read_data_next[279:272] = _050_ ? xram_data_in : sha_core_block[279:272];
  assign sha_core_block_read_data_next[287:280] = _051_ ? xram_data_in : sha_core_block[287:280];
  assign sha_core_block_read_data_next[295:288] = _052_ ? xram_data_in : sha_core_block[295:288];
  assign sha_core_block_read_data_next[303:296] = _053_ ? xram_data_in : sha_core_block[303:296];
  assign sha_core_block_read_data_next[311:304] = _054_ ? xram_data_in : sha_core_block[311:304];
  assign sha_core_block_read_data_next[319:312] = _055_ ? xram_data_in : sha_core_block[319:312];
  assign sha_core_block_read_data_next[327:320] = _056_ ? xram_data_in : sha_core_block[327:320];
  assign sha_core_block_read_data_next[335:328] = _057_ ? xram_data_in : sha_core_block[335:328];
  assign sha_core_block_read_data_next[343:336] = _058_ ? xram_data_in : sha_core_block[343:336];
  assign sha_core_block_read_data_next[351:344] = _059_ ? xram_data_in : sha_core_block[351:344];
  assign sha_core_block_read_data_next[359:352] = writing_last_byte ? xram_data_in : sha_core_block[359:352];
  assign sha_core_block_read_data_next[367:360] = _060_ ? xram_data_in : sha_core_block[367:360];
  assign sha_core_block_read_data_next[375:368] = _061_ ? xram_data_in : sha_core_block[375:368];
  assign sha_core_block_read_data_next[383:376] = _062_ ? xram_data_in : sha_core_block[383:376];
  assign sha_core_block_read_data_next[391:384] = _063_ ? xram_data_in : sha_core_block[391:384];
  assign sha_core_block_read_data_next[399:392] = _064_ ? xram_data_in : sha_core_block[399:392];
  assign sha_core_block_read_data_next[407:400] = _065_ ? xram_data_in : sha_core_block[407:400];
  assign sha_core_block_read_data_next[415:408] = _066_ ? xram_data_in : sha_core_block[415:408];
  assign sha_core_block_read_data_next[423:416] = _067_ ? xram_data_in : sha_core_block[423:416];
  assign sha_core_block_read_data_next[431:424] = _068_ ? xram_data_in : sha_core_block[431:424];
  assign sha_core_block_read_data_next[439:432] = _069_ ? xram_data_in : sha_core_block[439:432];
  assign sha_core_block_read_data_next[447:440] = _070_ ? xram_data_in : sha_core_block[447:440];
  assign sha_core_block_read_data_next[455:448] = _071_ ? xram_data_in : sha_core_block[455:448];
  assign sha_core_block_read_data_next[463:456] = _072_ ? xram_data_in : sha_core_block[463:456];
  assign sha_core_block_read_data_next[471:464] = _073_ ? xram_data_in : sha_core_block[471:464];
  assign sha_core_block_read_data_next[479:472] = _074_ ? xram_data_in : sha_core_block[479:472];
  assign sha_core_block_read_data_next[487:480] = _075_ ? xram_data_in : sha_core_block[487:480];
  assign sha_core_block_read_data_next[495:488] = _076_ ? xram_data_in : sha_core_block[495:488];
  assign sha_core_block_read_data_next[503:496] = _077_ ? xram_data_in : sha_core_block[503:496];
  assign sha_core_block_read_data_next[511:504] = _078_ ? xram_data_in : sha_core_block[511:504];
  assign _103_ = sha_state_read_data ? sha_core_block_read_data_next : sha_core_block;
  assign sha_core_block_next = sha_state_idle ? 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : _103_;
  assign _104_ = sel_reg_len ? data_out_len : 8'b00000000;
  assign _105_ = sel_reg_wr_addr ? data_out_wr_addr : _104_;
  assign _106_ = sel_reg_rd_addr ? data_out_rd_addr : _105_;
  assign data_out = sel_reg_state ? { 5'b00000, sha_reg_state } : _106_;
  assign { _014_[159:68], sha_reg_digest_next } = sha_core_digest_valid ? sha_core_digest : sha_reg_digest;
  assign _107_ = sha_state_write_data ? _012_ : 16'b0000000000000000;
  assign xram_addr = sha_state_read_data ? _011_ : _107_;
  assign _108_ = _078_ ? sha_reg_digest[159:152] : 8'b00000000;
  assign _109_ = _077_ ? sha_reg_digest[151:144] : _108_;
  assign _110_ = _076_ ? sha_reg_digest[143:136] : _109_;
  assign _111_ = _075_ ? sha_reg_digest[135:128] : _110_;
  assign _112_ = _074_ ? sha_reg_digest[127:120] : _111_;
  assign _113_ = _073_ ? sha_reg_digest[119:112] : _112_;
  assign _114_ = _072_ ? sha_reg_digest[111:104] : _113_;
  assign _115_ = _071_ ? sha_reg_digest[103:96] : _114_;
  assign _116_ = _070_ ? sha_reg_digest[95:88] : _115_;
  assign _117_ = _069_ ? sha_reg_digest[87:80] : _116_;
  assign _118_ = _068_ ? sha_reg_digest[79:72] : _117_;
  assign _119_ = _067_ ? sha_reg_digest[71:64] : _118_;
  assign _120_ = _066_ ? sha_reg_digest[63:56] : _119_;
  assign _121_ = _065_ ? sha_reg_digest[55:48] : _120_;
  assign _122_ = _064_ ? sha_reg_digest[47:40] : _121_;
  assign _123_ = _063_ ? sha_reg_digest[39:32] : _122_;
  assign _124_ = _062_ ? sha_reg_digest[31:24] : _123_;
  assign _125_ = _061_ ? sha_reg_digest[23:16] : _124_;
  assign _126_ = _060_ ? sha_reg_digest[15:8] : _125_;
  assign xram_data_out = writing_last_byte ? sha_reg_digest[7:0] : _126_;
  sha1_core sha1_core_i (
    .block(sha_core_block),
    .clk(clk),
    .digest(sha_core_digest),
    .digest_valid(sha_core_digest_valid),
    .init(sha_core_init),
    .next(sha_core_next),
    .ready(sha_core_ready),
    .reset_n(sha_core_rst_n)
  );
  reg2byte sha_reg_len_i (
    .addr(addr[0]),
    .clk(clk),
    .data_in(data_in),
    .data_out(data_out_len),
    .en(sel_reg_len),
    .reg_out(sha_reg_len),
    .rst(rst),
    .wr(_088_)
  );
  reg2byte sha_reg_rd_addr_i (
    .addr(addr[0]),
    .clk(clk),
    .data_in(data_in),
    .data_out(data_out_rd_addr),
    .en(sel_reg_rd_addr),
    .reg_out(sha_reg_rd_addr),
    .rst(rst),
    .wr(_086_)
  );
  reg2byte sha_reg_wr_addr_i (
    .addr(addr[0]),
    .clk(clk),
    .data_in(data_in),
    .data_out(data_out_wr_addr),
    .en(sel_reg_wr_addr),
    .reg_out(sha_reg_wr_addr),
    .rst(rst),
    .wr(_087_)
  );
  assign data_out_state = { 5'b00000, sha_reg_state };
  assign sha_len = sha_reg_len;
  assign sha_rdaddr = sha_reg_rd_addr;
  assign sha_state = sha_reg_state;
  assign sha_state_next_idle = start_op;
  assign sha_wraddr = sha_reg_wr_addr;
  assign xram_wr = sha_state_write_data;
endmodule
