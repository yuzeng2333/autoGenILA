module NV_NVDLA_RT_cmac_b2cacc(nvdla_core_clk, nvdla_core_rstn, mac2accu_src_pvld, mac2accu_src_mask, mac2accu_src_mode, mac2accu_src_data0, mac2accu_src_data1, mac2accu_src_data2, mac2accu_src_data3, mac2accu_src_data4, mac2accu_src_data5, mac2accu_src_data6, mac2accu_src_data7, mac2accu_src_pd, mac2accu_dst_pvld, mac2accu_dst_mask, mac2accu_dst_mode, mac2accu_dst_data0, mac2accu_dst_data1, mac2accu_dst_data2, mac2accu_dst_data3, mac2accu_dst_data4, mac2accu_dst_data5, mac2accu_dst_data6, mac2accu_dst_data7, mac2accu_dst_pd);
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:170" *)
  wire [131:0] _000_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:160" *)
  wire [43:0] _001_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:364" *)
  wire [131:0] _002_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:354" *)
  wire [43:0] _003_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:558" *)
  wire [131:0] _004_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:548" *)
  wire [43:0] _005_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:190" *)
  wire [131:0] _006_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:180" *)
  wire [43:0] _007_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:384" *)
  wire [131:0] _008_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:374" *)
  wire [43:0] _009_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:578" *)
  wire [131:0] _010_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:568" *)
  wire [43:0] _011_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:210" *)
  wire [131:0] _012_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:200" *)
  wire [43:0] _013_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:404" *)
  wire [131:0] _014_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:394" *)
  wire [43:0] _015_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:598" *)
  wire [131:0] _016_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:588" *)
  wire [43:0] _017_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:230" *)
  wire [131:0] _018_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:220" *)
  wire [43:0] _019_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:424" *)
  wire [131:0] _020_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:414" *)
  wire [43:0] _021_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:618" *)
  wire [131:0] _022_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:608" *)
  wire [43:0] _023_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:250" *)
  wire [131:0] _024_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:240" *)
  wire [43:0] _025_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:444" *)
  wire [131:0] _026_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:434" *)
  wire [43:0] _027_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:638" *)
  wire [131:0] _028_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:628" *)
  wire [43:0] _029_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:270" *)
  wire [131:0] _030_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:260" *)
  wire [43:0] _031_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:464" *)
  wire [131:0] _032_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:454" *)
  wire [43:0] _033_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:658" *)
  wire [131:0] _034_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:648" *)
  wire [43:0] _035_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:290" *)
  wire [131:0] _036_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:280" *)
  wire [43:0] _037_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:484" *)
  wire [131:0] _038_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:474" *)
  wire [43:0] _039_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:678" *)
  wire [131:0] _040_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:668" *)
  wire [43:0] _041_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:310" *)
  wire [131:0] _042_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:300" *)
  wire [43:0] _043_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:504" *)
  wire [131:0] _044_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:494" *)
  wire [43:0] _045_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:698" *)
  wire [131:0] _046_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:688" *)
  wire [43:0] _047_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:143" *)
  wire [7:0] _048_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:337" *)
  wire [7:0] _049_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:531" *)
  wire [7:0] _050_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:133" *)
  wire [8:0] _051_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:327" *)
  wire [8:0] _052_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:521" *)
  wire [8:0] _053_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:171" *)
  wire _054_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:191" *)
  wire _055_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:211" *)
  wire _056_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:231" *)
  wire _057_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:251" *)
  wire _058_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:271" *)
  wire _059_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:291" *)
  wire _060_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:311" *)
  wire _061_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:365" *)
  wire _062_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:385" *)
  wire _063_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:405" *)
  wire _064_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:425" *)
  wire _065_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:445" *)
  wire _066_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:465" *)
  wire _067_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:485" *)
  wire _068_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:505" *)
  wire _069_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:559" *)
  wire _070_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:579" *)
  wire _071_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:599" *)
  wire _072_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:619" *)
  wire _073_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:639" *)
  wire _074_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:659" *)
  wire _075_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:679" *)
  wire _076_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:699" *)
  wire _077_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:66" *)
  wire [175:0] mac2accu_data0_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:78" *)
  reg [175:0] mac2accu_data0_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:79" *)
  reg [175:0] mac2accu_data0_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:80" *)
  reg [175:0] mac2accu_data0_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:67" *)
  wire [175:0] mac2accu_data1_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:81" *)
  reg [175:0] mac2accu_data1_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:82" *)
  reg [175:0] mac2accu_data1_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:83" *)
  reg [175:0] mac2accu_data1_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:68" *)
  wire [175:0] mac2accu_data2_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:84" *)
  reg [175:0] mac2accu_data2_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:85" *)
  reg [175:0] mac2accu_data2_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:86" *)
  reg [175:0] mac2accu_data2_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:69" *)
  wire [175:0] mac2accu_data3_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:87" *)
  reg [175:0] mac2accu_data3_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:88" *)
  reg [175:0] mac2accu_data3_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:89" *)
  reg [175:0] mac2accu_data3_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:70" *)
  wire [175:0] mac2accu_data4_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:90" *)
  reg [175:0] mac2accu_data4_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:91" *)
  reg [175:0] mac2accu_data4_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:92" *)
  reg [175:0] mac2accu_data4_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:71" *)
  wire [175:0] mac2accu_data5_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:93" *)
  reg [175:0] mac2accu_data5_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:94" *)
  reg [175:0] mac2accu_data5_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:95" *)
  reg [175:0] mac2accu_data5_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:72" *)
  wire [175:0] mac2accu_data6_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:96" *)
  reg [175:0] mac2accu_data6_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:97" *)
  reg [175:0] mac2accu_data6_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:98" *)
  reg [175:0] mac2accu_data6_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:73" *)
  wire [175:0] mac2accu_data7_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:99" *)
  reg [175:0] mac2accu_data7_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:100" *)
  reg [175:0] mac2accu_data7_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:101" *)
  reg [175:0] mac2accu_data7_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:57" *)
  output [175:0] mac2accu_dst_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:58" *)
  output [175:0] mac2accu_dst_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:59" *)
  output [175:0] mac2accu_dst_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:60" *)
  output [175:0] mac2accu_dst_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:61" *)
  output [175:0] mac2accu_dst_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:62" *)
  output [175:0] mac2accu_dst_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:63" *)
  output [175:0] mac2accu_dst_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:64" *)
  output [175:0] mac2accu_dst_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:55" *)
  output [7:0] mac2accu_dst_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:56" *)
  output [7:0] mac2accu_dst_mode;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:65" *)
  output [8:0] mac2accu_dst_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:54" *)
  output mac2accu_dst_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:74" *)
  wire [7:0] mac2accu_mask_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:102" *)
  reg [7:0] mac2accu_mask_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:103" *)
  reg [7:0] mac2accu_mask_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:104" *)
  reg [7:0] mac2accu_mask_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:75" *)
  wire [7:0] mac2accu_mode_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:105" *)
  reg [7:0] mac2accu_mode_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:106" *)
  reg [7:0] mac2accu_mode_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:107" *)
  reg [7:0] mac2accu_mode_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:76" *)
  wire [8:0] mac2accu_pd_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:108" *)
  reg [8:0] mac2accu_pd_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:109" *)
  reg [8:0] mac2accu_pd_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:110" *)
  reg [8:0] mac2accu_pd_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:77" *)
  wire mac2accu_pvld_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:111" *)
  reg mac2accu_pvld_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:112" *)
  reg mac2accu_pvld_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:113" *)
  reg mac2accu_pvld_d3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:45" *)
  input [175:0] mac2accu_src_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:46" *)
  input [175:0] mac2accu_src_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:47" *)
  input [175:0] mac2accu_src_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:48" *)
  input [175:0] mac2accu_src_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:49" *)
  input [175:0] mac2accu_src_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:50" *)
  input [175:0] mac2accu_src_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:51" *)
  input [175:0] mac2accu_src_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:52" *)
  input [175:0] mac2accu_src_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:43" *)
  input [7:0] mac2accu_src_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:44" *)
  input [7:0] mac2accu_src_mode;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:53" *)
  input [8:0] mac2accu_src_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:42" *)
  input mac2accu_src_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:40" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:41" *)
  input nvdla_core_rstn;
  assign _054_ = mac2accu_src_mask[0] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:171" *) mac2accu_src_mode[0];
  assign _055_ = mac2accu_src_mask[1] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:191" *) mac2accu_src_mode[1];
  assign _056_ = mac2accu_src_mask[2] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:211" *) mac2accu_src_mode[2];
  assign _057_ = mac2accu_src_mask[3] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:231" *) mac2accu_src_mode[3];
  assign _058_ = mac2accu_src_mask[4] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:251" *) mac2accu_src_mode[4];
  assign _059_ = mac2accu_src_mask[5] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:271" *) mac2accu_src_mode[5];
  assign _060_ = mac2accu_src_mask[6] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:291" *) mac2accu_src_mode[6];
  assign _061_ = mac2accu_src_mask[7] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:311" *) mac2accu_src_mode[7];
  assign _062_ = mac2accu_mask_d1[0] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:365" *) mac2accu_mode_d1[0];
  assign _063_ = mac2accu_mask_d1[1] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:385" *) mac2accu_mode_d1[1];
  assign _064_ = mac2accu_mask_d1[2] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:405" *) mac2accu_mode_d1[2];
  assign _065_ = mac2accu_mask_d1[3] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:425" *) mac2accu_mode_d1[3];
  assign _066_ = mac2accu_mask_d1[4] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:445" *) mac2accu_mode_d1[4];
  assign _067_ = mac2accu_mask_d1[5] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:465" *) mac2accu_mode_d1[5];
  assign _068_ = mac2accu_mask_d1[6] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:485" *) mac2accu_mode_d1[6];
  assign _069_ = mac2accu_mask_d1[7] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:505" *) mac2accu_mode_d1[7];
  assign _070_ = mac2accu_mask_d2[0] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:559" *) mac2accu_mode_d2[0];
  assign _071_ = mac2accu_mask_d2[1] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:579" *) mac2accu_mode_d2[1];
  assign _072_ = mac2accu_mask_d2[2] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:599" *) mac2accu_mode_d2[2];
  assign _073_ = mac2accu_mask_d2[3] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:619" *) mac2accu_mode_d2[3];
  assign _074_ = mac2accu_mask_d2[4] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:639" *) mac2accu_mode_d2[4];
  assign _075_ = mac2accu_mask_d2[5] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:659" *) mac2accu_mode_d2[5];
  assign _076_ = mac2accu_mask_d2[6] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:679" *) mac2accu_mode_d2[6];
  assign _077_ = mac2accu_mask_d2[7] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:699" *) mac2accu_mode_d2[7];
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d3[175:44] <= _046_;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d3[43:0] <= _047_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d3[175:44] <= _040_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d3[43:0] <= _041_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d3[175:44] <= _034_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d3[43:0] <= _035_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d3[175:44] <= _028_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d3[43:0] <= _029_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d3[175:44] <= _022_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d3[43:0] <= _023_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d3[175:44] <= _016_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d3[43:0] <= _017_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d3[175:44] <= _010_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d3[43:0] <= _011_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d3[175:44] <= _004_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d3[43:0] <= _005_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_mask_d3 <= 8'b00000000;
    else
      mac2accu_mask_d3 <= mac2accu_mask_d2;
  always @(posedge nvdla_core_clk)
      mac2accu_mode_d3 <= _050_;
  always @(posedge nvdla_core_clk)
      mac2accu_pd_d3 <= _053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_pvld_d3 <= 1'b0;
    else
      mac2accu_pvld_d3 <= mac2accu_pvld_d2;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d2[175:44] <= _044_;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d2[43:0] <= _045_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d2[175:44] <= _038_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d2[43:0] <= _039_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d2[175:44] <= _032_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d2[43:0] <= _033_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d2[175:44] <= _026_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d2[43:0] <= _027_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d2[175:44] <= _020_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d2[43:0] <= _021_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d2[175:44] <= _014_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d2[43:0] <= _015_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d2[175:44] <= _008_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d2[43:0] <= _009_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d2[175:44] <= _002_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d2[43:0] <= _003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_mask_d2 <= 8'b00000000;
    else
      mac2accu_mask_d2 <= mac2accu_mask_d1;
  always @(posedge nvdla_core_clk)
      mac2accu_mode_d2 <= _049_;
  always @(posedge nvdla_core_clk)
      mac2accu_pd_d2 <= _052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_pvld_d2 <= 1'b0;
    else
      mac2accu_pvld_d2 <= mac2accu_pvld_d1;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d1[175:44] <= _042_;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d1[43:0] <= _043_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d1[175:44] <= _036_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d1[43:0] <= _037_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d1[175:44] <= _030_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d1[43:0] <= _031_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d1[175:44] <= _024_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d1[43:0] <= _025_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d1[175:44] <= _018_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d1[43:0] <= _019_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d1[175:44] <= _012_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d1[43:0] <= _013_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d1[175:44] <= _006_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d1[43:0] <= _007_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d1[175:44] <= _000_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d1[43:0] <= _001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_mask_d1 <= 8'b00000000;
    else
      mac2accu_mask_d1 <= mac2accu_src_mask;
  always @(posedge nvdla_core_clk)
      mac2accu_mode_d1 <= _048_;
  always @(posedge nvdla_core_clk)
      mac2accu_pd_d1 <= _051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_pvld_d1 <= 1'b0;
    else
      mac2accu_pvld_d1 <= mac2accu_src_pvld;
  assign _046_ = _077_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:699" *) mac2accu_data7_d2[175:44] : mac2accu_data7_d3[175:44];
  assign _047_ = mac2accu_mask_d2[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:689" *) mac2accu_data7_d2[43:0] : mac2accu_data7_d3[43:0];
  assign _040_ = _076_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:679" *) mac2accu_data6_d2[175:44] : mac2accu_data6_d3[175:44];
  assign _041_ = mac2accu_mask_d2[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:669" *) mac2accu_data6_d2[43:0] : mac2accu_data6_d3[43:0];
  assign _034_ = _075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:659" *) mac2accu_data5_d2[175:44] : mac2accu_data5_d3[175:44];
  assign _035_ = mac2accu_mask_d2[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:649" *) mac2accu_data5_d2[43:0] : mac2accu_data5_d3[43:0];
  assign _028_ = _074_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:639" *) mac2accu_data4_d2[175:44] : mac2accu_data4_d3[175:44];
  assign _029_ = mac2accu_mask_d2[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:629" *) mac2accu_data4_d2[43:0] : mac2accu_data4_d3[43:0];
  assign _022_ = _073_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:619" *) mac2accu_data3_d2[175:44] : mac2accu_data3_d3[175:44];
  assign _023_ = mac2accu_mask_d2[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:609" *) mac2accu_data3_d2[43:0] : mac2accu_data3_d3[43:0];
  assign _016_ = _072_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:599" *) mac2accu_data2_d2[175:44] : mac2accu_data2_d3[175:44];
  assign _017_ = mac2accu_mask_d2[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:589" *) mac2accu_data2_d2[43:0] : mac2accu_data2_d3[43:0];
  assign _010_ = _071_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:579" *) mac2accu_data1_d2[175:44] : mac2accu_data1_d3[175:44];
  assign _011_ = mac2accu_mask_d2[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:569" *) mac2accu_data1_d2[43:0] : mac2accu_data1_d3[43:0];
  assign _004_ = _070_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:559" *) mac2accu_data0_d2[175:44] : mac2accu_data0_d3[175:44];
  assign _005_ = mac2accu_mask_d2[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:549" *) mac2accu_data0_d2[43:0] : mac2accu_data0_d3[43:0];
  assign _050_ = mac2accu_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:532" *) mac2accu_mode_d2 : mac2accu_mode_d3;
  assign _053_ = mac2accu_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:522" *) mac2accu_pd_d2 : mac2accu_pd_d3;
  assign _044_ = _069_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:505" *) mac2accu_data7_d1[175:44] : mac2accu_data7_d2[175:44];
  assign _045_ = mac2accu_mask_d1[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:495" *) mac2accu_data7_d1[43:0] : mac2accu_data7_d2[43:0];
  assign _038_ = _068_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:485" *) mac2accu_data6_d1[175:44] : mac2accu_data6_d2[175:44];
  assign _039_ = mac2accu_mask_d1[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:475" *) mac2accu_data6_d1[43:0] : mac2accu_data6_d2[43:0];
  assign _032_ = _067_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:465" *) mac2accu_data5_d1[175:44] : mac2accu_data5_d2[175:44];
  assign _033_ = mac2accu_mask_d1[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:455" *) mac2accu_data5_d1[43:0] : mac2accu_data5_d2[43:0];
  assign _026_ = _066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:445" *) mac2accu_data4_d1[175:44] : mac2accu_data4_d2[175:44];
  assign _027_ = mac2accu_mask_d1[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:435" *) mac2accu_data4_d1[43:0] : mac2accu_data4_d2[43:0];
  assign _020_ = _065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:425" *) mac2accu_data3_d1[175:44] : mac2accu_data3_d2[175:44];
  assign _021_ = mac2accu_mask_d1[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:415" *) mac2accu_data3_d1[43:0] : mac2accu_data3_d2[43:0];
  assign _014_ = _064_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:405" *) mac2accu_data2_d1[175:44] : mac2accu_data2_d2[175:44];
  assign _015_ = mac2accu_mask_d1[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:395" *) mac2accu_data2_d1[43:0] : mac2accu_data2_d2[43:0];
  assign _008_ = _063_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:385" *) mac2accu_data1_d1[175:44] : mac2accu_data1_d2[175:44];
  assign _009_ = mac2accu_mask_d1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:375" *) mac2accu_data1_d1[43:0] : mac2accu_data1_d2[43:0];
  assign _002_ = _062_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:365" *) mac2accu_data0_d1[175:44] : mac2accu_data0_d2[175:44];
  assign _003_ = mac2accu_mask_d1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:355" *) mac2accu_data0_d1[43:0] : mac2accu_data0_d2[43:0];
  assign _049_ = mac2accu_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:338" *) mac2accu_mode_d1 : mac2accu_mode_d2;
  assign _052_ = mac2accu_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:328" *) mac2accu_pd_d1 : mac2accu_pd_d2;
  assign _042_ = _061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:311" *) mac2accu_src_data7[175:44] : mac2accu_data7_d1[175:44];
  assign _043_ = mac2accu_src_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:301" *) mac2accu_src_data7[43:0] : mac2accu_data7_d1[43:0];
  assign _036_ = _060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:291" *) mac2accu_src_data6[175:44] : mac2accu_data6_d1[175:44];
  assign _037_ = mac2accu_src_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:281" *) mac2accu_src_data6[43:0] : mac2accu_data6_d1[43:0];
  assign _030_ = _059_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:271" *) mac2accu_src_data5[175:44] : mac2accu_data5_d1[175:44];
  assign _031_ = mac2accu_src_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:261" *) mac2accu_src_data5[43:0] : mac2accu_data5_d1[43:0];
  assign _024_ = _058_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:251" *) mac2accu_src_data4[175:44] : mac2accu_data4_d1[175:44];
  assign _025_ = mac2accu_src_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:241" *) mac2accu_src_data4[43:0] : mac2accu_data4_d1[43:0];
  assign _018_ = _057_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:231" *) mac2accu_src_data3[175:44] : mac2accu_data3_d1[175:44];
  assign _019_ = mac2accu_src_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:221" *) mac2accu_src_data3[43:0] : mac2accu_data3_d1[43:0];
  assign _012_ = _056_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:211" *) mac2accu_src_data2[175:44] : mac2accu_data2_d1[175:44];
  assign _013_ = mac2accu_src_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:201" *) mac2accu_src_data2[43:0] : mac2accu_data2_d1[43:0];
  assign _006_ = _055_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:191" *) mac2accu_src_data1[175:44] : mac2accu_data1_d1[175:44];
  assign _007_ = mac2accu_src_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:181" *) mac2accu_src_data1[43:0] : mac2accu_data1_d1[43:0];
  assign _000_ = _054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:171" *) mac2accu_src_data0[175:44] : mac2accu_data0_d1[175:44];
  assign _001_ = mac2accu_src_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:161" *) mac2accu_src_data0[43:0] : mac2accu_data0_d1[43:0];
  assign _048_ = mac2accu_src_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:144" *) mac2accu_src_mode : mac2accu_mode_d1;
  assign _051_ = mac2accu_src_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_b2cacc.v:134" *) mac2accu_src_pd : mac2accu_pd_d1;
  assign mac2accu_data0_d0 = mac2accu_src_data0;
  assign mac2accu_data1_d0 = mac2accu_src_data1;
  assign mac2accu_data2_d0 = mac2accu_src_data2;
  assign mac2accu_data3_d0 = mac2accu_src_data3;
  assign mac2accu_data4_d0 = mac2accu_src_data4;
  assign mac2accu_data5_d0 = mac2accu_src_data5;
  assign mac2accu_data6_d0 = mac2accu_src_data6;
  assign mac2accu_data7_d0 = mac2accu_src_data7;
  assign mac2accu_dst_data0 = mac2accu_data0_d3;
  assign mac2accu_dst_data1 = mac2accu_data1_d3;
  assign mac2accu_dst_data2 = mac2accu_data2_d3;
  assign mac2accu_dst_data3 = mac2accu_data3_d3;
  assign mac2accu_dst_data4 = mac2accu_data4_d3;
  assign mac2accu_dst_data5 = mac2accu_data5_d3;
  assign mac2accu_dst_data6 = mac2accu_data6_d3;
  assign mac2accu_dst_data7 = mac2accu_data7_d3;
  assign mac2accu_dst_mask = mac2accu_mask_d3;
  assign mac2accu_dst_mode = mac2accu_mode_d3;
  assign mac2accu_dst_pd = mac2accu_pd_d3;
  assign mac2accu_dst_pvld = mac2accu_pvld_d3;
  assign mac2accu_mask_d0 = mac2accu_src_mask;
  assign mac2accu_mode_d0 = mac2accu_src_mode;
  assign mac2accu_pd_d0 = mac2accu_src_pd;
  assign mac2accu_pvld_d0 = mac2accu_src_pvld;
endmodule
