module memory_to_color(color_depth_i, mem_i, mem_lsb_i, color_o, sel_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire [3:0] _13_;
  wire [31:0] _14_;
  wire [31:0] _15_;
  wire [31:0] _16_;
  wire [31:0] _17_;
  wire [31:0] _18_;
  input [1:0] color_depth_i;
  output [31:0] color_o;
  input [31:0] mem_i;
  input [1:0] mem_lsb_i;
  output [3:0] sel_o;
  assign _00_ = ! color_depth_i;
  assign _01_ = color_depth_i == 1'b1;
  assign _02_ = ! mem_lsb_i;
  assign _03_ = mem_lsb_i == 1'b1;
  assign _04_ = mem_lsb_i == 2'b10;
  assign _05_ = mem_lsb_i == 2'b11;
  assign _06_ = ~ mem_lsb_i[0];
  assign _07_ = _00_ && _02_;
  assign _08_ = _00_ && _03_;
  assign _09_ = _00_ && _04_;
  assign _10_ = _00_ && _05_;
  assign _11_ = _01_ && _06_;
  assign _12_ = _01_ && mem_lsb_i[0];
  assign _13_ = _01_ ? 4'b0011 : 4'b1111;
  assign sel_o = _00_ ? 4'b0001 : _13_;
  assign _14_ = _12_ ? { 16'b0000000000000000, mem_i[15:0] } : mem_i;
  assign _15_ = _11_ ? { 16'b0000000000000000, mem_i[31:16] } : _14_;
  assign _16_ = _10_ ? { 24'b000000000000000000000000, mem_i[7:0] } : _15_;
  assign _17_ = _09_ ? { 24'b000000000000000000000000, mem_i[15:8] } : _16_;
  assign _18_ = _08_ ? { 24'b000000000000000000000000, mem_i[23:16] } : _17_;
  assign color_o = _07_ ? { 24'b000000000000000000000000, mem_i[31:24] } : _18_;
endmodule
