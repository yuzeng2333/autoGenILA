module FP32_SUB_chn_b_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_sub.v:352" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_sub.v:353" *)
  output outsig;
  assign outsig = in_0;
endmodule
