module HLS_fp17_add_core_chn_a_rsci_chn_a_wait_ctrl(nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, core_wen, chn_a_rsci_iswt0, chn_a_rsci_ld_core_psct, core_wten, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_ld_core_sct, chn_a_rsci_vd);
  (* src = "./vmod/vlibs/HLS_fp17_add.v:606" *)
  wire _00_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:601" *)
  wire _01_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:611" *)
  wire _02_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:611" *)
  wire _03_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:593" *)
  output chn_a_rsci_bdwt;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:592" *)
  output chn_a_rsci_biwt;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:599" *)
  reg chn_a_rsci_icwt;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:589" *)
  input chn_a_rsci_iswt0;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:590" *)
  input chn_a_rsci_ld_core_psct;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:594" *)
  output chn_a_rsci_ld_core_sct;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:597" *)
  wire chn_a_rsci_ogwt;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:587" *)
  input chn_a_rsci_oswt;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:598" *)
  wire chn_a_rsci_pdswt0;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:595" *)
  input chn_a_rsci_vd;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:588" *)
  input core_wen;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:591" *)
  input core_wten;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:585" *)
  input nvdla_core_clk;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:586" *)
  input nvdla_core_rstn;
  assign chn_a_rsci_pdswt0 = _01_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:601" *) chn_a_rsci_iswt0;
  assign chn_a_rsci_biwt = chn_a_rsci_ogwt & (* src = "./vmod/vlibs/HLS_fp17_add.v:602" *) chn_a_rsci_vd;
  assign chn_a_rsci_bdwt = chn_a_rsci_oswt & (* src = "./vmod/vlibs/HLS_fp17_add.v:604" *) core_wen;
  assign chn_a_rsci_ld_core_sct = chn_a_rsci_ld_core_psct & (* src = "./vmod/vlibs/HLS_fp17_add.v:605" *) chn_a_rsci_ogwt;
  assign _01_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:601" *) core_wten;
  assign _02_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:611" *) chn_a_rsci_ogwt;
  assign _00_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:611" *) _03_;
  assign chn_a_rsci_ogwt = chn_a_rsci_pdswt0 | (* src = "./vmod/vlibs/HLS_fp17_add.v:603" *) chn_a_rsci_icwt;
  assign _03_ = _02_ | (* src = "./vmod/vlibs/HLS_fp17_add.v:611" *) chn_a_rsci_biwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_a_rsci_icwt <= 1'b0;
    else
      chn_a_rsci_icwt <= _00_;
endmodule
