module bar__DOT__i1(
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
in,
out,
__COUNTER_start__n0
);
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg      [7:0] in;
output reg      [7:0] out;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire      [7:0] bv_8_0_n406;
wire      [7:0] bv_8_100_n298;
wire      [7:0] bv_8_101_n190;
wire      [7:0] bv_8_102_n128;
wire      [7:0] bv_8_103_n369;
wire      [7:0] bv_8_104_n27;
wire      [7:0] bv_8_105_n82;
wire      [7:0] bv_8_106_n363;
wire      [7:0] bv_8_107_n361;
wire      [7:0] bv_8_108_n197;
wire      [7:0] bv_8_109_n209;
wire      [7:0] bv_8_10_n247;
wire      [7:0] bv_8_110_n355;
wire      [7:0] bv_8_111_n353;
wire      [7:0] bv_8_112_n137;
wire      [7:0] bv_8_113_n349;
wire      [7:0] bv_8_114_n346;
wire      [7:0] bv_8_115_n292;
wire      [7:0] bv_8_116_n154;
wire      [7:0] bv_8_117_n342;
wire      [7:0] bv_8_118_n339;
wire      [7:0] bv_8_119_n337;
wire      [7:0] bv_8_11_n258;
wire      [7:0] bv_8_120_n177;
wire      [7:0] bv_8_121_n218;
wire      [7:0] bv_8_122_n187;
wire      [7:0] bv_8_123_n331;
wire      [7:0] bv_8_124_n328;
wire      [7:0] bv_8_125_n326;
wire      [7:0] bv_8_126_n302;
wire      [7:0] bv_8_127_n323;
wire      [7:0] bv_8_128_n321;
wire      [7:0] bv_8_129_n287;
wire      [7:0] bv_8_12_n320;
wire      [7:0] bv_8_130_n316;
wire      [7:0] bv_8_131_n314;
wire      [7:0] bv_8_132_n311;
wire      [7:0] bv_8_133_n309;
wire      [7:0] bv_8_134_n103;
wire      [7:0] bv_8_135_n66;
wire      [7:0] bv_8_136_n273;
wire      [7:0] bv_8_137_n42;
wire      [7:0] bv_8_138_n140;
wire      [7:0] bv_8_139_n142;
wire      [7:0] bv_8_13_n39;
wire      [7:0] bv_8_140_n48;
wire      [7:0] bv_8_141_n206;
wire      [7:0] bv_8_142_n76;
wire      [7:0] bv_8_143_n290;
wire      [7:0] bv_8_144_n276;
wire      [7:0] bv_8_145_n225;
wire      [7:0] bv_8_146_n283;
wire      [7:0] bv_8_147_n281;
wire      [7:0] bv_8_148_n74;
wire      [7:0] bv_8_149_n222;
wire      [7:0] bv_8_14_n117;
wire      [7:0] bv_8_150_n274;
wire      [7:0] bv_8_151_n271;
wire      [7:0] bv_8_152_n88;
wire      [7:0] bv_8_153_n21;
wire      [7:0] bv_8_154_n266;
wire      [7:0] bv_8_155_n71;
wire      [7:0] bv_8_156_n262;
wire      [7:0] bv_8_157_n259;
wire      [7:0] bv_8_158_n94;
wire      [7:0] bv_8_159_n255;
wire      [7:0] bv_8_15_n15;
wire      [7:0] bv_8_160_n253;
wire      [7:0] bv_8_161_n45;
wire      [7:0] bv_8_162_n248;
wire      [7:0] bv_8_163_n245;
wire      [7:0] bv_8_164_n242;
wire      [7:0] bv_8_165_n239;
wire      [7:0] bv_8_166_n166;
wire      [7:0] bv_8_167_n234;
wire      [7:0] bv_8_168_n232;
wire      [7:0] bv_8_169_n200;
wire      [7:0] bv_8_16_n330;
wire      [7:0] bv_8_170_n229;
wire      [7:0] bv_8_171_n226;
wire      [7:0] bv_8_172_n223;
wire      [7:0] bv_8_173_n220;
wire      [7:0] bv_8_174_n185;
wire      [7:0] bv_8_175_n216;
wire      [7:0] bv_8_176_n12;
wire      [7:0] bv_8_177_n213;
wire      [7:0] bv_8_178_n210;
wire      [7:0] bv_8_179_n207;
wire      [7:0] bv_8_17_n85;
wire      [7:0] bv_8_180_n163;
wire      [7:0] bv_8_181_n131;
wire      [7:0] bv_8_182_n201;
wire      [7:0] bv_8_183_n198;
wire      [7:0] bv_8_184_n195;
wire      [7:0] bv_8_185_n106;
wire      [7:0] bv_8_186_n180;
wire      [7:0] bv_8_187_n6;
wire      [7:0] bv_8_188_n188;
wire      [7:0] bv_8_189_n145;
wire      [7:0] bv_8_18_n442;
wire      [7:0] bv_8_190_n183;
wire      [7:0] bv_8_191_n36;
wire      [7:0] bv_8_192_n178;
wire      [7:0] bv_8_193_n100;
wire      [7:0] bv_8_194_n173;
wire      [7:0] bv_8_195_n170;
wire      [7:0] bv_8_196_n167;
wire      [7:0] bv_8_197_n164;
wire      [7:0] bv_8_198_n161;
wire      [7:0] bv_8_199_n159;
wire      [7:0] bv_8_19_n318;
wire      [7:0] bv_8_1_n503;
wire      [7:0] bv_8_200_n157;
wire      [7:0] bv_8_201_n155;
wire      [7:0] bv_8_202_n152;
wire      [7:0] bv_8_203_n149;
wire      [7:0] bv_8_204_n146;
wire      [7:0] bv_8_205_n143;
wire      [7:0] bv_8_206_n60;
wire      [7:0] bv_8_207_n138;
wire      [7:0] bv_8_208_n135;
wire      [7:0] bv_8_209_n132;
wire      [7:0] bv_8_20_n265;
wire      [7:0] bv_8_210_n129;
wire      [7:0] bv_8_211_n126;
wire      [7:0] bv_8_212_n123;
wire      [7:0] bv_8_213_n120;
wire      [7:0] bv_8_214_n118;
wire      [7:0] bv_8_215_n115;
wire      [7:0] bv_8_216_n112;
wire      [7:0] bv_8_217_n79;
wire      [7:0] bv_8_218_n107;
wire      [7:0] bv_8_219_n104;
wire      [7:0] bv_8_21_n462;
wire      [7:0] bv_8_220_n101;
wire      [7:0] bv_8_221_n98;
wire      [7:0] bv_8_222_n95;
wire      [7:0] bv_8_223_n51;
wire      [7:0] bv_8_224_n91;
wire      [7:0] bv_8_225_n89;
wire      [7:0] bv_8_226_n86;
wire      [7:0] bv_8_227_n83;
wire      [7:0] bv_8_228_n80;
wire      [7:0] bv_8_229_n77;
wire      [7:0] bv_8_22_n3;
wire      [7:0] bv_8_230_n33;
wire      [7:0] bv_8_231_n72;
wire      [7:0] bv_8_232_n69;
wire      [7:0] bv_8_233_n63;
wire      [7:0] bv_8_234_n64;
wire      [7:0] bv_8_235_n61;
wire      [7:0] bv_8_236_n58;
wire      [7:0] bv_8_237_n55;
wire      [7:0] bv_8_238_n52;
wire      [7:0] bv_8_239_n49;
wire      [7:0] bv_8_23_n306;
wire      [7:0] bv_8_240_n46;
wire      [7:0] bv_8_241_n43;
wire      [7:0] bv_8_242_n40;
wire      [7:0] bv_8_243_n37;
wire      [7:0] bv_8_244_n34;
wire      [7:0] bv_8_245_n31;
wire      [7:0] bv_8_246_n28;
wire      [7:0] bv_8_247_n25;
wire      [7:0] bv_8_248_n22;
wire      [7:0] bv_8_249_n19;
wire      [7:0] bv_8_24_n452;
wire      [7:0] bv_8_250_n16;
wire      [7:0] bv_8_251_n13;
wire      [7:0] bv_8_252_n10;
wire      [7:0] bv_8_253_n7;
wire      [7:0] bv_8_254_n4;
wire      [7:0] bv_8_255_n1;
wire      [7:0] bv_8_25_n294;
wire      [7:0] bv_8_26_n427;
wire      [7:0] bv_8_27_n425;
wire      [7:0] bv_8_28_n169;
wire      [7:0] bv_8_29_n97;
wire      [7:0] bv_8_2_n365;
wire      [7:0] bv_8_30_n68;
wire      [7:0] bv_8_31_n151;
wire      [7:0] bv_8_32_n401;
wire      [7:0] bv_8_33_n333;
wire      [7:0] bv_8_34_n280;
wire      [7:0] bv_8_35_n455;
wire      [7:0] bv_8_36_n238;
wire      [7:0] bv_8_37_n175;
wire      [7:0] bv_8_38_n472;
wire      [7:0] bv_8_39_n437;
wire      [7:0] bv_8_3_n122;
wire      [7:0] bv_8_40_n54;
wire      [7:0] bv_8_41_n414;
wire      [7:0] bv_8_42_n278;
wire      [7:0] bv_8_43_n466;
wire      [7:0] bv_8_44_n429;
wire      [7:0] bv_8_45_n18;
wire      [7:0] bv_8_46_n172;
wire      [7:0] bv_8_47_n411;
wire      [7:0] bv_8_48_n458;
wire      [7:0] bv_8_49_n456;
wire      [7:0] bv_8_4_n460;
wire      [7:0] bv_8_50_n252;
wire      [7:0] bv_8_51_n372;
wire      [7:0] bv_8_52_n450;
wire      [7:0] bv_8_53_n111;
wire      [7:0] bv_8_54_n446;
wire      [7:0] bv_8_55_n212;
wire      [7:0] bv_8_56_n341;
wire      [7:0] bv_8_57_n391;
wire      [7:0] bv_8_58_n250;
wire      [7:0] bv_8_59_n418;
wire      [7:0] bv_8_5_n448;
wire      [7:0] bv_8_60_n358;
wire      [7:0] bv_8_61_n300;
wire      [7:0] bv_8_62_n134;
wire      [7:0] bv_8_63_n433;
wire      [7:0] bv_8_64_n348;
wire      [7:0] bv_8_65_n24;
wire      [7:0] bv_8_66_n30;
wire      [7:0] bv_8_67_n376;
wire      [7:0] bv_8_68_n308;
wire      [7:0] bv_8_69_n368;
wire      [7:0] bv_8_6_n241;
wire      [7:0] bv_8_70_n270;
wire      [7:0] bv_8_71_n420;
wire      [7:0] bv_8_72_n125;
wire      [7:0] bv_8_73_n244;
wire      [7:0] bv_8_74_n388;
wire      [7:0] bv_8_75_n148;
wire      [7:0] bv_8_76_n386;
wire      [7:0] bv_8_77_n374;
wire      [7:0] bv_8_78_n203;
wire      [7:0] bv_8_79_n285;
wire      [7:0] bv_8_7_n444;
wire      [7:0] bv_8_80_n360;
wire      [7:0] bv_8_81_n352;
wire      [7:0] bv_8_82_n404;
wire      [7:0] bv_8_83_n402;
wire      [7:0] bv_8_84_n9;
wire      [7:0] bv_8_85_n57;
wire      [7:0] bv_8_86_n194;
wire      [7:0] bv_8_87_n109;
wire      [7:0] bv_8_88_n384;
wire      [7:0] bv_8_89_n394;
wire      [7:0] bv_8_8_n182;
wire      [7:0] bv_8_90_n392;
wire      [7:0] bv_8_91_n389;
wire      [7:0] bv_8_92_n236;
wire      [7:0] bv_8_93_n296;
wire      [7:0] bv_8_94_n261;
wire      [7:0] bv_8_95_n313;
wire      [7:0] bv_8_96_n289;
wire      [7:0] bv_8_97_n114;
wire      [7:0] bv_8_98_n228;
wire      [7:0] bv_8_99_n377;
wire      [7:0] bv_8_9_n432;
wire            clk;
wire            n102;
wire            n105;
wire            n108;
wire            n11;
wire            n110;
wire            n113;
wire            n116;
wire            n119;
wire            n121;
wire            n124;
wire            n127;
wire            n130;
wire            n133;
wire            n136;
wire            n139;
wire            n14;
wire            n141;
wire            n144;
wire            n147;
wire            n150;
wire            n153;
wire            n156;
wire            n158;
wire            n160;
wire            n162;
wire            n165;
wire            n168;
wire            n17;
wire            n171;
wire            n174;
wire            n176;
wire            n179;
wire            n181;
wire            n184;
wire            n186;
wire            n189;
wire            n191;
wire            n192;
wire            n193;
wire            n196;
wire            n199;
wire            n2;
wire            n20;
wire            n202;
wire            n204;
wire            n205;
wire            n208;
wire            n211;
wire            n214;
wire            n215;
wire            n217;
wire            n219;
wire            n221;
wire            n224;
wire            n227;
wire            n23;
wire            n230;
wire            n231;
wire            n233;
wire            n235;
wire            n237;
wire            n240;
wire            n243;
wire            n246;
wire            n249;
wire            n251;
wire            n254;
wire            n256;
wire            n257;
wire            n26;
wire            n260;
wire            n263;
wire            n264;
wire            n267;
wire            n268;
wire            n269;
wire            n272;
wire            n275;
wire            n277;
wire            n279;
wire            n282;
wire            n284;
wire            n286;
wire            n288;
wire            n29;
wire            n291;
wire            n293;
wire            n295;
wire            n297;
wire            n299;
wire            n301;
wire            n303;
wire            n304;
wire            n305;
wire            n307;
wire            n310;
wire            n312;
wire            n315;
wire            n317;
wire            n319;
wire            n32;
wire            n322;
wire            n324;
wire            n325;
wire            n327;
wire            n329;
wire            n332;
wire            n334;
wire            n335;
wire            n336;
wire            n338;
wire            n340;
wire            n343;
wire            n344;
wire            n345;
wire            n347;
wire            n35;
wire            n350;
wire            n351;
wire            n354;
wire            n356;
wire            n357;
wire            n359;
wire            n362;
wire            n364;
wire            n366;
wire            n367;
wire            n370;
wire            n371;
wire            n373;
wire            n375;
wire            n378;
wire            n379;
wire            n38;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n385;
wire            n387;
wire            n390;
wire            n393;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire            n399;
wire            n400;
wire            n403;
wire            n405;
wire            n407;
wire            n408;
wire            n409;
wire            n41;
wire            n410;
wire            n412;
wire            n413;
wire            n415;
wire            n416;
wire            n417;
wire            n419;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n426;
wire            n428;
wire            n430;
wire            n431;
wire            n434;
wire            n435;
wire            n436;
wire            n438;
wire            n439;
wire            n44;
wire            n440;
wire            n441;
wire            n443;
wire            n445;
wire            n447;
wire            n449;
wire            n451;
wire            n453;
wire            n454;
wire            n457;
wire            n459;
wire            n461;
wire            n463;
wire            n464;
wire            n465;
wire            n467;
wire            n468;
wire            n469;
wire            n47;
wire            n470;
wire            n471;
wire            n473;
wire            n474;
wire            n475;
wire            n476;
wire            n477;
wire            n478;
wire            n479;
wire            n480;
wire            n481;
wire            n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n490;
wire            n491;
wire            n492;
wire            n493;
wire            n494;
wire            n495;
wire            n496;
wire            n497;
wire            n498;
wire            n499;
wire            n5;
wire            n50;
wire            n500;
wire            n501;
wire            n502;
wire            n504;
wire            n505;
wire            n506;
wire            n507;
wire            n508;
wire            n509;
wire            n510;
wire            n511;
wire            n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire            n53;
wire      [7:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire      [7:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire      [7:0] n552;
wire      [7:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire            n56;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire      [7:0] n565;
wire      [7:0] n566;
wire      [7:0] n567;
wire      [7:0] n568;
wire      [7:0] n569;
wire      [7:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire      [7:0] n581;
wire      [7:0] n582;
wire      [7:0] n583;
wire      [7:0] n584;
wire      [7:0] n585;
wire      [7:0] n586;
wire      [7:0] n587;
wire      [7:0] n588;
wire      [7:0] n589;
wire            n59;
wire      [7:0] n590;
wire      [7:0] n591;
wire      [7:0] n592;
wire      [7:0] n593;
wire      [7:0] n594;
wire      [7:0] n595;
wire      [7:0] n596;
wire      [7:0] n597;
wire      [7:0] n598;
wire      [7:0] n599;
wire      [7:0] n600;
wire      [7:0] n601;
wire      [7:0] n602;
wire      [7:0] n603;
wire      [7:0] n604;
wire      [7:0] n605;
wire      [7:0] n606;
wire      [7:0] n607;
wire      [7:0] n608;
wire      [7:0] n609;
wire      [7:0] n610;
wire      [7:0] n611;
wire      [7:0] n612;
wire      [7:0] n613;
wire      [7:0] n614;
wire      [7:0] n615;
wire      [7:0] n616;
wire      [7:0] n617;
wire      [7:0] n618;
wire      [7:0] n619;
wire            n62;
wire      [7:0] n620;
wire      [7:0] n621;
wire      [7:0] n622;
wire      [7:0] n623;
wire      [7:0] n624;
wire      [7:0] n625;
wire      [7:0] n626;
wire      [7:0] n627;
wire      [7:0] n628;
wire      [7:0] n629;
wire      [7:0] n630;
wire      [7:0] n631;
wire      [7:0] n632;
wire      [7:0] n633;
wire      [7:0] n634;
wire      [7:0] n635;
wire      [7:0] n636;
wire      [7:0] n637;
wire      [7:0] n638;
wire      [7:0] n639;
wire      [7:0] n640;
wire      [7:0] n641;
wire      [7:0] n642;
wire      [7:0] n643;
wire      [7:0] n644;
wire      [7:0] n645;
wire      [7:0] n646;
wire      [7:0] n647;
wire      [7:0] n648;
wire      [7:0] n649;
wire            n65;
wire      [7:0] n650;
wire      [7:0] n651;
wire      [7:0] n652;
wire      [7:0] n653;
wire      [7:0] n654;
wire      [7:0] n655;
wire      [7:0] n656;
wire      [7:0] n657;
wire      [7:0] n658;
wire      [7:0] n659;
wire      [7:0] n660;
wire      [7:0] n661;
wire      [7:0] n662;
wire      [7:0] n663;
wire      [7:0] n664;
wire      [7:0] n665;
wire      [7:0] n666;
wire      [7:0] n667;
wire      [7:0] n668;
wire      [7:0] n669;
wire            n67;
wire      [7:0] n670;
wire      [7:0] n671;
wire      [7:0] n672;
wire      [7:0] n673;
wire      [7:0] n674;
wire      [7:0] n675;
wire      [7:0] n676;
wire      [7:0] n677;
wire      [7:0] n678;
wire      [7:0] n679;
wire      [7:0] n680;
wire      [7:0] n681;
wire      [7:0] n682;
wire      [7:0] n683;
wire      [7:0] n684;
wire      [7:0] n685;
wire      [7:0] n686;
wire      [7:0] n687;
wire      [7:0] n688;
wire      [7:0] n689;
wire      [7:0] n690;
wire      [7:0] n691;
wire      [7:0] n692;
wire      [7:0] n693;
wire      [7:0] n694;
wire      [7:0] n695;
wire      [7:0] n696;
wire      [7:0] n697;
wire      [7:0] n698;
wire      [7:0] n699;
wire            n70;
wire      [7:0] n700;
wire      [7:0] n701;
wire      [7:0] n702;
wire      [7:0] n703;
wire      [7:0] n704;
wire      [7:0] n705;
wire      [7:0] n706;
wire      [7:0] n707;
wire      [7:0] n708;
wire      [7:0] n709;
wire      [7:0] n710;
wire      [7:0] n711;
wire      [7:0] n712;
wire      [7:0] n713;
wire      [7:0] n714;
wire      [7:0] n715;
wire      [7:0] n716;
wire      [7:0] n717;
wire      [7:0] n718;
wire      [7:0] n719;
wire      [7:0] n720;
wire      [7:0] n721;
wire      [7:0] n722;
wire      [7:0] n723;
wire      [7:0] n724;
wire      [7:0] n725;
wire      [7:0] n726;
wire      [7:0] n727;
wire      [7:0] n728;
wire      [7:0] n729;
wire            n73;
wire      [7:0] n730;
wire      [7:0] n731;
wire      [7:0] n732;
wire      [7:0] n733;
wire      [7:0] n734;
wire      [7:0] n735;
wire      [7:0] n736;
wire      [7:0] n737;
wire      [7:0] n738;
wire      [7:0] n739;
wire      [7:0] n740;
wire      [7:0] n741;
wire      [7:0] n742;
wire      [7:0] n743;
wire      [7:0] n744;
wire      [7:0] n745;
wire      [7:0] n746;
wire      [7:0] n747;
wire      [7:0] n748;
wire      [7:0] n749;
wire            n75;
wire      [7:0] n750;
wire      [7:0] n751;
wire      [7:0] n752;
wire      [7:0] n753;
wire      [7:0] n754;
wire      [7:0] n755;
wire      [7:0] n756;
wire      [7:0] n757;
wire      [7:0] n758;
wire      [7:0] n759;
wire      [7:0] n760;
wire      [7:0] n761;
wire      [7:0] n762;
wire      [7:0] n763;
wire      [7:0] n764;
wire      [7:0] n765;
wire      [7:0] n766;
wire      [7:0] n767;
wire      [7:0] n768;
wire            n78;
wire            n8;
wire            n81;
wire            n84;
wire            n87;
wire            n90;
wire            n92;
wire            n93;
wire            n96;
wire            n99;
wire            rst;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign bv_8_255_n1 = 8'hff ;
assign n2 =  ( in ) == ( bv_8_255_n1 )  ;
assign bv_8_22_n3 = 8'h16 ;
assign bv_8_254_n4 = 8'hfe ;
assign n5 =  ( in ) == ( bv_8_254_n4 )  ;
assign bv_8_187_n6 = 8'hbb ;
assign bv_8_253_n7 = 8'hfd ;
assign n8 =  ( in ) == ( bv_8_253_n7 )  ;
assign bv_8_84_n9 = 8'h54 ;
assign bv_8_252_n10 = 8'hfc ;
assign n11 =  ( in ) == ( bv_8_252_n10 )  ;
assign bv_8_176_n12 = 8'hb0 ;
assign bv_8_251_n13 = 8'hfb ;
assign n14 =  ( in ) == ( bv_8_251_n13 )  ;
assign bv_8_15_n15 = 8'hf ;
assign bv_8_250_n16 = 8'hfa ;
assign n17 =  ( in ) == ( bv_8_250_n16 )  ;
assign bv_8_45_n18 = 8'h2d ;
assign bv_8_249_n19 = 8'hf9 ;
assign n20 =  ( in ) == ( bv_8_249_n19 )  ;
assign bv_8_153_n21 = 8'h99 ;
assign bv_8_248_n22 = 8'hf8 ;
assign n23 =  ( in ) == ( bv_8_248_n22 )  ;
assign bv_8_65_n24 = 8'h41 ;
assign bv_8_247_n25 = 8'hf7 ;
assign n26 =  ( in ) == ( bv_8_247_n25 )  ;
assign bv_8_104_n27 = 8'h68 ;
assign bv_8_246_n28 = 8'hf6 ;
assign n29 =  ( in ) == ( bv_8_246_n28 )  ;
assign bv_8_66_n30 = 8'h42 ;
assign bv_8_245_n31 = 8'hf5 ;
assign n32 =  ( in ) == ( bv_8_245_n31 )  ;
assign bv_8_230_n33 = 8'he6 ;
assign bv_8_244_n34 = 8'hf4 ;
assign n35 =  ( in ) == ( bv_8_244_n34 )  ;
assign bv_8_191_n36 = 8'hbf ;
assign bv_8_243_n37 = 8'hf3 ;
assign n38 =  ( in ) == ( bv_8_243_n37 )  ;
assign bv_8_13_n39 = 8'hd ;
assign bv_8_242_n40 = 8'hf2 ;
assign n41 =  ( in ) == ( bv_8_242_n40 )  ;
assign bv_8_137_n42 = 8'h89 ;
assign bv_8_241_n43 = 8'hf1 ;
assign n44 =  ( in ) == ( bv_8_241_n43 )  ;
assign bv_8_161_n45 = 8'ha1 ;
assign bv_8_240_n46 = 8'hf0 ;
assign n47 =  ( in ) == ( bv_8_240_n46 )  ;
assign bv_8_140_n48 = 8'h8c ;
assign bv_8_239_n49 = 8'hef ;
assign n50 =  ( in ) == ( bv_8_239_n49 )  ;
assign bv_8_223_n51 = 8'hdf ;
assign bv_8_238_n52 = 8'hee ;
assign n53 =  ( in ) == ( bv_8_238_n52 )  ;
assign bv_8_40_n54 = 8'h28 ;
assign bv_8_237_n55 = 8'hed ;
assign n56 =  ( in ) == ( bv_8_237_n55 )  ;
assign bv_8_85_n57 = 8'h55 ;
assign bv_8_236_n58 = 8'hec ;
assign n59 =  ( in ) == ( bv_8_236_n58 )  ;
assign bv_8_206_n60 = 8'hce ;
assign bv_8_235_n61 = 8'heb ;
assign n62 =  ( in ) == ( bv_8_235_n61 )  ;
assign bv_8_233_n63 = 8'he9 ;
assign bv_8_234_n64 = 8'hea ;
assign n65 =  ( in ) == ( bv_8_234_n64 )  ;
assign bv_8_135_n66 = 8'h87 ;
assign n67 =  ( in ) == ( bv_8_233_n63 )  ;
assign bv_8_30_n68 = 8'h1e ;
assign bv_8_232_n69 = 8'he8 ;
assign n70 =  ( in ) == ( bv_8_232_n69 )  ;
assign bv_8_155_n71 = 8'h9b ;
assign bv_8_231_n72 = 8'he7 ;
assign n73 =  ( in ) == ( bv_8_231_n72 )  ;
assign bv_8_148_n74 = 8'h94 ;
assign n75 =  ( in ) == ( bv_8_230_n33 )  ;
assign bv_8_142_n76 = 8'h8e ;
assign bv_8_229_n77 = 8'he5 ;
assign n78 =  ( in ) == ( bv_8_229_n77 )  ;
assign bv_8_217_n79 = 8'hd9 ;
assign bv_8_228_n80 = 8'he4 ;
assign n81 =  ( in ) == ( bv_8_228_n80 )  ;
assign bv_8_105_n82 = 8'h69 ;
assign bv_8_227_n83 = 8'he3 ;
assign n84 =  ( in ) == ( bv_8_227_n83 )  ;
assign bv_8_17_n85 = 8'h11 ;
assign bv_8_226_n86 = 8'he2 ;
assign n87 =  ( in ) == ( bv_8_226_n86 )  ;
assign bv_8_152_n88 = 8'h98 ;
assign bv_8_225_n89 = 8'he1 ;
assign n90 =  ( in ) == ( bv_8_225_n89 )  ;
assign bv_8_224_n91 = 8'he0 ;
assign n92 =  ( in ) == ( bv_8_224_n91 )  ;
assign n93 =  ( in ) == ( bv_8_223_n51 )  ;
assign bv_8_158_n94 = 8'h9e ;
assign bv_8_222_n95 = 8'hde ;
assign n96 =  ( in ) == ( bv_8_222_n95 )  ;
assign bv_8_29_n97 = 8'h1d ;
assign bv_8_221_n98 = 8'hdd ;
assign n99 =  ( in ) == ( bv_8_221_n98 )  ;
assign bv_8_193_n100 = 8'hc1 ;
assign bv_8_220_n101 = 8'hdc ;
assign n102 =  ( in ) == ( bv_8_220_n101 )  ;
assign bv_8_134_n103 = 8'h86 ;
assign bv_8_219_n104 = 8'hdb ;
assign n105 =  ( in ) == ( bv_8_219_n104 )  ;
assign bv_8_185_n106 = 8'hb9 ;
assign bv_8_218_n107 = 8'hda ;
assign n108 =  ( in ) == ( bv_8_218_n107 )  ;
assign bv_8_87_n109 = 8'h57 ;
assign n110 =  ( in ) == ( bv_8_217_n79 )  ;
assign bv_8_53_n111 = 8'h35 ;
assign bv_8_216_n112 = 8'hd8 ;
assign n113 =  ( in ) == ( bv_8_216_n112 )  ;
assign bv_8_97_n114 = 8'h61 ;
assign bv_8_215_n115 = 8'hd7 ;
assign n116 =  ( in ) == ( bv_8_215_n115 )  ;
assign bv_8_14_n117 = 8'he ;
assign bv_8_214_n118 = 8'hd6 ;
assign n119 =  ( in ) == ( bv_8_214_n118 )  ;
assign bv_8_213_n120 = 8'hd5 ;
assign n121 =  ( in ) == ( bv_8_213_n120 )  ;
assign bv_8_3_n122 = 8'h3 ;
assign bv_8_212_n123 = 8'hd4 ;
assign n124 =  ( in ) == ( bv_8_212_n123 )  ;
assign bv_8_72_n125 = 8'h48 ;
assign bv_8_211_n126 = 8'hd3 ;
assign n127 =  ( in ) == ( bv_8_211_n126 )  ;
assign bv_8_102_n128 = 8'h66 ;
assign bv_8_210_n129 = 8'hd2 ;
assign n130 =  ( in ) == ( bv_8_210_n129 )  ;
assign bv_8_181_n131 = 8'hb5 ;
assign bv_8_209_n132 = 8'hd1 ;
assign n133 =  ( in ) == ( bv_8_209_n132 )  ;
assign bv_8_62_n134 = 8'h3e ;
assign bv_8_208_n135 = 8'hd0 ;
assign n136 =  ( in ) == ( bv_8_208_n135 )  ;
assign bv_8_112_n137 = 8'h70 ;
assign bv_8_207_n138 = 8'hcf ;
assign n139 =  ( in ) == ( bv_8_207_n138 )  ;
assign bv_8_138_n140 = 8'h8a ;
assign n141 =  ( in ) == ( bv_8_206_n60 )  ;
assign bv_8_139_n142 = 8'h8b ;
assign bv_8_205_n143 = 8'hcd ;
assign n144 =  ( in ) == ( bv_8_205_n143 )  ;
assign bv_8_189_n145 = 8'hbd ;
assign bv_8_204_n146 = 8'hcc ;
assign n147 =  ( in ) == ( bv_8_204_n146 )  ;
assign bv_8_75_n148 = 8'h4b ;
assign bv_8_203_n149 = 8'hcb ;
assign n150 =  ( in ) == ( bv_8_203_n149 )  ;
assign bv_8_31_n151 = 8'h1f ;
assign bv_8_202_n152 = 8'hca ;
assign n153 =  ( in ) == ( bv_8_202_n152 )  ;
assign bv_8_116_n154 = 8'h74 ;
assign bv_8_201_n155 = 8'hc9 ;
assign n156 =  ( in ) == ( bv_8_201_n155 )  ;
assign bv_8_200_n157 = 8'hc8 ;
assign n158 =  ( in ) == ( bv_8_200_n157 )  ;
assign bv_8_199_n159 = 8'hc7 ;
assign n160 =  ( in ) == ( bv_8_199_n159 )  ;
assign bv_8_198_n161 = 8'hc6 ;
assign n162 =  ( in ) == ( bv_8_198_n161 )  ;
assign bv_8_180_n163 = 8'hb4 ;
assign bv_8_197_n164 = 8'hc5 ;
assign n165 =  ( in ) == ( bv_8_197_n164 )  ;
assign bv_8_166_n166 = 8'ha6 ;
assign bv_8_196_n167 = 8'hc4 ;
assign n168 =  ( in ) == ( bv_8_196_n167 )  ;
assign bv_8_28_n169 = 8'h1c ;
assign bv_8_195_n170 = 8'hc3 ;
assign n171 =  ( in ) == ( bv_8_195_n170 )  ;
assign bv_8_46_n172 = 8'h2e ;
assign bv_8_194_n173 = 8'hc2 ;
assign n174 =  ( in ) == ( bv_8_194_n173 )  ;
assign bv_8_37_n175 = 8'h25 ;
assign n176 =  ( in ) == ( bv_8_193_n100 )  ;
assign bv_8_120_n177 = 8'h78 ;
assign bv_8_192_n178 = 8'hc0 ;
assign n179 =  ( in ) == ( bv_8_192_n178 )  ;
assign bv_8_186_n180 = 8'hba ;
assign n181 =  ( in ) == ( bv_8_191_n36 )  ;
assign bv_8_8_n182 = 8'h8 ;
assign bv_8_190_n183 = 8'hbe ;
assign n184 =  ( in ) == ( bv_8_190_n183 )  ;
assign bv_8_174_n185 = 8'hae ;
assign n186 =  ( in ) == ( bv_8_189_n145 )  ;
assign bv_8_122_n187 = 8'h7a ;
assign bv_8_188_n188 = 8'hbc ;
assign n189 =  ( in ) == ( bv_8_188_n188 )  ;
assign bv_8_101_n190 = 8'h65 ;
assign n191 =  ( in ) == ( bv_8_187_n6 )  ;
assign n192 =  ( in ) == ( bv_8_186_n180 )  ;
assign n193 =  ( in ) == ( bv_8_185_n106 )  ;
assign bv_8_86_n194 = 8'h56 ;
assign bv_8_184_n195 = 8'hb8 ;
assign n196 =  ( in ) == ( bv_8_184_n195 )  ;
assign bv_8_108_n197 = 8'h6c ;
assign bv_8_183_n198 = 8'hb7 ;
assign n199 =  ( in ) == ( bv_8_183_n198 )  ;
assign bv_8_169_n200 = 8'ha9 ;
assign bv_8_182_n201 = 8'hb6 ;
assign n202 =  ( in ) == ( bv_8_182_n201 )  ;
assign bv_8_78_n203 = 8'h4e ;
assign n204 =  ( in ) == ( bv_8_181_n131 )  ;
assign n205 =  ( in ) == ( bv_8_180_n163 )  ;
assign bv_8_141_n206 = 8'h8d ;
assign bv_8_179_n207 = 8'hb3 ;
assign n208 =  ( in ) == ( bv_8_179_n207 )  ;
assign bv_8_109_n209 = 8'h6d ;
assign bv_8_178_n210 = 8'hb2 ;
assign n211 =  ( in ) == ( bv_8_178_n210 )  ;
assign bv_8_55_n212 = 8'h37 ;
assign bv_8_177_n213 = 8'hb1 ;
assign n214 =  ( in ) == ( bv_8_177_n213 )  ;
assign n215 =  ( in ) == ( bv_8_176_n12 )  ;
assign bv_8_175_n216 = 8'haf ;
assign n217 =  ( in ) == ( bv_8_175_n216 )  ;
assign bv_8_121_n218 = 8'h79 ;
assign n219 =  ( in ) == ( bv_8_174_n185 )  ;
assign bv_8_173_n220 = 8'had ;
assign n221 =  ( in ) == ( bv_8_173_n220 )  ;
assign bv_8_149_n222 = 8'h95 ;
assign bv_8_172_n223 = 8'hac ;
assign n224 =  ( in ) == ( bv_8_172_n223 )  ;
assign bv_8_145_n225 = 8'h91 ;
assign bv_8_171_n226 = 8'hab ;
assign n227 =  ( in ) == ( bv_8_171_n226 )  ;
assign bv_8_98_n228 = 8'h62 ;
assign bv_8_170_n229 = 8'haa ;
assign n230 =  ( in ) == ( bv_8_170_n229 )  ;
assign n231 =  ( in ) == ( bv_8_169_n200 )  ;
assign bv_8_168_n232 = 8'ha8 ;
assign n233 =  ( in ) == ( bv_8_168_n232 )  ;
assign bv_8_167_n234 = 8'ha7 ;
assign n235 =  ( in ) == ( bv_8_167_n234 )  ;
assign bv_8_92_n236 = 8'h5c ;
assign n237 =  ( in ) == ( bv_8_166_n166 )  ;
assign bv_8_36_n238 = 8'h24 ;
assign bv_8_165_n239 = 8'ha5 ;
assign n240 =  ( in ) == ( bv_8_165_n239 )  ;
assign bv_8_6_n241 = 8'h6 ;
assign bv_8_164_n242 = 8'ha4 ;
assign n243 =  ( in ) == ( bv_8_164_n242 )  ;
assign bv_8_73_n244 = 8'h49 ;
assign bv_8_163_n245 = 8'ha3 ;
assign n246 =  ( in ) == ( bv_8_163_n245 )  ;
assign bv_8_10_n247 = 8'ha ;
assign bv_8_162_n248 = 8'ha2 ;
assign n249 =  ( in ) == ( bv_8_162_n248 )  ;
assign bv_8_58_n250 = 8'h3a ;
assign n251 =  ( in ) == ( bv_8_161_n45 )  ;
assign bv_8_50_n252 = 8'h32 ;
assign bv_8_160_n253 = 8'ha0 ;
assign n254 =  ( in ) == ( bv_8_160_n253 )  ;
assign bv_8_159_n255 = 8'h9f ;
assign n256 =  ( in ) == ( bv_8_159_n255 )  ;
assign n257 =  ( in ) == ( bv_8_158_n94 )  ;
assign bv_8_11_n258 = 8'hb ;
assign bv_8_157_n259 = 8'h9d ;
assign n260 =  ( in ) == ( bv_8_157_n259 )  ;
assign bv_8_94_n261 = 8'h5e ;
assign bv_8_156_n262 = 8'h9c ;
assign n263 =  ( in ) == ( bv_8_156_n262 )  ;
assign n264 =  ( in ) == ( bv_8_155_n71 )  ;
assign bv_8_20_n265 = 8'h14 ;
assign bv_8_154_n266 = 8'h9a ;
assign n267 =  ( in ) == ( bv_8_154_n266 )  ;
assign n268 =  ( in ) == ( bv_8_153_n21 )  ;
assign n269 =  ( in ) == ( bv_8_152_n88 )  ;
assign bv_8_70_n270 = 8'h46 ;
assign bv_8_151_n271 = 8'h97 ;
assign n272 =  ( in ) == ( bv_8_151_n271 )  ;
assign bv_8_136_n273 = 8'h88 ;
assign bv_8_150_n274 = 8'h96 ;
assign n275 =  ( in ) == ( bv_8_150_n274 )  ;
assign bv_8_144_n276 = 8'h90 ;
assign n277 =  ( in ) == ( bv_8_149_n222 )  ;
assign bv_8_42_n278 = 8'h2a ;
assign n279 =  ( in ) == ( bv_8_148_n74 )  ;
assign bv_8_34_n280 = 8'h22 ;
assign bv_8_147_n281 = 8'h93 ;
assign n282 =  ( in ) == ( bv_8_147_n281 )  ;
assign bv_8_146_n283 = 8'h92 ;
assign n284 =  ( in ) == ( bv_8_146_n283 )  ;
assign bv_8_79_n285 = 8'h4f ;
assign n286 =  ( in ) == ( bv_8_145_n225 )  ;
assign bv_8_129_n287 = 8'h81 ;
assign n288 =  ( in ) == ( bv_8_144_n276 )  ;
assign bv_8_96_n289 = 8'h60 ;
assign bv_8_143_n290 = 8'h8f ;
assign n291 =  ( in ) == ( bv_8_143_n290 )  ;
assign bv_8_115_n292 = 8'h73 ;
assign n293 =  ( in ) == ( bv_8_142_n76 )  ;
assign bv_8_25_n294 = 8'h19 ;
assign n295 =  ( in ) == ( bv_8_141_n206 )  ;
assign bv_8_93_n296 = 8'h5d ;
assign n297 =  ( in ) == ( bv_8_140_n48 )  ;
assign bv_8_100_n298 = 8'h64 ;
assign n299 =  ( in ) == ( bv_8_139_n142 )  ;
assign bv_8_61_n300 = 8'h3d ;
assign n301 =  ( in ) == ( bv_8_138_n140 )  ;
assign bv_8_126_n302 = 8'h7e ;
assign n303 =  ( in ) == ( bv_8_137_n42 )  ;
assign n304 =  ( in ) == ( bv_8_136_n273 )  ;
assign n305 =  ( in ) == ( bv_8_135_n66 )  ;
assign bv_8_23_n306 = 8'h17 ;
assign n307 =  ( in ) == ( bv_8_134_n103 )  ;
assign bv_8_68_n308 = 8'h44 ;
assign bv_8_133_n309 = 8'h85 ;
assign n310 =  ( in ) == ( bv_8_133_n309 )  ;
assign bv_8_132_n311 = 8'h84 ;
assign n312 =  ( in ) == ( bv_8_132_n311 )  ;
assign bv_8_95_n313 = 8'h5f ;
assign bv_8_131_n314 = 8'h83 ;
assign n315 =  ( in ) == ( bv_8_131_n314 )  ;
assign bv_8_130_n316 = 8'h82 ;
assign n317 =  ( in ) == ( bv_8_130_n316 )  ;
assign bv_8_19_n318 = 8'h13 ;
assign n319 =  ( in ) == ( bv_8_129_n287 )  ;
assign bv_8_12_n320 = 8'hc ;
assign bv_8_128_n321 = 8'h80 ;
assign n322 =  ( in ) == ( bv_8_128_n321 )  ;
assign bv_8_127_n323 = 8'h7f ;
assign n324 =  ( in ) == ( bv_8_127_n323 )  ;
assign n325 =  ( in ) == ( bv_8_126_n302 )  ;
assign bv_8_125_n326 = 8'h7d ;
assign n327 =  ( in ) == ( bv_8_125_n326 )  ;
assign bv_8_124_n328 = 8'h7c ;
assign n329 =  ( in ) == ( bv_8_124_n328 )  ;
assign bv_8_16_n330 = 8'h10 ;
assign bv_8_123_n331 = 8'h7b ;
assign n332 =  ( in ) == ( bv_8_123_n331 )  ;
assign bv_8_33_n333 = 8'h21 ;
assign n334 =  ( in ) == ( bv_8_122_n187 )  ;
assign n335 =  ( in ) == ( bv_8_121_n218 )  ;
assign n336 =  ( in ) == ( bv_8_120_n177 )  ;
assign bv_8_119_n337 = 8'h77 ;
assign n338 =  ( in ) == ( bv_8_119_n337 )  ;
assign bv_8_118_n339 = 8'h76 ;
assign n340 =  ( in ) == ( bv_8_118_n339 )  ;
assign bv_8_56_n341 = 8'h38 ;
assign bv_8_117_n342 = 8'h75 ;
assign n343 =  ( in ) == ( bv_8_117_n342 )  ;
assign n344 =  ( in ) == ( bv_8_116_n154 )  ;
assign n345 =  ( in ) == ( bv_8_115_n292 )  ;
assign bv_8_114_n346 = 8'h72 ;
assign n347 =  ( in ) == ( bv_8_114_n346 )  ;
assign bv_8_64_n348 = 8'h40 ;
assign bv_8_113_n349 = 8'h71 ;
assign n350 =  ( in ) == ( bv_8_113_n349 )  ;
assign n351 =  ( in ) == ( bv_8_112_n137 )  ;
assign bv_8_81_n352 = 8'h51 ;
assign bv_8_111_n353 = 8'h6f ;
assign n354 =  ( in ) == ( bv_8_111_n353 )  ;
assign bv_8_110_n355 = 8'h6e ;
assign n356 =  ( in ) == ( bv_8_110_n355 )  ;
assign n357 =  ( in ) == ( bv_8_109_n209 )  ;
assign bv_8_60_n358 = 8'h3c ;
assign n359 =  ( in ) == ( bv_8_108_n197 )  ;
assign bv_8_80_n360 = 8'h50 ;
assign bv_8_107_n361 = 8'h6b ;
assign n362 =  ( in ) == ( bv_8_107_n361 )  ;
assign bv_8_106_n363 = 8'h6a ;
assign n364 =  ( in ) == ( bv_8_106_n363 )  ;
assign bv_8_2_n365 = 8'h2 ;
assign n366 =  ( in ) == ( bv_8_105_n82 )  ;
assign n367 =  ( in ) == ( bv_8_104_n27 )  ;
assign bv_8_69_n368 = 8'h45 ;
assign bv_8_103_n369 = 8'h67 ;
assign n370 =  ( in ) == ( bv_8_103_n369 )  ;
assign n371 =  ( in ) == ( bv_8_102_n128 )  ;
assign bv_8_51_n372 = 8'h33 ;
assign n373 =  ( in ) == ( bv_8_101_n190 )  ;
assign bv_8_77_n374 = 8'h4d ;
assign n375 =  ( in ) == ( bv_8_100_n298 )  ;
assign bv_8_67_n376 = 8'h43 ;
assign bv_8_99_n377 = 8'h63 ;
assign n378 =  ( in ) == ( bv_8_99_n377 )  ;
assign n379 =  ( in ) == ( bv_8_98_n228 )  ;
assign n380 =  ( in ) == ( bv_8_97_n114 )  ;
assign n381 =  ( in ) == ( bv_8_96_n289 )  ;
assign n382 =  ( in ) == ( bv_8_95_n313 )  ;
assign n383 =  ( in ) == ( bv_8_94_n261 )  ;
assign bv_8_88_n384 = 8'h58 ;
assign n385 =  ( in ) == ( bv_8_93_n296 )  ;
assign bv_8_76_n386 = 8'h4c ;
assign n387 =  ( in ) == ( bv_8_92_n236 )  ;
assign bv_8_74_n388 = 8'h4a ;
assign bv_8_91_n389 = 8'h5b ;
assign n390 =  ( in ) == ( bv_8_91_n389 )  ;
assign bv_8_57_n391 = 8'h39 ;
assign bv_8_90_n392 = 8'h5a ;
assign n393 =  ( in ) == ( bv_8_90_n392 )  ;
assign bv_8_89_n394 = 8'h59 ;
assign n395 =  ( in ) == ( bv_8_89_n394 )  ;
assign n396 =  ( in ) == ( bv_8_88_n384 )  ;
assign n397 =  ( in ) == ( bv_8_87_n109 )  ;
assign n398 =  ( in ) == ( bv_8_86_n194 )  ;
assign n399 =  ( in ) == ( bv_8_85_n57 )  ;
assign n400 =  ( in ) == ( bv_8_84_n9 )  ;
assign bv_8_32_n401 = 8'h20 ;
assign bv_8_83_n402 = 8'h53 ;
assign n403 =  ( in ) == ( bv_8_83_n402 )  ;
assign bv_8_82_n404 = 8'h52 ;
assign n405 =  ( in ) == ( bv_8_82_n404 )  ;
assign bv_8_0_n406 = 8'h0 ;
assign n407 =  ( in ) == ( bv_8_81_n352 )  ;
assign n408 =  ( in ) == ( bv_8_80_n360 )  ;
assign n409 =  ( in ) == ( bv_8_79_n285 )  ;
assign n410 =  ( in ) == ( bv_8_78_n203 )  ;
assign bv_8_47_n411 = 8'h2f ;
assign n412 =  ( in ) == ( bv_8_77_n374 )  ;
assign n413 =  ( in ) == ( bv_8_76_n386 )  ;
assign bv_8_41_n414 = 8'h29 ;
assign n415 =  ( in ) == ( bv_8_75_n148 )  ;
assign n416 =  ( in ) == ( bv_8_74_n388 )  ;
assign n417 =  ( in ) == ( bv_8_73_n244 )  ;
assign bv_8_59_n418 = 8'h3b ;
assign n419 =  ( in ) == ( bv_8_72_n125 )  ;
assign bv_8_71_n420 = 8'h47 ;
assign n421 =  ( in ) == ( bv_8_71_n420 )  ;
assign n422 =  ( in ) == ( bv_8_70_n270 )  ;
assign n423 =  ( in ) == ( bv_8_69_n368 )  ;
assign n424 =  ( in ) == ( bv_8_68_n308 )  ;
assign bv_8_27_n425 = 8'h1b ;
assign n426 =  ( in ) == ( bv_8_67_n376 )  ;
assign bv_8_26_n427 = 8'h1a ;
assign n428 =  ( in ) == ( bv_8_66_n30 )  ;
assign bv_8_44_n429 = 8'h2c ;
assign n430 =  ( in ) == ( bv_8_65_n24 )  ;
assign n431 =  ( in ) == ( bv_8_64_n348 )  ;
assign bv_8_9_n432 = 8'h9 ;
assign bv_8_63_n433 = 8'h3f ;
assign n434 =  ( in ) == ( bv_8_63_n433 )  ;
assign n435 =  ( in ) == ( bv_8_62_n134 )  ;
assign n436 =  ( in ) == ( bv_8_61_n300 )  ;
assign bv_8_39_n437 = 8'h27 ;
assign n438 =  ( in ) == ( bv_8_60_n358 )  ;
assign n439 =  ( in ) == ( bv_8_59_n418 )  ;
assign n440 =  ( in ) == ( bv_8_58_n250 )  ;
assign n441 =  ( in ) == ( bv_8_57_n391 )  ;
assign bv_8_18_n442 = 8'h12 ;
assign n443 =  ( in ) == ( bv_8_56_n341 )  ;
assign bv_8_7_n444 = 8'h7 ;
assign n445 =  ( in ) == ( bv_8_55_n212 )  ;
assign bv_8_54_n446 = 8'h36 ;
assign n447 =  ( in ) == ( bv_8_54_n446 )  ;
assign bv_8_5_n448 = 8'h5 ;
assign n449 =  ( in ) == ( bv_8_53_n111 )  ;
assign bv_8_52_n450 = 8'h34 ;
assign n451 =  ( in ) == ( bv_8_52_n450 )  ;
assign bv_8_24_n452 = 8'h18 ;
assign n453 =  ( in ) == ( bv_8_51_n372 )  ;
assign n454 =  ( in ) == ( bv_8_50_n252 )  ;
assign bv_8_35_n455 = 8'h23 ;
assign bv_8_49_n456 = 8'h31 ;
assign n457 =  ( in ) == ( bv_8_49_n456 )  ;
assign bv_8_48_n458 = 8'h30 ;
assign n459 =  ( in ) == ( bv_8_48_n458 )  ;
assign bv_8_4_n460 = 8'h4 ;
assign n461 =  ( in ) == ( bv_8_47_n411 )  ;
assign bv_8_21_n462 = 8'h15 ;
assign n463 =  ( in ) == ( bv_8_46_n172 )  ;
assign n464 =  ( in ) == ( bv_8_45_n18 )  ;
assign n465 =  ( in ) == ( bv_8_44_n429 )  ;
assign bv_8_43_n466 = 8'h2b ;
assign n467 =  ( in ) == ( bv_8_43_n466 )  ;
assign n468 =  ( in ) == ( bv_8_42_n278 )  ;
assign n469 =  ( in ) == ( bv_8_41_n414 )  ;
assign n470 =  ( in ) == ( bv_8_40_n54 )  ;
assign n471 =  ( in ) == ( bv_8_39_n437 )  ;
assign bv_8_38_n472 = 8'h26 ;
assign n473 =  ( in ) == ( bv_8_38_n472 )  ;
assign n474 =  ( in ) == ( bv_8_37_n175 )  ;
assign n475 =  ( in ) == ( bv_8_36_n238 )  ;
assign n476 =  ( in ) == ( bv_8_35_n455 )  ;
assign n477 =  ( in ) == ( bv_8_34_n280 )  ;
assign n478 =  ( in ) == ( bv_8_33_n333 )  ;
assign n479 =  ( in ) == ( bv_8_32_n401 )  ;
assign n480 =  ( in ) == ( bv_8_31_n151 )  ;
assign n481 =  ( in ) == ( bv_8_30_n68 )  ;
assign n482 =  ( in ) == ( bv_8_29_n97 )  ;
assign n483 =  ( in ) == ( bv_8_28_n169 )  ;
assign n484 =  ( in ) == ( bv_8_27_n425 )  ;
assign n485 =  ( in ) == ( bv_8_26_n427 )  ;
assign n486 =  ( in ) == ( bv_8_25_n294 )  ;
assign n487 =  ( in ) == ( bv_8_24_n452 )  ;
assign n488 =  ( in ) == ( bv_8_23_n306 )  ;
assign n489 =  ( in ) == ( bv_8_22_n3 )  ;
assign n490 =  ( in ) == ( bv_8_21_n462 )  ;
assign n491 =  ( in ) == ( bv_8_20_n265 )  ;
assign n492 =  ( in ) == ( bv_8_19_n318 )  ;
assign n493 =  ( in ) == ( bv_8_18_n442 )  ;
assign n494 =  ( in ) == ( bv_8_17_n85 )  ;
assign n495 =  ( in ) == ( bv_8_16_n330 )  ;
assign n496 =  ( in ) == ( bv_8_15_n15 )  ;
assign n497 =  ( in ) == ( bv_8_14_n117 )  ;
assign n498 =  ( in ) == ( bv_8_13_n39 )  ;
assign n499 =  ( in ) == ( bv_8_12_n320 )  ;
assign n500 =  ( in ) == ( bv_8_11_n258 )  ;
assign n501 =  ( in ) == ( bv_8_10_n247 )  ;
assign n502 =  ( in ) == ( bv_8_9_n432 )  ;
assign bv_8_1_n503 = 8'h1 ;
assign n504 =  ( in ) == ( bv_8_8_n182 )  ;
assign n505 =  ( in ) == ( bv_8_7_n444 )  ;
assign n506 =  ( in ) == ( bv_8_6_n241 )  ;
assign n507 =  ( in ) == ( bv_8_5_n448 )  ;
assign n508 =  ( in ) == ( bv_8_4_n460 )  ;
assign n509 =  ( in ) == ( bv_8_3_n122 )  ;
assign n510 =  ( in ) == ( bv_8_2_n365 )  ;
assign n511 =  ( in ) == ( bv_8_1_n503 )  ;
assign n512 =  ( in ) == ( bv_8_0_n406 )  ;
assign n513 =  ( n512 ) ? ( bv_8_99_n377 ) : ( out ) ;
assign n514 =  ( n511 ) ? ( bv_8_124_n328 ) : ( n513 ) ;
assign n515 =  ( n510 ) ? ( bv_8_119_n337 ) : ( n514 ) ;
assign n516 =  ( n509 ) ? ( bv_8_123_n331 ) : ( n515 ) ;
assign n517 =  ( n508 ) ? ( bv_8_242_n40 ) : ( n516 ) ;
assign n518 =  ( n507 ) ? ( bv_8_107_n361 ) : ( n517 ) ;
assign n519 =  ( n506 ) ? ( bv_8_111_n353 ) : ( n518 ) ;
assign n520 =  ( n505 ) ? ( bv_8_197_n164 ) : ( n519 ) ;
assign n521 =  ( n504 ) ? ( bv_8_48_n458 ) : ( n520 ) ;
assign n522 =  ( n502 ) ? ( bv_8_1_n503 ) : ( n521 ) ;
assign n523 =  ( n501 ) ? ( bv_8_103_n369 ) : ( n522 ) ;
assign n524 =  ( n500 ) ? ( bv_8_43_n466 ) : ( n523 ) ;
assign n525 =  ( n499 ) ? ( bv_8_254_n4 ) : ( n524 ) ;
assign n526 =  ( n498 ) ? ( bv_8_215_n115 ) : ( n525 ) ;
assign n527 =  ( n497 ) ? ( bv_8_171_n226 ) : ( n526 ) ;
assign n528 =  ( n496 ) ? ( bv_8_118_n339 ) : ( n527 ) ;
assign n529 =  ( n495 ) ? ( bv_8_202_n152 ) : ( n528 ) ;
assign n530 =  ( n494 ) ? ( bv_8_130_n316 ) : ( n529 ) ;
assign n531 =  ( n493 ) ? ( bv_8_201_n155 ) : ( n530 ) ;
assign n532 =  ( n492 ) ? ( bv_8_125_n326 ) : ( n531 ) ;
assign n533 =  ( n491 ) ? ( bv_8_250_n16 ) : ( n532 ) ;
assign n534 =  ( n490 ) ? ( bv_8_89_n394 ) : ( n533 ) ;
assign n535 =  ( n489 ) ? ( bv_8_71_n420 ) : ( n534 ) ;
assign n536 =  ( n488 ) ? ( bv_8_240_n46 ) : ( n535 ) ;
assign n537 =  ( n487 ) ? ( bv_8_173_n220 ) : ( n536 ) ;
assign n538 =  ( n486 ) ? ( bv_8_212_n123 ) : ( n537 ) ;
assign n539 =  ( n485 ) ? ( bv_8_162_n248 ) : ( n538 ) ;
assign n540 =  ( n484 ) ? ( bv_8_175_n216 ) : ( n539 ) ;
assign n541 =  ( n483 ) ? ( bv_8_156_n262 ) : ( n540 ) ;
assign n542 =  ( n482 ) ? ( bv_8_164_n242 ) : ( n541 ) ;
assign n543 =  ( n481 ) ? ( bv_8_114_n346 ) : ( n542 ) ;
assign n544 =  ( n480 ) ? ( bv_8_192_n178 ) : ( n543 ) ;
assign n545 =  ( n479 ) ? ( bv_8_183_n198 ) : ( n544 ) ;
assign n546 =  ( n478 ) ? ( bv_8_253_n7 ) : ( n545 ) ;
assign n547 =  ( n477 ) ? ( bv_8_147_n281 ) : ( n546 ) ;
assign n548 =  ( n476 ) ? ( bv_8_38_n472 ) : ( n547 ) ;
assign n549 =  ( n475 ) ? ( bv_8_54_n446 ) : ( n548 ) ;
assign n550 =  ( n474 ) ? ( bv_8_63_n433 ) : ( n549 ) ;
assign n551 =  ( n473 ) ? ( bv_8_247_n25 ) : ( n550 ) ;
assign n552 =  ( n471 ) ? ( bv_8_204_n146 ) : ( n551 ) ;
assign n553 =  ( n470 ) ? ( bv_8_52_n450 ) : ( n552 ) ;
assign n554 =  ( n469 ) ? ( bv_8_165_n239 ) : ( n553 ) ;
assign n555 =  ( n468 ) ? ( bv_8_229_n77 ) : ( n554 ) ;
assign n556 =  ( n467 ) ? ( bv_8_241_n43 ) : ( n555 ) ;
assign n557 =  ( n465 ) ? ( bv_8_113_n349 ) : ( n556 ) ;
assign n558 =  ( n464 ) ? ( bv_8_216_n112 ) : ( n557 ) ;
assign n559 =  ( n463 ) ? ( bv_8_49_n456 ) : ( n558 ) ;
assign n560 =  ( n461 ) ? ( bv_8_21_n462 ) : ( n559 ) ;
assign n561 =  ( n459 ) ? ( bv_8_4_n460 ) : ( n560 ) ;
assign n562 =  ( n457 ) ? ( bv_8_199_n159 ) : ( n561 ) ;
assign n563 =  ( n454 ) ? ( bv_8_35_n455 ) : ( n562 ) ;
assign n564 =  ( n453 ) ? ( bv_8_195_n170 ) : ( n563 ) ;
assign n565 =  ( n451 ) ? ( bv_8_24_n452 ) : ( n564 ) ;
assign n566 =  ( n449 ) ? ( bv_8_150_n274 ) : ( n565 ) ;
assign n567 =  ( n447 ) ? ( bv_8_5_n448 ) : ( n566 ) ;
assign n568 =  ( n445 ) ? ( bv_8_154_n266 ) : ( n567 ) ;
assign n569 =  ( n443 ) ? ( bv_8_7_n444 ) : ( n568 ) ;
assign n570 =  ( n441 ) ? ( bv_8_18_n442 ) : ( n569 ) ;
assign n571 =  ( n440 ) ? ( bv_8_128_n321 ) : ( n570 ) ;
assign n572 =  ( n439 ) ? ( bv_8_226_n86 ) : ( n571 ) ;
assign n573 =  ( n438 ) ? ( bv_8_235_n61 ) : ( n572 ) ;
assign n574 =  ( n436 ) ? ( bv_8_39_n437 ) : ( n573 ) ;
assign n575 =  ( n435 ) ? ( bv_8_178_n210 ) : ( n574 ) ;
assign n576 =  ( n434 ) ? ( bv_8_117_n342 ) : ( n575 ) ;
assign n577 =  ( n431 ) ? ( bv_8_9_n432 ) : ( n576 ) ;
assign n578 =  ( n430 ) ? ( bv_8_131_n314 ) : ( n577 ) ;
assign n579 =  ( n428 ) ? ( bv_8_44_n429 ) : ( n578 ) ;
assign n580 =  ( n426 ) ? ( bv_8_26_n427 ) : ( n579 ) ;
assign n581 =  ( n424 ) ? ( bv_8_27_n425 ) : ( n580 ) ;
assign n582 =  ( n423 ) ? ( bv_8_110_n355 ) : ( n581 ) ;
assign n583 =  ( n422 ) ? ( bv_8_90_n392 ) : ( n582 ) ;
assign n584 =  ( n421 ) ? ( bv_8_160_n253 ) : ( n583 ) ;
assign n585 =  ( n419 ) ? ( bv_8_82_n404 ) : ( n584 ) ;
assign n586 =  ( n417 ) ? ( bv_8_59_n418 ) : ( n585 ) ;
assign n587 =  ( n416 ) ? ( bv_8_214_n118 ) : ( n586 ) ;
assign n588 =  ( n415 ) ? ( bv_8_179_n207 ) : ( n587 ) ;
assign n589 =  ( n413 ) ? ( bv_8_41_n414 ) : ( n588 ) ;
assign n590 =  ( n412 ) ? ( bv_8_227_n83 ) : ( n589 ) ;
assign n591 =  ( n410 ) ? ( bv_8_47_n411 ) : ( n590 ) ;
assign n592 =  ( n409 ) ? ( bv_8_132_n311 ) : ( n591 ) ;
assign n593 =  ( n408 ) ? ( bv_8_83_n402 ) : ( n592 ) ;
assign n594 =  ( n407 ) ? ( bv_8_209_n132 ) : ( n593 ) ;
assign n595 =  ( n405 ) ? ( bv_8_0_n406 ) : ( n594 ) ;
assign n596 =  ( n403 ) ? ( bv_8_237_n55 ) : ( n595 ) ;
assign n597 =  ( n400 ) ? ( bv_8_32_n401 ) : ( n596 ) ;
assign n598 =  ( n399 ) ? ( bv_8_252_n10 ) : ( n597 ) ;
assign n599 =  ( n398 ) ? ( bv_8_177_n213 ) : ( n598 ) ;
assign n600 =  ( n397 ) ? ( bv_8_91_n389 ) : ( n599 ) ;
assign n601 =  ( n396 ) ? ( bv_8_106_n363 ) : ( n600 ) ;
assign n602 =  ( n395 ) ? ( bv_8_203_n149 ) : ( n601 ) ;
assign n603 =  ( n393 ) ? ( bv_8_190_n183 ) : ( n602 ) ;
assign n604 =  ( n390 ) ? ( bv_8_57_n391 ) : ( n603 ) ;
assign n605 =  ( n387 ) ? ( bv_8_74_n388 ) : ( n604 ) ;
assign n606 =  ( n385 ) ? ( bv_8_76_n386 ) : ( n605 ) ;
assign n607 =  ( n383 ) ? ( bv_8_88_n384 ) : ( n606 ) ;
assign n608 =  ( n382 ) ? ( bv_8_207_n138 ) : ( n607 ) ;
assign n609 =  ( n381 ) ? ( bv_8_208_n135 ) : ( n608 ) ;
assign n610 =  ( n380 ) ? ( bv_8_239_n49 ) : ( n609 ) ;
assign n611 =  ( n379 ) ? ( bv_8_170_n229 ) : ( n610 ) ;
assign n612 =  ( n378 ) ? ( bv_8_251_n13 ) : ( n611 ) ;
assign n613 =  ( n375 ) ? ( bv_8_67_n376 ) : ( n612 ) ;
assign n614 =  ( n373 ) ? ( bv_8_77_n374 ) : ( n613 ) ;
assign n615 =  ( n371 ) ? ( bv_8_51_n372 ) : ( n614 ) ;
assign n616 =  ( n370 ) ? ( bv_8_133_n309 ) : ( n615 ) ;
assign n617 =  ( n367 ) ? ( bv_8_69_n368 ) : ( n616 ) ;
assign n618 =  ( n366 ) ? ( bv_8_249_n19 ) : ( n617 ) ;
assign n619 =  ( n364 ) ? ( bv_8_2_n365 ) : ( n618 ) ;
assign n620 =  ( n362 ) ? ( bv_8_127_n323 ) : ( n619 ) ;
assign n621 =  ( n359 ) ? ( bv_8_80_n360 ) : ( n620 ) ;
assign n622 =  ( n357 ) ? ( bv_8_60_n358 ) : ( n621 ) ;
assign n623 =  ( n356 ) ? ( bv_8_159_n255 ) : ( n622 ) ;
assign n624 =  ( n354 ) ? ( bv_8_168_n232 ) : ( n623 ) ;
assign n625 =  ( n351 ) ? ( bv_8_81_n352 ) : ( n624 ) ;
assign n626 =  ( n350 ) ? ( bv_8_163_n245 ) : ( n625 ) ;
assign n627 =  ( n347 ) ? ( bv_8_64_n348 ) : ( n626 ) ;
assign n628 =  ( n345 ) ? ( bv_8_143_n290 ) : ( n627 ) ;
assign n629 =  ( n344 ) ? ( bv_8_146_n283 ) : ( n628 ) ;
assign n630 =  ( n343 ) ? ( bv_8_157_n259 ) : ( n629 ) ;
assign n631 =  ( n340 ) ? ( bv_8_56_n341 ) : ( n630 ) ;
assign n632 =  ( n338 ) ? ( bv_8_245_n31 ) : ( n631 ) ;
assign n633 =  ( n336 ) ? ( bv_8_188_n188 ) : ( n632 ) ;
assign n634 =  ( n335 ) ? ( bv_8_182_n201 ) : ( n633 ) ;
assign n635 =  ( n334 ) ? ( bv_8_218_n107 ) : ( n634 ) ;
assign n636 =  ( n332 ) ? ( bv_8_33_n333 ) : ( n635 ) ;
assign n637 =  ( n329 ) ? ( bv_8_16_n330 ) : ( n636 ) ;
assign n638 =  ( n327 ) ? ( bv_8_255_n1 ) : ( n637 ) ;
assign n639 =  ( n325 ) ? ( bv_8_243_n37 ) : ( n638 ) ;
assign n640 =  ( n324 ) ? ( bv_8_210_n129 ) : ( n639 ) ;
assign n641 =  ( n322 ) ? ( bv_8_205_n143 ) : ( n640 ) ;
assign n642 =  ( n319 ) ? ( bv_8_12_n320 ) : ( n641 ) ;
assign n643 =  ( n317 ) ? ( bv_8_19_n318 ) : ( n642 ) ;
assign n644 =  ( n315 ) ? ( bv_8_236_n58 ) : ( n643 ) ;
assign n645 =  ( n312 ) ? ( bv_8_95_n313 ) : ( n644 ) ;
assign n646 =  ( n310 ) ? ( bv_8_151_n271 ) : ( n645 ) ;
assign n647 =  ( n307 ) ? ( bv_8_68_n308 ) : ( n646 ) ;
assign n648 =  ( n305 ) ? ( bv_8_23_n306 ) : ( n647 ) ;
assign n649 =  ( n304 ) ? ( bv_8_196_n167 ) : ( n648 ) ;
assign n650 =  ( n303 ) ? ( bv_8_167_n234 ) : ( n649 ) ;
assign n651 =  ( n301 ) ? ( bv_8_126_n302 ) : ( n650 ) ;
assign n652 =  ( n299 ) ? ( bv_8_61_n300 ) : ( n651 ) ;
assign n653 =  ( n297 ) ? ( bv_8_100_n298 ) : ( n652 ) ;
assign n654 =  ( n295 ) ? ( bv_8_93_n296 ) : ( n653 ) ;
assign n655 =  ( n293 ) ? ( bv_8_25_n294 ) : ( n654 ) ;
assign n656 =  ( n291 ) ? ( bv_8_115_n292 ) : ( n655 ) ;
assign n657 =  ( n288 ) ? ( bv_8_96_n289 ) : ( n656 ) ;
assign n658 =  ( n286 ) ? ( bv_8_129_n287 ) : ( n657 ) ;
assign n659 =  ( n284 ) ? ( bv_8_79_n285 ) : ( n658 ) ;
assign n660 =  ( n282 ) ? ( bv_8_220_n101 ) : ( n659 ) ;
assign n661 =  ( n279 ) ? ( bv_8_34_n280 ) : ( n660 ) ;
assign n662 =  ( n277 ) ? ( bv_8_42_n278 ) : ( n661 ) ;
assign n663 =  ( n275 ) ? ( bv_8_144_n276 ) : ( n662 ) ;
assign n664 =  ( n272 ) ? ( bv_8_136_n273 ) : ( n663 ) ;
assign n665 =  ( n269 ) ? ( bv_8_70_n270 ) : ( n664 ) ;
assign n666 =  ( n268 ) ? ( bv_8_238_n52 ) : ( n665 ) ;
assign n667 =  ( n267 ) ? ( bv_8_184_n195 ) : ( n666 ) ;
assign n668 =  ( n264 ) ? ( bv_8_20_n265 ) : ( n667 ) ;
assign n669 =  ( n263 ) ? ( bv_8_222_n95 ) : ( n668 ) ;
assign n670 =  ( n260 ) ? ( bv_8_94_n261 ) : ( n669 ) ;
assign n671 =  ( n257 ) ? ( bv_8_11_n258 ) : ( n670 ) ;
assign n672 =  ( n256 ) ? ( bv_8_219_n104 ) : ( n671 ) ;
assign n673 =  ( n254 ) ? ( bv_8_224_n91 ) : ( n672 ) ;
assign n674 =  ( n251 ) ? ( bv_8_50_n252 ) : ( n673 ) ;
assign n675 =  ( n249 ) ? ( bv_8_58_n250 ) : ( n674 ) ;
assign n676 =  ( n246 ) ? ( bv_8_10_n247 ) : ( n675 ) ;
assign n677 =  ( n243 ) ? ( bv_8_73_n244 ) : ( n676 ) ;
assign n678 =  ( n240 ) ? ( bv_8_6_n241 ) : ( n677 ) ;
assign n679 =  ( n237 ) ? ( bv_8_36_n238 ) : ( n678 ) ;
assign n680 =  ( n235 ) ? ( bv_8_92_n236 ) : ( n679 ) ;
assign n681 =  ( n233 ) ? ( bv_8_194_n173 ) : ( n680 ) ;
assign n682 =  ( n231 ) ? ( bv_8_211_n126 ) : ( n681 ) ;
assign n683 =  ( n230 ) ? ( bv_8_172_n223 ) : ( n682 ) ;
assign n684 =  ( n227 ) ? ( bv_8_98_n228 ) : ( n683 ) ;
assign n685 =  ( n224 ) ? ( bv_8_145_n225 ) : ( n684 ) ;
assign n686 =  ( n221 ) ? ( bv_8_149_n222 ) : ( n685 ) ;
assign n687 =  ( n219 ) ? ( bv_8_228_n80 ) : ( n686 ) ;
assign n688 =  ( n217 ) ? ( bv_8_121_n218 ) : ( n687 ) ;
assign n689 =  ( n215 ) ? ( bv_8_231_n72 ) : ( n688 ) ;
assign n690 =  ( n214 ) ? ( bv_8_200_n157 ) : ( n689 ) ;
assign n691 =  ( n211 ) ? ( bv_8_55_n212 ) : ( n690 ) ;
assign n692 =  ( n208 ) ? ( bv_8_109_n209 ) : ( n691 ) ;
assign n693 =  ( n205 ) ? ( bv_8_141_n206 ) : ( n692 ) ;
assign n694 =  ( n204 ) ? ( bv_8_213_n120 ) : ( n693 ) ;
assign n695 =  ( n202 ) ? ( bv_8_78_n203 ) : ( n694 ) ;
assign n696 =  ( n199 ) ? ( bv_8_169_n200 ) : ( n695 ) ;
assign n697 =  ( n196 ) ? ( bv_8_108_n197 ) : ( n696 ) ;
assign n698 =  ( n193 ) ? ( bv_8_86_n194 ) : ( n697 ) ;
assign n699 =  ( n192 ) ? ( bv_8_244_n34 ) : ( n698 ) ;
assign n700 =  ( n191 ) ? ( bv_8_234_n64 ) : ( n699 ) ;
assign n701 =  ( n189 ) ? ( bv_8_101_n190 ) : ( n700 ) ;
assign n702 =  ( n186 ) ? ( bv_8_122_n187 ) : ( n701 ) ;
assign n703 =  ( n184 ) ? ( bv_8_174_n185 ) : ( n702 ) ;
assign n704 =  ( n181 ) ? ( bv_8_8_n182 ) : ( n703 ) ;
assign n705 =  ( n179 ) ? ( bv_8_186_n180 ) : ( n704 ) ;
assign n706 =  ( n176 ) ? ( bv_8_120_n177 ) : ( n705 ) ;
assign n707 =  ( n174 ) ? ( bv_8_37_n175 ) : ( n706 ) ;
assign n708 =  ( n171 ) ? ( bv_8_46_n172 ) : ( n707 ) ;
assign n709 =  ( n168 ) ? ( bv_8_28_n169 ) : ( n708 ) ;
assign n710 =  ( n165 ) ? ( bv_8_166_n166 ) : ( n709 ) ;
assign n711 =  ( n162 ) ? ( bv_8_180_n163 ) : ( n710 ) ;
assign n712 =  ( n160 ) ? ( bv_8_198_n161 ) : ( n711 ) ;
assign n713 =  ( n158 ) ? ( bv_8_232_n69 ) : ( n712 ) ;
assign n714 =  ( n156 ) ? ( bv_8_221_n98 ) : ( n713 ) ;
assign n715 =  ( n153 ) ? ( bv_8_116_n154 ) : ( n714 ) ;
assign n716 =  ( n150 ) ? ( bv_8_31_n151 ) : ( n715 ) ;
assign n717 =  ( n147 ) ? ( bv_8_75_n148 ) : ( n716 ) ;
assign n718 =  ( n144 ) ? ( bv_8_189_n145 ) : ( n717 ) ;
assign n719 =  ( n141 ) ? ( bv_8_139_n142 ) : ( n718 ) ;
assign n720 =  ( n139 ) ? ( bv_8_138_n140 ) : ( n719 ) ;
assign n721 =  ( n136 ) ? ( bv_8_112_n137 ) : ( n720 ) ;
assign n722 =  ( n133 ) ? ( bv_8_62_n134 ) : ( n721 ) ;
assign n723 =  ( n130 ) ? ( bv_8_181_n131 ) : ( n722 ) ;
assign n724 =  ( n127 ) ? ( bv_8_102_n128 ) : ( n723 ) ;
assign n725 =  ( n124 ) ? ( bv_8_72_n125 ) : ( n724 ) ;
assign n726 =  ( n121 ) ? ( bv_8_3_n122 ) : ( n725 ) ;
assign n727 =  ( n119 ) ? ( bv_8_246_n28 ) : ( n726 ) ;
assign n728 =  ( n116 ) ? ( bv_8_14_n117 ) : ( n727 ) ;
assign n729 =  ( n113 ) ? ( bv_8_97_n114 ) : ( n728 ) ;
assign n730 =  ( n110 ) ? ( bv_8_53_n111 ) : ( n729 ) ;
assign n731 =  ( n108 ) ? ( bv_8_87_n109 ) : ( n730 ) ;
assign n732 =  ( n105 ) ? ( bv_8_185_n106 ) : ( n731 ) ;
assign n733 =  ( n102 ) ? ( bv_8_134_n103 ) : ( n732 ) ;
assign n734 =  ( n99 ) ? ( bv_8_193_n100 ) : ( n733 ) ;
assign n735 =  ( n96 ) ? ( bv_8_29_n97 ) : ( n734 ) ;
assign n736 =  ( n93 ) ? ( bv_8_158_n94 ) : ( n735 ) ;
assign n737 =  ( n92 ) ? ( bv_8_225_n89 ) : ( n736 ) ;
assign n738 =  ( n90 ) ? ( bv_8_248_n22 ) : ( n737 ) ;
assign n739 =  ( n87 ) ? ( bv_8_152_n88 ) : ( n738 ) ;
assign n740 =  ( n84 ) ? ( bv_8_17_n85 ) : ( n739 ) ;
assign n741 =  ( n81 ) ? ( bv_8_105_n82 ) : ( n740 ) ;
assign n742 =  ( n78 ) ? ( bv_8_217_n79 ) : ( n741 ) ;
assign n743 =  ( n75 ) ? ( bv_8_142_n76 ) : ( n742 ) ;
assign n744 =  ( n73 ) ? ( bv_8_148_n74 ) : ( n743 ) ;
assign n745 =  ( n70 ) ? ( bv_8_155_n71 ) : ( n744 ) ;
assign n746 =  ( n67 ) ? ( bv_8_30_n68 ) : ( n745 ) ;
assign n747 =  ( n65 ) ? ( bv_8_135_n66 ) : ( n746 ) ;
assign n748 =  ( n62 ) ? ( bv_8_233_n63 ) : ( n747 ) ;
assign n749 =  ( n59 ) ? ( bv_8_206_n60 ) : ( n748 ) ;
assign n750 =  ( n56 ) ? ( bv_8_85_n57 ) : ( n749 ) ;
assign n751 =  ( n53 ) ? ( bv_8_40_n54 ) : ( n750 ) ;
assign n752 =  ( n50 ) ? ( bv_8_223_n51 ) : ( n751 ) ;
assign n753 =  ( n47 ) ? ( bv_8_140_n48 ) : ( n752 ) ;
assign n754 =  ( n44 ) ? ( bv_8_161_n45 ) : ( n753 ) ;
assign n755 =  ( n41 ) ? ( bv_8_137_n42 ) : ( n754 ) ;
assign n756 =  ( n38 ) ? ( bv_8_13_n39 ) : ( n755 ) ;
assign n757 =  ( n35 ) ? ( bv_8_191_n36 ) : ( n756 ) ;
assign n758 =  ( n32 ) ? ( bv_8_230_n33 ) : ( n757 ) ;
assign n759 =  ( n29 ) ? ( bv_8_66_n30 ) : ( n758 ) ;
assign n760 =  ( n26 ) ? ( bv_8_104_n27 ) : ( n759 ) ;
assign n761 =  ( n23 ) ? ( bv_8_65_n24 ) : ( n760 ) ;
assign n762 =  ( n20 ) ? ( bv_8_153_n21 ) : ( n761 ) ;
assign n763 =  ( n17 ) ? ( bv_8_45_n18 ) : ( n762 ) ;
assign n764 =  ( n14 ) ? ( bv_8_15_n15 ) : ( n763 ) ;
assign n765 =  ( n11 ) ? ( bv_8_176_n12 ) : ( n764 ) ;
assign n766 =  ( n8 ) ? ( bv_8_84_n9 ) : ( n765 ) ;
assign n767 =  ( n5 ) ? ( bv_8_187_n6 ) : ( n766 ) ;
assign n768 =  ( n2 ) ? ( bv_8_22_n3 ) : ( n767 ) ;
always @(posedge clk) begin
   if(rst) begin
       __COUNTER_start__n0 <= 0;
   end
   else if(__ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           in <= in ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           out <= n768 ;
       end
   end
end
endmodule
