module \$paramod\CDP_ICVT_mgc_in_wire_v1\rscid=5\width=2 (d, z);
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:78" *)
  output [1:0] d;
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:79" *)
  input [1:0] z;
  assign d = z;
endmodule
