module NV_NVDLA_CMAC_CORE_MAC_nan(nvdla_core_clk, nvdla_core_rstn, cfg_is_fp16, cfg_reg_en, dat_actv_data, dat_actv_nan, wt_actv_data, wt_actv_nan, out_nan_mts, out_nan_pvld);
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:308" *)
  wire [32:0] _000_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1086" *)
  wire _001_;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:23" *)
  input cfg_is_fp16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:31" *)
  reg [32:0] cfg_is_fp16_d1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:24" *)
  input cfg_reg_en;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:32" *)
  (* unused_bits = "0 1 2 13 14 16 17 18 29 30 32 33 34 45 46 48 49 50 61 62 64 65 66 77 78 80 81 82 93 94 96 97 98 109 110 112 113 114 125 126 128 129 130 141 142 144 145 146 157 158 160 161 162 173 174 176 177 178 189 190 192 193 194 205 206 208 209 210 221 222 224 225 226 237 238 240 241 242 253 254 256 257 258 269 270 272 273 274 285 286 288 289 290 301 302 304 305 306 317 318 320 321 322 333 334 336 337 338 349 350 352 353 354 365 366 368 369 370 381 382 384 385 386 397 398 400 401 402 413 414 416 417 418 429 430 432 433 434 445 446 448 449 450 461 462 464 465 466 477 478 480 481 482 493 494 496 497 498 509 510 512 513 514 525 526 528 529 530 541 542 544 545 546 557 558 560 561 562 573 574 576 577 578 589 590 592 593 594 605 606 608 609 610 621 622 624 625 626 637 638 640 641 642 653 654 656 657 658 669 670 672 673 674 685 686 688 689 690 701 702 704 705 706 717 718 720 721 722 733 734 736 737 738 749 750 752 753 754 765 766 768 769 770 781 782 784 785 786 797 798 800 801 802 813 814 816 817 818 829 830 832 833 834 845 846 848 849 850 861 862 864 865 866 877 878 880 881 882 893 894 896 897 898 909 910 912 913 914 925 926 928 929 930 941 942 944 945 946 957 958 960 961 962 973 974 976 977 978 989 990 992 993 994 1005 1006 1008 1009 1010 1021 1022 1024 1025 1026 1037 1038 1040 1041 1042 1053 1054 1056 1057 1058 1069 1070 1072 1073 1074 1085 1086 1088 1089 1090 1101 1102 1104 1105 1106 1117 1118 1120 1121 1122 1133 1134 1136 1137 1138 1149 1150 1152 1153 1154 1165 1166 1168 1169 1170 1181 1182 1184 1185 1186 1197 1198 1200 1201 1202 1213 1214 1216 1217 1218 1229 1230 1232 1233 1234 1245 1246 1248 1249 1250 1261 1262 1264 1265 1266 1277 1278 1280 1281 1282 1293 1294 1296 1297 1298 1309 1310 1312 1313 1314 1325 1326 1328 1329 1330 1341 1342 1344 1345 1346 1357 1358 1360 1361 1362 1373 1374 1376 1377 1378 1389 1390 1392 1393 1394 1405 1406 1408 1409 1410 1421 1422 1424 1425 1426 1437 1438 1440 1441 1442 1453 1454 1456 1457 1458 1469 1470 1472 1473 1474 1485 1486 1488 1489 1490 1501 1502 1504 1505 1506 1517 1518 1520 1521 1522 1533 1534 1536 1537 1538 1549 1550 1552 1553 1554 1565 1566 1568 1569 1570 1581 1582 1584 1585 1586 1597 1598 1600 1601 1602 1613 1614 1616 1617 1618 1629 1630 1632 1633 1634 1645 1646 1648 1649 1650 1661 1662 1664 1665 1666 1677 1678 1680 1681 1682 1693 1694 1696 1697 1698 1709 1710 1712 1713 1714 1725 1726 1728 1729 1730 1741 1742 1744 1745 1746 1757 1758 1760 1761 1762 1773 1774 1776 1777 1778 1789 1790 1792 1793 1794 1805 1806 1808 1809 1810 1821 1822 1824 1825 1826 1837 1838 1840 1841 1842 1853 1854 1856 1857 1858 1869 1870 1872 1873 1874 1885 1886 1888 1889 1890 1901 1902 1904 1905 1906 1917 1918 1920 1921 1922 1933 1934 1936 1937 1938 1949 1950 1952 1953 1954 1965 1966 1968 1969 1970 1981 1982 1984 1985 1986 1997 1998 2000 2001 2002 2013 2014 2016 2017 2018 2029 2030 2032 2033 2034 2045 2046" *)
  wire [2047:0] cur_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:25" *)
  input [1023:0] dat_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:26" *)
  input [63:0] dat_actv_nan;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:33" *)
  wire [127:0] nan_flag_l0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:34" *)
  wire [63:0] nan_flag_l1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:35" *)
  wire [31:0] nan_flag_l2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:36" *)
  wire [15:0] nan_flag_l3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:37" *)
  wire [7:0] nan_flag_l4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:38" *)
  wire [3:0] nan_flag_l5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:39" *)
  wire [1:0] nan_flag_l6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:40" *)
  wire nan_flag_l7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:41" *)
  wire [10:0] nan_mts_l0n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:42" *)
  wire [10:0] nan_mts_l0n1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:43" *)
  wire [10:0] nan_mts_l0n10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:44" *)
  wire [10:0] nan_mts_l0n100;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:45" *)
  wire [10:0] nan_mts_l0n101;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:46" *)
  wire [10:0] nan_mts_l0n102;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:47" *)
  wire [10:0] nan_mts_l0n103;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:48" *)
  wire [10:0] nan_mts_l0n104;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:49" *)
  wire [10:0] nan_mts_l0n105;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:50" *)
  wire [10:0] nan_mts_l0n106;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:51" *)
  wire [10:0] nan_mts_l0n107;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:52" *)
  wire [10:0] nan_mts_l0n108;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:53" *)
  wire [10:0] nan_mts_l0n109;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:54" *)
  wire [10:0] nan_mts_l0n11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:55" *)
  wire [10:0] nan_mts_l0n110;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:56" *)
  wire [10:0] nan_mts_l0n111;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:57" *)
  wire [10:0] nan_mts_l0n112;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:58" *)
  wire [10:0] nan_mts_l0n113;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:59" *)
  wire [10:0] nan_mts_l0n114;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:60" *)
  wire [10:0] nan_mts_l0n115;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:61" *)
  wire [10:0] nan_mts_l0n116;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:62" *)
  wire [10:0] nan_mts_l0n117;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:63" *)
  wire [10:0] nan_mts_l0n118;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:64" *)
  wire [10:0] nan_mts_l0n119;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:65" *)
  wire [10:0] nan_mts_l0n12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:66" *)
  wire [10:0] nan_mts_l0n120;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:67" *)
  wire [10:0] nan_mts_l0n121;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:68" *)
  wire [10:0] nan_mts_l0n122;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:69" *)
  wire [10:0] nan_mts_l0n123;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:70" *)
  wire [10:0] nan_mts_l0n124;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:71" *)
  wire [10:0] nan_mts_l0n125;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:72" *)
  wire [10:0] nan_mts_l0n126;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:73" *)
  wire [10:0] nan_mts_l0n127;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:74" *)
  wire [10:0] nan_mts_l0n13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:75" *)
  wire [10:0] nan_mts_l0n14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:76" *)
  wire [10:0] nan_mts_l0n15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:77" *)
  wire [10:0] nan_mts_l0n16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:78" *)
  wire [10:0] nan_mts_l0n17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:79" *)
  wire [10:0] nan_mts_l0n18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:80" *)
  wire [10:0] nan_mts_l0n19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:81" *)
  wire [10:0] nan_mts_l0n2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:82" *)
  wire [10:0] nan_mts_l0n20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:83" *)
  wire [10:0] nan_mts_l0n21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:84" *)
  wire [10:0] nan_mts_l0n22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:85" *)
  wire [10:0] nan_mts_l0n23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:86" *)
  wire [10:0] nan_mts_l0n24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:87" *)
  wire [10:0] nan_mts_l0n25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:88" *)
  wire [10:0] nan_mts_l0n26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:89" *)
  wire [10:0] nan_mts_l0n27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:90" *)
  wire [10:0] nan_mts_l0n28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:91" *)
  wire [10:0] nan_mts_l0n29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:92" *)
  wire [10:0] nan_mts_l0n3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:93" *)
  wire [10:0] nan_mts_l0n30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:94" *)
  wire [10:0] nan_mts_l0n31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:95" *)
  wire [10:0] nan_mts_l0n32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:96" *)
  wire [10:0] nan_mts_l0n33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:97" *)
  wire [10:0] nan_mts_l0n34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:98" *)
  wire [10:0] nan_mts_l0n35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:99" *)
  wire [10:0] nan_mts_l0n36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:100" *)
  wire [10:0] nan_mts_l0n37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:101" *)
  wire [10:0] nan_mts_l0n38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:102" *)
  wire [10:0] nan_mts_l0n39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:103" *)
  wire [10:0] nan_mts_l0n4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:104" *)
  wire [10:0] nan_mts_l0n40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:105" *)
  wire [10:0] nan_mts_l0n41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:106" *)
  wire [10:0] nan_mts_l0n42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:107" *)
  wire [10:0] nan_mts_l0n43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:108" *)
  wire [10:0] nan_mts_l0n44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:109" *)
  wire [10:0] nan_mts_l0n45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:110" *)
  wire [10:0] nan_mts_l0n46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:111" *)
  wire [10:0] nan_mts_l0n47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:112" *)
  wire [10:0] nan_mts_l0n48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:113" *)
  wire [10:0] nan_mts_l0n49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:114" *)
  wire [10:0] nan_mts_l0n5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:115" *)
  wire [10:0] nan_mts_l0n50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:116" *)
  wire [10:0] nan_mts_l0n51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:117" *)
  wire [10:0] nan_mts_l0n52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:118" *)
  wire [10:0] nan_mts_l0n53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:119" *)
  wire [10:0] nan_mts_l0n54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:120" *)
  wire [10:0] nan_mts_l0n55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:121" *)
  wire [10:0] nan_mts_l0n56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:122" *)
  wire [10:0] nan_mts_l0n57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:123" *)
  wire [10:0] nan_mts_l0n58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:124" *)
  wire [10:0] nan_mts_l0n59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:125" *)
  wire [10:0] nan_mts_l0n6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:126" *)
  wire [10:0] nan_mts_l0n60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:127" *)
  wire [10:0] nan_mts_l0n61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:128" *)
  wire [10:0] nan_mts_l0n62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:129" *)
  wire [10:0] nan_mts_l0n63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:130" *)
  wire [10:0] nan_mts_l0n64;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:131" *)
  wire [10:0] nan_mts_l0n65;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:132" *)
  wire [10:0] nan_mts_l0n66;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:133" *)
  wire [10:0] nan_mts_l0n67;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:134" *)
  wire [10:0] nan_mts_l0n68;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:135" *)
  wire [10:0] nan_mts_l0n69;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:136" *)
  wire [10:0] nan_mts_l0n7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:137" *)
  wire [10:0] nan_mts_l0n70;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:138" *)
  wire [10:0] nan_mts_l0n71;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:139" *)
  wire [10:0] nan_mts_l0n72;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:140" *)
  wire [10:0] nan_mts_l0n73;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:141" *)
  wire [10:0] nan_mts_l0n74;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:142" *)
  wire [10:0] nan_mts_l0n75;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:143" *)
  wire [10:0] nan_mts_l0n76;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:144" *)
  wire [10:0] nan_mts_l0n77;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:145" *)
  wire [10:0] nan_mts_l0n78;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:146" *)
  wire [10:0] nan_mts_l0n79;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:147" *)
  wire [10:0] nan_mts_l0n8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:148" *)
  wire [10:0] nan_mts_l0n80;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:149" *)
  wire [10:0] nan_mts_l0n81;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:150" *)
  wire [10:0] nan_mts_l0n82;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:151" *)
  wire [10:0] nan_mts_l0n83;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:152" *)
  wire [10:0] nan_mts_l0n84;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:153" *)
  wire [10:0] nan_mts_l0n85;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:154" *)
  wire [10:0] nan_mts_l0n86;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:155" *)
  wire [10:0] nan_mts_l0n87;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:156" *)
  wire [10:0] nan_mts_l0n88;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:157" *)
  wire [10:0] nan_mts_l0n89;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:158" *)
  wire [10:0] nan_mts_l0n9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:159" *)
  wire [10:0] nan_mts_l0n90;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:160" *)
  wire [10:0] nan_mts_l0n91;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:161" *)
  wire [10:0] nan_mts_l0n92;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:162" *)
  wire [10:0] nan_mts_l0n93;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:163" *)
  wire [10:0] nan_mts_l0n94;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:164" *)
  wire [10:0] nan_mts_l0n95;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:165" *)
  wire [10:0] nan_mts_l0n96;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:166" *)
  wire [10:0] nan_mts_l0n97;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:167" *)
  wire [10:0] nan_mts_l0n98;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:168" *)
  wire [10:0] nan_mts_l0n99;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:169" *)
  wire [10:0] nan_mts_l1n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:170" *)
  wire [10:0] nan_mts_l1n1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:171" *)
  wire [10:0] nan_mts_l1n10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:172" *)
  wire [10:0] nan_mts_l1n11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:173" *)
  wire [10:0] nan_mts_l1n12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:174" *)
  wire [10:0] nan_mts_l1n13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:175" *)
  wire [10:0] nan_mts_l1n14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:176" *)
  wire [10:0] nan_mts_l1n15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:177" *)
  wire [10:0] nan_mts_l1n16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:178" *)
  wire [10:0] nan_mts_l1n17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:179" *)
  wire [10:0] nan_mts_l1n18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:180" *)
  wire [10:0] nan_mts_l1n19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:181" *)
  wire [10:0] nan_mts_l1n2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:182" *)
  wire [10:0] nan_mts_l1n20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:183" *)
  wire [10:0] nan_mts_l1n21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:184" *)
  wire [10:0] nan_mts_l1n22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:185" *)
  wire [10:0] nan_mts_l1n23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:186" *)
  wire [10:0] nan_mts_l1n24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:187" *)
  wire [10:0] nan_mts_l1n25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:188" *)
  wire [10:0] nan_mts_l1n26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:189" *)
  wire [10:0] nan_mts_l1n27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:190" *)
  wire [10:0] nan_mts_l1n28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:191" *)
  wire [10:0] nan_mts_l1n29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:192" *)
  wire [10:0] nan_mts_l1n3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:193" *)
  wire [10:0] nan_mts_l1n30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:194" *)
  wire [10:0] nan_mts_l1n31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:195" *)
  wire [10:0] nan_mts_l1n32;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:196" *)
  wire [10:0] nan_mts_l1n33;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:197" *)
  wire [10:0] nan_mts_l1n34;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:198" *)
  wire [10:0] nan_mts_l1n35;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:199" *)
  wire [10:0] nan_mts_l1n36;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:200" *)
  wire [10:0] nan_mts_l1n37;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:201" *)
  wire [10:0] nan_mts_l1n38;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:202" *)
  wire [10:0] nan_mts_l1n39;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:203" *)
  wire [10:0] nan_mts_l1n4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:204" *)
  wire [10:0] nan_mts_l1n40;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:205" *)
  wire [10:0] nan_mts_l1n41;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:206" *)
  wire [10:0] nan_mts_l1n42;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:207" *)
  wire [10:0] nan_mts_l1n43;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:208" *)
  wire [10:0] nan_mts_l1n44;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:209" *)
  wire [10:0] nan_mts_l1n45;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:210" *)
  wire [10:0] nan_mts_l1n46;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:211" *)
  wire [10:0] nan_mts_l1n47;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:212" *)
  wire [10:0] nan_mts_l1n48;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:213" *)
  wire [10:0] nan_mts_l1n49;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:214" *)
  wire [10:0] nan_mts_l1n5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:215" *)
  wire [10:0] nan_mts_l1n50;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:216" *)
  wire [10:0] nan_mts_l1n51;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:217" *)
  wire [10:0] nan_mts_l1n52;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:218" *)
  wire [10:0] nan_mts_l1n53;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:219" *)
  wire [10:0] nan_mts_l1n54;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:220" *)
  wire [10:0] nan_mts_l1n55;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:221" *)
  wire [10:0] nan_mts_l1n56;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:222" *)
  wire [10:0] nan_mts_l1n57;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:223" *)
  wire [10:0] nan_mts_l1n58;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:224" *)
  wire [10:0] nan_mts_l1n59;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:225" *)
  wire [10:0] nan_mts_l1n6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:226" *)
  wire [10:0] nan_mts_l1n60;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:227" *)
  wire [10:0] nan_mts_l1n61;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:228" *)
  wire [10:0] nan_mts_l1n62;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:229" *)
  wire [10:0] nan_mts_l1n63;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:230" *)
  wire [10:0] nan_mts_l1n7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:231" *)
  wire [10:0] nan_mts_l1n8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:232" *)
  wire [10:0] nan_mts_l1n9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:233" *)
  wire [10:0] nan_mts_l2n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:234" *)
  wire [10:0] nan_mts_l2n1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:235" *)
  wire [10:0] nan_mts_l2n10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:236" *)
  wire [10:0] nan_mts_l2n11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:237" *)
  wire [10:0] nan_mts_l2n12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:238" *)
  wire [10:0] nan_mts_l2n13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:239" *)
  wire [10:0] nan_mts_l2n14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:240" *)
  wire [10:0] nan_mts_l2n15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:241" *)
  wire [10:0] nan_mts_l2n16;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:242" *)
  wire [10:0] nan_mts_l2n17;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:243" *)
  wire [10:0] nan_mts_l2n18;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:244" *)
  wire [10:0] nan_mts_l2n19;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:245" *)
  wire [10:0] nan_mts_l2n2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:246" *)
  wire [10:0] nan_mts_l2n20;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:247" *)
  wire [10:0] nan_mts_l2n21;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:248" *)
  wire [10:0] nan_mts_l2n22;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:249" *)
  wire [10:0] nan_mts_l2n23;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:250" *)
  wire [10:0] nan_mts_l2n24;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:251" *)
  wire [10:0] nan_mts_l2n25;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:252" *)
  wire [10:0] nan_mts_l2n26;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:253" *)
  wire [10:0] nan_mts_l2n27;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:254" *)
  wire [10:0] nan_mts_l2n28;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:255" *)
  wire [10:0] nan_mts_l2n29;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:256" *)
  wire [10:0] nan_mts_l2n3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:257" *)
  wire [10:0] nan_mts_l2n30;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:258" *)
  wire [10:0] nan_mts_l2n31;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:259" *)
  wire [10:0] nan_mts_l2n4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:260" *)
  wire [10:0] nan_mts_l2n5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:261" *)
  wire [10:0] nan_mts_l2n6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:262" *)
  wire [10:0] nan_mts_l2n7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:263" *)
  wire [10:0] nan_mts_l2n8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:264" *)
  wire [10:0] nan_mts_l2n9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:265" *)
  wire [10:0] nan_mts_l3n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:266" *)
  wire [10:0] nan_mts_l3n1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:267" *)
  wire [10:0] nan_mts_l3n10;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:268" *)
  wire [10:0] nan_mts_l3n11;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:269" *)
  wire [10:0] nan_mts_l3n12;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:270" *)
  wire [10:0] nan_mts_l3n13;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:271" *)
  wire [10:0] nan_mts_l3n14;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:272" *)
  wire [10:0] nan_mts_l3n15;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:273" *)
  wire [10:0] nan_mts_l3n2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:274" *)
  wire [10:0] nan_mts_l3n3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:275" *)
  wire [10:0] nan_mts_l3n4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:276" *)
  wire [10:0] nan_mts_l3n5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:277" *)
  wire [10:0] nan_mts_l3n6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:278" *)
  wire [10:0] nan_mts_l3n7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:279" *)
  wire [10:0] nan_mts_l3n8;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:280" *)
  wire [10:0] nan_mts_l3n9;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:281" *)
  wire [10:0] nan_mts_l4n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:282" *)
  wire [10:0] nan_mts_l4n1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:283" *)
  wire [10:0] nan_mts_l4n2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:284" *)
  wire [10:0] nan_mts_l4n3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:285" *)
  wire [10:0] nan_mts_l4n4;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:286" *)
  wire [10:0] nan_mts_l4n5;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:287" *)
  wire [10:0] nan_mts_l4n6;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:288" *)
  wire [10:0] nan_mts_l4n7;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:289" *)
  wire [10:0] nan_mts_l5n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:290" *)
  wire [10:0] nan_mts_l5n1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:291" *)
  wire [10:0] nan_mts_l5n2;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:292" *)
  wire [10:0] nan_mts_l5n3;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:293" *)
  wire [10:0] nan_mts_l6n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:294" *)
  wire [10:0] nan_mts_l6n1;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:295" *)
  wire [10:0] nan_mts_l7n0;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:21" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:22" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:29" *)
  output [10:0] out_nan_mts;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:30" *)
  output out_nan_pvld;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:27" *)
  input [1023:0] wt_actv_data;
  (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:28" *)
  input [63:0] wt_actv_nan;
  assign out_nan_pvld = cfg_is_fp16_d1[32] & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1086" *) _001_;
  assign out_nan_mts = nan_mts_l7n0 & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1088" *) { nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7, nan_flag_l7 };
  assign nan_flag_l0 = { cfg_is_fp16_d1[31:0], cfg_is_fp16_d1[31:0], cfg_is_fp16_d1[31:0], cfg_is_fp16_d1[31:0] } & (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:377" *) { dat_actv_nan, wt_actv_nan };
  assign nan_flag_l4[0] = nan_flag_l3[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1020" *) nan_flag_l3[1];
  assign nan_flag_l4[1] = nan_flag_l3[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1021" *) nan_flag_l3[3];
  assign nan_flag_l4[2] = nan_flag_l3[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1022" *) nan_flag_l3[5];
  assign nan_flag_l4[3] = nan_flag_l3[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1023" *) nan_flag_l3[7];
  assign nan_flag_l4[4] = nan_flag_l3[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1024" *) nan_flag_l3[9];
  assign nan_flag_l4[5] = nan_flag_l3[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1025" *) nan_flag_l3[11];
  assign nan_flag_l4[6] = nan_flag_l3[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1026" *) nan_flag_l3[13];
  assign nan_flag_l4[7] = nan_flag_l3[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1027" *) nan_flag_l3[15];
  assign nan_flag_l5[0] = nan_flag_l4[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1048" *) nan_flag_l4[1];
  assign nan_flag_l5[1] = nan_flag_l4[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1049" *) nan_flag_l4[3];
  assign nan_flag_l5[2] = nan_flag_l4[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1050" *) nan_flag_l4[5];
  assign nan_flag_l5[3] = nan_flag_l4[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1051" *) nan_flag_l4[7];
  assign nan_flag_l6[0] = nan_flag_l5[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1066" *) nan_flag_l5[1];
  assign nan_flag_l6[1] = nan_flag_l5[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1067" *) nan_flag_l5[3];
  assign nan_flag_l7 = nan_flag_l6[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1079" *) nan_flag_l6[1];
  assign nan_flag_l1[0] = nan_flag_l0[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:716" *) nan_flag_l0[1];
  assign nan_flag_l1[1] = nan_flag_l0[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:717" *) nan_flag_l0[3];
  assign nan_flag_l1[2] = nan_flag_l0[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:718" *) nan_flag_l0[5];
  assign nan_flag_l1[3] = nan_flag_l0[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:719" *) nan_flag_l0[7];
  assign nan_flag_l1[4] = nan_flag_l0[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:720" *) nan_flag_l0[9];
  assign nan_flag_l1[5] = nan_flag_l0[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:721" *) nan_flag_l0[11];
  assign nan_flag_l1[6] = nan_flag_l0[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:722" *) nan_flag_l0[13];
  assign nan_flag_l1[7] = nan_flag_l0[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:723" *) nan_flag_l0[15];
  assign nan_flag_l1[8] = nan_flag_l0[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:724" *) nan_flag_l0[17];
  assign nan_flag_l1[9] = nan_flag_l0[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:725" *) nan_flag_l0[19];
  assign nan_flag_l1[10] = nan_flag_l0[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:726" *) nan_flag_l0[21];
  assign nan_flag_l1[11] = nan_flag_l0[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:727" *) nan_flag_l0[23];
  assign nan_flag_l1[12] = nan_flag_l0[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:728" *) nan_flag_l0[25];
  assign nan_flag_l1[13] = nan_flag_l0[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:729" *) nan_flag_l0[27];
  assign nan_flag_l1[14] = nan_flag_l0[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:730" *) nan_flag_l0[29];
  assign nan_flag_l1[15] = nan_flag_l0[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:731" *) nan_flag_l0[31];
  assign nan_flag_l1[16] = nan_flag_l0[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:732" *) nan_flag_l0[33];
  assign nan_flag_l1[17] = nan_flag_l0[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:733" *) nan_flag_l0[35];
  assign nan_flag_l1[18] = nan_flag_l0[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:734" *) nan_flag_l0[37];
  assign nan_flag_l1[19] = nan_flag_l0[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:735" *) nan_flag_l0[39];
  assign nan_flag_l1[20] = nan_flag_l0[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:736" *) nan_flag_l0[41];
  assign nan_flag_l1[21] = nan_flag_l0[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:737" *) nan_flag_l0[43];
  assign nan_flag_l1[22] = nan_flag_l0[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:738" *) nan_flag_l0[45];
  assign nan_flag_l1[23] = nan_flag_l0[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:739" *) nan_flag_l0[47];
  assign nan_flag_l1[24] = nan_flag_l0[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:740" *) nan_flag_l0[49];
  assign nan_flag_l1[25] = nan_flag_l0[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:741" *) nan_flag_l0[51];
  assign nan_flag_l1[26] = nan_flag_l0[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:742" *) nan_flag_l0[53];
  assign nan_flag_l1[27] = nan_flag_l0[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:743" *) nan_flag_l0[55];
  assign nan_flag_l1[28] = nan_flag_l0[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:744" *) nan_flag_l0[57];
  assign nan_flag_l1[29] = nan_flag_l0[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:745" *) nan_flag_l0[59];
  assign nan_flag_l1[30] = nan_flag_l0[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:746" *) nan_flag_l0[61];
  assign nan_flag_l1[31] = nan_flag_l0[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:747" *) nan_flag_l0[63];
  assign nan_flag_l1[32] = nan_flag_l0[64] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:748" *) nan_flag_l0[65];
  assign nan_flag_l1[33] = nan_flag_l0[66] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:749" *) nan_flag_l0[67];
  assign nan_flag_l1[34] = nan_flag_l0[68] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:750" *) nan_flag_l0[69];
  assign nan_flag_l1[35] = nan_flag_l0[70] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:751" *) nan_flag_l0[71];
  assign nan_flag_l1[36] = nan_flag_l0[72] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:752" *) nan_flag_l0[73];
  assign nan_flag_l1[37] = nan_flag_l0[74] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:753" *) nan_flag_l0[75];
  assign nan_flag_l1[38] = nan_flag_l0[76] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:754" *) nan_flag_l0[77];
  assign nan_flag_l1[39] = nan_flag_l0[78] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:755" *) nan_flag_l0[79];
  assign nan_flag_l1[40] = nan_flag_l0[80] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:756" *) nan_flag_l0[81];
  assign nan_flag_l1[41] = nan_flag_l0[82] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:757" *) nan_flag_l0[83];
  assign nan_flag_l1[42] = nan_flag_l0[84] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:758" *) nan_flag_l0[85];
  assign nan_flag_l1[43] = nan_flag_l0[86] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:759" *) nan_flag_l0[87];
  assign nan_flag_l1[44] = nan_flag_l0[88] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:760" *) nan_flag_l0[89];
  assign nan_flag_l1[45] = nan_flag_l0[90] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:761" *) nan_flag_l0[91];
  assign nan_flag_l1[46] = nan_flag_l0[92] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:762" *) nan_flag_l0[93];
  assign nan_flag_l1[47] = nan_flag_l0[94] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:763" *) nan_flag_l0[95];
  assign nan_flag_l1[48] = nan_flag_l0[96] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:764" *) nan_flag_l0[97];
  assign nan_flag_l1[49] = nan_flag_l0[98] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:765" *) nan_flag_l0[99];
  assign nan_flag_l1[50] = nan_flag_l0[100] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:766" *) nan_flag_l0[101];
  assign nan_flag_l1[51] = nan_flag_l0[102] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:767" *) nan_flag_l0[103];
  assign nan_flag_l1[52] = nan_flag_l0[104] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:768" *) nan_flag_l0[105];
  assign nan_flag_l1[53] = nan_flag_l0[106] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:769" *) nan_flag_l0[107];
  assign nan_flag_l1[54] = nan_flag_l0[108] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:770" *) nan_flag_l0[109];
  assign nan_flag_l1[55] = nan_flag_l0[110] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:771" *) nan_flag_l0[111];
  assign nan_flag_l1[56] = nan_flag_l0[112] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:772" *) nan_flag_l0[113];
  assign nan_flag_l1[57] = nan_flag_l0[114] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:773" *) nan_flag_l0[115];
  assign nan_flag_l1[58] = nan_flag_l0[116] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:774" *) nan_flag_l0[117];
  assign nan_flag_l1[59] = nan_flag_l0[118] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:775" *) nan_flag_l0[119];
  assign nan_flag_l1[60] = nan_flag_l0[120] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:776" *) nan_flag_l0[121];
  assign nan_flag_l1[61] = nan_flag_l0[122] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:777" *) nan_flag_l0[123];
  assign nan_flag_l1[62] = nan_flag_l0[124] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:778" *) nan_flag_l0[125];
  assign nan_flag_l1[63] = nan_flag_l0[126] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:779" *) nan_flag_l0[127];
  assign nan_flag_l2[0] = nan_flag_l1[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:884" *) nan_flag_l1[1];
  assign nan_flag_l2[1] = nan_flag_l1[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:885" *) nan_flag_l1[3];
  assign nan_flag_l2[2] = nan_flag_l1[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:886" *) nan_flag_l1[5];
  assign nan_flag_l2[3] = nan_flag_l1[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:887" *) nan_flag_l1[7];
  assign nan_flag_l2[4] = nan_flag_l1[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:888" *) nan_flag_l1[9];
  assign nan_flag_l2[5] = nan_flag_l1[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:889" *) nan_flag_l1[11];
  assign nan_flag_l2[6] = nan_flag_l1[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:890" *) nan_flag_l1[13];
  assign nan_flag_l2[7] = nan_flag_l1[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:891" *) nan_flag_l1[15];
  assign nan_flag_l2[8] = nan_flag_l1[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:892" *) nan_flag_l1[17];
  assign nan_flag_l2[9] = nan_flag_l1[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:893" *) nan_flag_l1[19];
  assign nan_flag_l2[10] = nan_flag_l1[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:894" *) nan_flag_l1[21];
  assign nan_flag_l2[11] = nan_flag_l1[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:895" *) nan_flag_l1[23];
  assign nan_flag_l2[12] = nan_flag_l1[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:896" *) nan_flag_l1[25];
  assign nan_flag_l2[13] = nan_flag_l1[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:897" *) nan_flag_l1[27];
  assign nan_flag_l2[14] = nan_flag_l1[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:898" *) nan_flag_l1[29];
  assign nan_flag_l2[15] = nan_flag_l1[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:899" *) nan_flag_l1[31];
  assign nan_flag_l2[16] = nan_flag_l1[32] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:900" *) nan_flag_l1[33];
  assign nan_flag_l2[17] = nan_flag_l1[34] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:901" *) nan_flag_l1[35];
  assign nan_flag_l2[18] = nan_flag_l1[36] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:902" *) nan_flag_l1[37];
  assign nan_flag_l2[19] = nan_flag_l1[38] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:903" *) nan_flag_l1[39];
  assign nan_flag_l2[20] = nan_flag_l1[40] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:904" *) nan_flag_l1[41];
  assign nan_flag_l2[21] = nan_flag_l1[42] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:905" *) nan_flag_l1[43];
  assign nan_flag_l2[22] = nan_flag_l1[44] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:906" *) nan_flag_l1[45];
  assign nan_flag_l2[23] = nan_flag_l1[46] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:907" *) nan_flag_l1[47];
  assign nan_flag_l2[24] = nan_flag_l1[48] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:908" *) nan_flag_l1[49];
  assign nan_flag_l2[25] = nan_flag_l1[50] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:909" *) nan_flag_l1[51];
  assign nan_flag_l2[26] = nan_flag_l1[52] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:910" *) nan_flag_l1[53];
  assign nan_flag_l2[27] = nan_flag_l1[54] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:911" *) nan_flag_l1[55];
  assign nan_flag_l2[28] = nan_flag_l1[56] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:912" *) nan_flag_l1[57];
  assign nan_flag_l2[29] = nan_flag_l1[58] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:913" *) nan_flag_l1[59];
  assign nan_flag_l2[30] = nan_flag_l1[60] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:914" *) nan_flag_l1[61];
  assign nan_flag_l2[31] = nan_flag_l1[62] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:915" *) nan_flag_l1[63];
  assign nan_flag_l3[0] = nan_flag_l2[0] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:972" *) nan_flag_l2[1];
  assign nan_flag_l3[1] = nan_flag_l2[2] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:973" *) nan_flag_l2[3];
  assign nan_flag_l3[2] = nan_flag_l2[4] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:974" *) nan_flag_l2[5];
  assign nan_flag_l3[3] = nan_flag_l2[6] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:975" *) nan_flag_l2[7];
  assign nan_flag_l3[4] = nan_flag_l2[8] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:976" *) nan_flag_l2[9];
  assign nan_flag_l3[5] = nan_flag_l2[10] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:977" *) nan_flag_l2[11];
  assign nan_flag_l3[6] = nan_flag_l2[12] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:978" *) nan_flag_l2[13];
  assign nan_flag_l3[7] = nan_flag_l2[14] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:979" *) nan_flag_l2[15];
  assign nan_flag_l3[8] = nan_flag_l2[16] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:980" *) nan_flag_l2[17];
  assign nan_flag_l3[9] = nan_flag_l2[18] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:981" *) nan_flag_l2[19];
  assign nan_flag_l3[10] = nan_flag_l2[20] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:982" *) nan_flag_l2[21];
  assign nan_flag_l3[11] = nan_flag_l2[22] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:983" *) nan_flag_l2[23];
  assign nan_flag_l3[12] = nan_flag_l2[24] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:984" *) nan_flag_l2[25];
  assign nan_flag_l3[13] = nan_flag_l2[26] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:985" *) nan_flag_l2[27];
  assign nan_flag_l3[14] = nan_flag_l2[28] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:986" *) nan_flag_l2[29];
  assign nan_flag_l3[15] = nan_flag_l2[30] | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:987" *) nan_flag_l2[31];
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_is_fp16_d1 <= 33'b000000000000000000000000000000000;
    else
      cfg_is_fp16_d1 <= _000_;
  assign _000_ = cfg_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:312" *) { cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16, cfg_is_fp16 } : cfg_is_fp16_d1;
  assign _001_ = | (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1086" *) { dat_actv_nan[0], dat_actv_nan[1], dat_actv_nan[2], dat_actv_nan[3], dat_actv_nan[4], dat_actv_nan[5], dat_actv_nan[6], dat_actv_nan[7], dat_actv_nan[8], dat_actv_nan[9], dat_actv_nan[10], dat_actv_nan[11], dat_actv_nan[12], dat_actv_nan[13], dat_actv_nan[14], dat_actv_nan[15], dat_actv_nan[16], dat_actv_nan[17], dat_actv_nan[18], dat_actv_nan[19], dat_actv_nan[20], dat_actv_nan[21], dat_actv_nan[22], dat_actv_nan[23], dat_actv_nan[24], dat_actv_nan[25], dat_actv_nan[26], dat_actv_nan[27], dat_actv_nan[28], dat_actv_nan[29], dat_actv_nan[30], dat_actv_nan[31], dat_actv_nan[32], dat_actv_nan[33], dat_actv_nan[34], dat_actv_nan[35], dat_actv_nan[36], dat_actv_nan[37], dat_actv_nan[38], dat_actv_nan[39], dat_actv_nan[40], dat_actv_nan[41], dat_actv_nan[42], dat_actv_nan[43], dat_actv_nan[44], dat_actv_nan[45], dat_actv_nan[46], dat_actv_nan[47], dat_actv_nan[48], dat_actv_nan[49], dat_actv_nan[50], dat_actv_nan[51], dat_actv_nan[52], dat_actv_nan[53], dat_actv_nan[54], dat_actv_nan[55], dat_actv_nan[56], dat_actv_nan[57], dat_actv_nan[58], dat_actv_nan[59], dat_actv_nan[60], dat_actv_nan[61], dat_actv_nan[62], dat_actv_nan[63], wt_actv_nan[0], wt_actv_nan[1], wt_actv_nan[2], wt_actv_nan[3], wt_actv_nan[4], wt_actv_nan[5], wt_actv_nan[6], wt_actv_nan[7], wt_actv_nan[8], wt_actv_nan[9], wt_actv_nan[10], wt_actv_nan[11], wt_actv_nan[12], wt_actv_nan[13], wt_actv_nan[14], wt_actv_nan[15], wt_actv_nan[16], wt_actv_nan[17], wt_actv_nan[18], wt_actv_nan[19], wt_actv_nan[20], wt_actv_nan[21], wt_actv_nan[22], wt_actv_nan[23], wt_actv_nan[24], wt_actv_nan[25], wt_actv_nan[26], wt_actv_nan[27], wt_actv_nan[28], wt_actv_nan[29], wt_actv_nan[30], wt_actv_nan[31], wt_actv_nan[32], wt_actv_nan[33], wt_actv_nan[34], wt_actv_nan[35], wt_actv_nan[36], wt_actv_nan[37], wt_actv_nan[38], wt_actv_nan[39], wt_actv_nan[40], wt_actv_nan[41], wt_actv_nan[42], wt_actv_nan[43], wt_actv_nan[44], wt_actv_nan[45], wt_actv_nan[46], wt_actv_nan[47], wt_actv_nan[48], wt_actv_nan[49], wt_actv_nan[50], wt_actv_nan[51], wt_actv_nan[52], wt_actv_nan[53], wt_actv_nan[54], wt_actv_nan[55], wt_actv_nan[56], wt_actv_nan[57], wt_actv_nan[58], wt_actv_nan[59], wt_actv_nan[60], wt_actv_nan[61], wt_actv_nan[62], wt_actv_nan[63] };
  assign nan_mts_l4n0 = nan_flag_l3[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1008" *) nan_mts_l3n0 : nan_mts_l3n1;
  assign nan_mts_l4n1 = nan_flag_l3[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1009" *) nan_mts_l3n2 : nan_mts_l3n3;
  assign nan_mts_l4n2 = nan_flag_l3[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1010" *) nan_mts_l3n4 : nan_mts_l3n5;
  assign nan_mts_l4n3 = nan_flag_l3[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1011" *) nan_mts_l3n6 : nan_mts_l3n7;
  assign nan_mts_l4n4 = nan_flag_l3[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1012" *) nan_mts_l3n8 : nan_mts_l3n9;
  assign nan_mts_l4n5 = nan_flag_l3[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1013" *) nan_mts_l3n10 : nan_mts_l3n11;
  assign nan_mts_l4n6 = nan_flag_l3[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1014" *) nan_mts_l3n12 : nan_mts_l3n13;
  assign nan_mts_l4n7 = nan_flag_l3[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1015" *) nan_mts_l3n14 : nan_mts_l3n15;
  assign nan_mts_l5n0 = nan_flag_l4[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1040" *) nan_mts_l4n0 : nan_mts_l4n1;
  assign nan_mts_l5n1 = nan_flag_l4[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1041" *) nan_mts_l4n2 : nan_mts_l4n3;
  assign nan_mts_l5n2 = nan_flag_l4[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1042" *) nan_mts_l4n4 : nan_mts_l4n5;
  assign nan_mts_l5n3 = nan_flag_l4[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1043" *) nan_mts_l4n6 : nan_mts_l4n7;
  assign nan_mts_l6n0 = nan_flag_l5[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1060" *) nan_mts_l5n0 : nan_mts_l5n1;
  assign nan_mts_l6n1 = nan_flag_l5[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1061" *) nan_mts_l5n2 : nan_mts_l5n3;
  assign nan_mts_l7n0 = nan_flag_l6[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:1074" *) nan_mts_l6n0 : nan_mts_l6n1;
  assign nan_mts_l1n0 = nan_flag_l0[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:648" *) { wt_actv_data[15], wt_actv_data[12:3] } : { wt_actv_data[31], wt_actv_data[28:19] };
  assign nan_mts_l1n1 = nan_flag_l0[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:649" *) { wt_actv_data[47], wt_actv_data[44:35] } : { wt_actv_data[63], wt_actv_data[60:51] };
  assign nan_mts_l1n2 = nan_flag_l0[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:650" *) { wt_actv_data[79], wt_actv_data[76:67] } : { wt_actv_data[95], wt_actv_data[92:83] };
  assign nan_mts_l1n3 = nan_flag_l0[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:651" *) { wt_actv_data[111], wt_actv_data[108:99] } : { wt_actv_data[127], wt_actv_data[124:115] };
  assign nan_mts_l1n4 = nan_flag_l0[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:652" *) { wt_actv_data[143], wt_actv_data[140:131] } : { wt_actv_data[159], wt_actv_data[156:147] };
  assign nan_mts_l1n5 = nan_flag_l0[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:653" *) { wt_actv_data[175], wt_actv_data[172:163] } : { wt_actv_data[191], wt_actv_data[188:179] };
  assign nan_mts_l1n6 = nan_flag_l0[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:654" *) { wt_actv_data[207], wt_actv_data[204:195] } : { wt_actv_data[223], wt_actv_data[220:211] };
  assign nan_mts_l1n7 = nan_flag_l0[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:655" *) { wt_actv_data[239], wt_actv_data[236:227] } : { wt_actv_data[255], wt_actv_data[252:243] };
  assign nan_mts_l1n8 = nan_flag_l0[16] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:656" *) { wt_actv_data[271], wt_actv_data[268:259] } : { wt_actv_data[287], wt_actv_data[284:275] };
  assign nan_mts_l1n9 = nan_flag_l0[18] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:657" *) { wt_actv_data[303], wt_actv_data[300:291] } : { wt_actv_data[319], wt_actv_data[316:307] };
  assign nan_mts_l1n10 = nan_flag_l0[20] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:658" *) { wt_actv_data[335], wt_actv_data[332:323] } : { wt_actv_data[351], wt_actv_data[348:339] };
  assign nan_mts_l1n11 = nan_flag_l0[22] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:659" *) { wt_actv_data[367], wt_actv_data[364:355] } : { wt_actv_data[383], wt_actv_data[380:371] };
  assign nan_mts_l1n12 = nan_flag_l0[24] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:660" *) { wt_actv_data[399], wt_actv_data[396:387] } : { wt_actv_data[415], wt_actv_data[412:403] };
  assign nan_mts_l1n13 = nan_flag_l0[26] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:661" *) { wt_actv_data[431], wt_actv_data[428:419] } : { wt_actv_data[447], wt_actv_data[444:435] };
  assign nan_mts_l1n14 = nan_flag_l0[28] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:662" *) { wt_actv_data[463], wt_actv_data[460:451] } : { wt_actv_data[479], wt_actv_data[476:467] };
  assign nan_mts_l1n15 = nan_flag_l0[30] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:663" *) { wt_actv_data[495], wt_actv_data[492:483] } : { wt_actv_data[511], wt_actv_data[508:499] };
  assign nan_mts_l1n16 = nan_flag_l0[32] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:664" *) { wt_actv_data[527], wt_actv_data[524:515] } : { wt_actv_data[543], wt_actv_data[540:531] };
  assign nan_mts_l1n17 = nan_flag_l0[34] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:665" *) { wt_actv_data[559], wt_actv_data[556:547] } : { wt_actv_data[575], wt_actv_data[572:563] };
  assign nan_mts_l1n18 = nan_flag_l0[36] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:666" *) { wt_actv_data[591], wt_actv_data[588:579] } : { wt_actv_data[607], wt_actv_data[604:595] };
  assign nan_mts_l1n19 = nan_flag_l0[38] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:667" *) { wt_actv_data[623], wt_actv_data[620:611] } : { wt_actv_data[639], wt_actv_data[636:627] };
  assign nan_mts_l1n20 = nan_flag_l0[40] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:668" *) { wt_actv_data[655], wt_actv_data[652:643] } : { wt_actv_data[671], wt_actv_data[668:659] };
  assign nan_mts_l1n21 = nan_flag_l0[42] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:669" *) { wt_actv_data[687], wt_actv_data[684:675] } : { wt_actv_data[703], wt_actv_data[700:691] };
  assign nan_mts_l1n22 = nan_flag_l0[44] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:670" *) { wt_actv_data[719], wt_actv_data[716:707] } : { wt_actv_data[735], wt_actv_data[732:723] };
  assign nan_mts_l1n23 = nan_flag_l0[46] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:671" *) { wt_actv_data[751], wt_actv_data[748:739] } : { wt_actv_data[767], wt_actv_data[764:755] };
  assign nan_mts_l1n24 = nan_flag_l0[48] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:672" *) { wt_actv_data[783], wt_actv_data[780:771] } : { wt_actv_data[799], wt_actv_data[796:787] };
  assign nan_mts_l1n25 = nan_flag_l0[50] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:673" *) { wt_actv_data[815], wt_actv_data[812:803] } : { wt_actv_data[831], wt_actv_data[828:819] };
  assign nan_mts_l1n26 = nan_flag_l0[52] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:674" *) { wt_actv_data[847], wt_actv_data[844:835] } : { wt_actv_data[863], wt_actv_data[860:851] };
  assign nan_mts_l1n27 = nan_flag_l0[54] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:675" *) { wt_actv_data[879], wt_actv_data[876:867] } : { wt_actv_data[895], wt_actv_data[892:883] };
  assign nan_mts_l1n28 = nan_flag_l0[56] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:676" *) { wt_actv_data[911], wt_actv_data[908:899] } : { wt_actv_data[927], wt_actv_data[924:915] };
  assign nan_mts_l1n29 = nan_flag_l0[58] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:677" *) { wt_actv_data[943], wt_actv_data[940:931] } : { wt_actv_data[959], wt_actv_data[956:947] };
  assign nan_mts_l1n30 = nan_flag_l0[60] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:678" *) { wt_actv_data[975], wt_actv_data[972:963] } : { wt_actv_data[991], wt_actv_data[988:979] };
  assign nan_mts_l1n31 = nan_flag_l0[62] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:679" *) { wt_actv_data[1007], wt_actv_data[1004:995] } : { wt_actv_data[1023], wt_actv_data[1020:1011] };
  assign nan_mts_l1n32 = nan_flag_l0[64] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:680" *) { dat_actv_data[15], dat_actv_data[12:3] } : { dat_actv_data[31], dat_actv_data[28:19] };
  assign nan_mts_l1n33 = nan_flag_l0[66] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:681" *) { dat_actv_data[47], dat_actv_data[44:35] } : { dat_actv_data[63], dat_actv_data[60:51] };
  assign nan_mts_l1n34 = nan_flag_l0[68] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:682" *) { dat_actv_data[79], dat_actv_data[76:67] } : { dat_actv_data[95], dat_actv_data[92:83] };
  assign nan_mts_l1n35 = nan_flag_l0[70] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:683" *) { dat_actv_data[111], dat_actv_data[108:99] } : { dat_actv_data[127], dat_actv_data[124:115] };
  assign nan_mts_l1n36 = nan_flag_l0[72] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:684" *) { dat_actv_data[143], dat_actv_data[140:131] } : { dat_actv_data[159], dat_actv_data[156:147] };
  assign nan_mts_l1n37 = nan_flag_l0[74] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:685" *) { dat_actv_data[175], dat_actv_data[172:163] } : { dat_actv_data[191], dat_actv_data[188:179] };
  assign nan_mts_l1n38 = nan_flag_l0[76] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:686" *) { dat_actv_data[207], dat_actv_data[204:195] } : { dat_actv_data[223], dat_actv_data[220:211] };
  assign nan_mts_l1n39 = nan_flag_l0[78] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:687" *) { dat_actv_data[239], dat_actv_data[236:227] } : { dat_actv_data[255], dat_actv_data[252:243] };
  assign nan_mts_l1n40 = nan_flag_l0[80] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:688" *) { dat_actv_data[271], dat_actv_data[268:259] } : { dat_actv_data[287], dat_actv_data[284:275] };
  assign nan_mts_l1n41 = nan_flag_l0[82] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:689" *) { dat_actv_data[303], dat_actv_data[300:291] } : { dat_actv_data[319], dat_actv_data[316:307] };
  assign nan_mts_l1n42 = nan_flag_l0[84] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:690" *) { dat_actv_data[335], dat_actv_data[332:323] } : { dat_actv_data[351], dat_actv_data[348:339] };
  assign nan_mts_l1n43 = nan_flag_l0[86] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:691" *) { dat_actv_data[367], dat_actv_data[364:355] } : { dat_actv_data[383], dat_actv_data[380:371] };
  assign nan_mts_l1n44 = nan_flag_l0[88] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:692" *) { dat_actv_data[399], dat_actv_data[396:387] } : { dat_actv_data[415], dat_actv_data[412:403] };
  assign nan_mts_l1n45 = nan_flag_l0[90] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:693" *) { dat_actv_data[431], dat_actv_data[428:419] } : { dat_actv_data[447], dat_actv_data[444:435] };
  assign nan_mts_l1n46 = nan_flag_l0[92] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:694" *) { dat_actv_data[463], dat_actv_data[460:451] } : { dat_actv_data[479], dat_actv_data[476:467] };
  assign nan_mts_l1n47 = nan_flag_l0[94] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:695" *) { dat_actv_data[495], dat_actv_data[492:483] } : { dat_actv_data[511], dat_actv_data[508:499] };
  assign nan_mts_l1n48 = nan_flag_l0[96] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:696" *) { dat_actv_data[527], dat_actv_data[524:515] } : { dat_actv_data[543], dat_actv_data[540:531] };
  assign nan_mts_l1n49 = nan_flag_l0[98] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:697" *) { dat_actv_data[559], dat_actv_data[556:547] } : { dat_actv_data[575], dat_actv_data[572:563] };
  assign nan_mts_l1n50 = nan_flag_l0[100] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:698" *) { dat_actv_data[591], dat_actv_data[588:579] } : { dat_actv_data[607], dat_actv_data[604:595] };
  assign nan_mts_l1n51 = nan_flag_l0[102] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:699" *) { dat_actv_data[623], dat_actv_data[620:611] } : { dat_actv_data[639], dat_actv_data[636:627] };
  assign nan_mts_l1n52 = nan_flag_l0[104] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:700" *) { dat_actv_data[655], dat_actv_data[652:643] } : { dat_actv_data[671], dat_actv_data[668:659] };
  assign nan_mts_l1n53 = nan_flag_l0[106] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:701" *) { dat_actv_data[687], dat_actv_data[684:675] } : { dat_actv_data[703], dat_actv_data[700:691] };
  assign nan_mts_l1n54 = nan_flag_l0[108] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:702" *) { dat_actv_data[719], dat_actv_data[716:707] } : { dat_actv_data[735], dat_actv_data[732:723] };
  assign nan_mts_l1n55 = nan_flag_l0[110] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:703" *) { dat_actv_data[751], dat_actv_data[748:739] } : { dat_actv_data[767], dat_actv_data[764:755] };
  assign nan_mts_l1n56 = nan_flag_l0[112] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:704" *) { dat_actv_data[783], dat_actv_data[780:771] } : { dat_actv_data[799], dat_actv_data[796:787] };
  assign nan_mts_l1n57 = nan_flag_l0[114] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:705" *) { dat_actv_data[815], dat_actv_data[812:803] } : { dat_actv_data[831], dat_actv_data[828:819] };
  assign nan_mts_l1n58 = nan_flag_l0[116] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:706" *) { dat_actv_data[847], dat_actv_data[844:835] } : { dat_actv_data[863], dat_actv_data[860:851] };
  assign nan_mts_l1n59 = nan_flag_l0[118] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:707" *) { dat_actv_data[879], dat_actv_data[876:867] } : { dat_actv_data[895], dat_actv_data[892:883] };
  assign nan_mts_l1n60 = nan_flag_l0[120] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:708" *) { dat_actv_data[911], dat_actv_data[908:899] } : { dat_actv_data[927], dat_actv_data[924:915] };
  assign nan_mts_l1n61 = nan_flag_l0[122] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:709" *) { dat_actv_data[943], dat_actv_data[940:931] } : { dat_actv_data[959], dat_actv_data[956:947] };
  assign nan_mts_l1n62 = nan_flag_l0[124] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:710" *) { dat_actv_data[975], dat_actv_data[972:963] } : { dat_actv_data[991], dat_actv_data[988:979] };
  assign nan_mts_l1n63 = nan_flag_l0[126] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:711" *) { dat_actv_data[1007], dat_actv_data[1004:995] } : { dat_actv_data[1023], dat_actv_data[1020:1011] };
  assign nan_mts_l2n0 = nan_flag_l1[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:848" *) nan_mts_l1n0 : nan_mts_l1n1;
  assign nan_mts_l2n1 = nan_flag_l1[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:849" *) nan_mts_l1n2 : nan_mts_l1n3;
  assign nan_mts_l2n2 = nan_flag_l1[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:850" *) nan_mts_l1n4 : nan_mts_l1n5;
  assign nan_mts_l2n3 = nan_flag_l1[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:851" *) nan_mts_l1n6 : nan_mts_l1n7;
  assign nan_mts_l2n4 = nan_flag_l1[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:852" *) nan_mts_l1n8 : nan_mts_l1n9;
  assign nan_mts_l2n5 = nan_flag_l1[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:853" *) nan_mts_l1n10 : nan_mts_l1n11;
  assign nan_mts_l2n6 = nan_flag_l1[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:854" *) nan_mts_l1n12 : nan_mts_l1n13;
  assign nan_mts_l2n7 = nan_flag_l1[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:855" *) nan_mts_l1n14 : nan_mts_l1n15;
  assign nan_mts_l2n8 = nan_flag_l1[16] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:856" *) nan_mts_l1n16 : nan_mts_l1n17;
  assign nan_mts_l2n9 = nan_flag_l1[18] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:857" *) nan_mts_l1n18 : nan_mts_l1n19;
  assign nan_mts_l2n10 = nan_flag_l1[20] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:858" *) nan_mts_l1n20 : nan_mts_l1n21;
  assign nan_mts_l2n11 = nan_flag_l1[22] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:859" *) nan_mts_l1n22 : nan_mts_l1n23;
  assign nan_mts_l2n12 = nan_flag_l1[24] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:860" *) nan_mts_l1n24 : nan_mts_l1n25;
  assign nan_mts_l2n13 = nan_flag_l1[26] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:861" *) nan_mts_l1n26 : nan_mts_l1n27;
  assign nan_mts_l2n14 = nan_flag_l1[28] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:862" *) nan_mts_l1n28 : nan_mts_l1n29;
  assign nan_mts_l2n15 = nan_flag_l1[30] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:863" *) nan_mts_l1n30 : nan_mts_l1n31;
  assign nan_mts_l2n16 = nan_flag_l1[32] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:864" *) nan_mts_l1n32 : nan_mts_l1n33;
  assign nan_mts_l2n17 = nan_flag_l1[34] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:865" *) nan_mts_l1n34 : nan_mts_l1n35;
  assign nan_mts_l2n18 = nan_flag_l1[36] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:866" *) nan_mts_l1n36 : nan_mts_l1n37;
  assign nan_mts_l2n19 = nan_flag_l1[38] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:867" *) nan_mts_l1n38 : nan_mts_l1n39;
  assign nan_mts_l2n20 = nan_flag_l1[40] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:868" *) nan_mts_l1n40 : nan_mts_l1n41;
  assign nan_mts_l2n21 = nan_flag_l1[42] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:869" *) nan_mts_l1n42 : nan_mts_l1n43;
  assign nan_mts_l2n22 = nan_flag_l1[44] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:870" *) nan_mts_l1n44 : nan_mts_l1n45;
  assign nan_mts_l2n23 = nan_flag_l1[46] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:871" *) nan_mts_l1n46 : nan_mts_l1n47;
  assign nan_mts_l2n24 = nan_flag_l1[48] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:872" *) nan_mts_l1n48 : nan_mts_l1n49;
  assign nan_mts_l2n25 = nan_flag_l1[50] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:873" *) nan_mts_l1n50 : nan_mts_l1n51;
  assign nan_mts_l2n26 = nan_flag_l1[52] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:874" *) nan_mts_l1n52 : nan_mts_l1n53;
  assign nan_mts_l2n27 = nan_flag_l1[54] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:875" *) nan_mts_l1n54 : nan_mts_l1n55;
  assign nan_mts_l2n28 = nan_flag_l1[56] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:876" *) nan_mts_l1n56 : nan_mts_l1n57;
  assign nan_mts_l2n29 = nan_flag_l1[58] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:877" *) nan_mts_l1n58 : nan_mts_l1n59;
  assign nan_mts_l2n30 = nan_flag_l1[60] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:878" *) nan_mts_l1n60 : nan_mts_l1n61;
  assign nan_mts_l2n31 = nan_flag_l1[62] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:879" *) nan_mts_l1n62 : nan_mts_l1n63;
  assign nan_mts_l3n0 = nan_flag_l2[0] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:952" *) nan_mts_l2n0 : nan_mts_l2n1;
  assign nan_mts_l3n1 = nan_flag_l2[2] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:953" *) nan_mts_l2n2 : nan_mts_l2n3;
  assign nan_mts_l3n2 = nan_flag_l2[4] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:954" *) nan_mts_l2n4 : nan_mts_l2n5;
  assign nan_mts_l3n3 = nan_flag_l2[6] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:955" *) nan_mts_l2n6 : nan_mts_l2n7;
  assign nan_mts_l3n4 = nan_flag_l2[8] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:956" *) nan_mts_l2n8 : nan_mts_l2n9;
  assign nan_mts_l3n5 = nan_flag_l2[10] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:957" *) nan_mts_l2n10 : nan_mts_l2n11;
  assign nan_mts_l3n6 = nan_flag_l2[12] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:958" *) nan_mts_l2n12 : nan_mts_l2n13;
  assign nan_mts_l3n7 = nan_flag_l2[14] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:959" *) nan_mts_l2n14 : nan_mts_l2n15;
  assign nan_mts_l3n8 = nan_flag_l2[16] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:960" *) nan_mts_l2n16 : nan_mts_l2n17;
  assign nan_mts_l3n9 = nan_flag_l2[18] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:961" *) nan_mts_l2n18 : nan_mts_l2n19;
  assign nan_mts_l3n10 = nan_flag_l2[20] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:962" *) nan_mts_l2n20 : nan_mts_l2n21;
  assign nan_mts_l3n11 = nan_flag_l2[22] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:963" *) nan_mts_l2n22 : nan_mts_l2n23;
  assign nan_mts_l3n12 = nan_flag_l2[24] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:964" *) nan_mts_l2n24 : nan_mts_l2n25;
  assign nan_mts_l3n13 = nan_flag_l2[26] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:965" *) nan_mts_l2n26 : nan_mts_l2n27;
  assign nan_mts_l3n14 = nan_flag_l2[28] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:966" *) nan_mts_l2n28 : nan_mts_l2n29;
  assign nan_mts_l3n15 = nan_flag_l2[30] ? (* src = "./vmod/nvdla/cmac/NV_NVDLA_CMAC_CORE_MAC_nan.v:967" *) nan_mts_l2n30 : nan_mts_l2n31;
  assign cur_data = { dat_actv_data, wt_actv_data };
  assign nan_mts_l0n0 = { wt_actv_data[15], wt_actv_data[12:3] };
  assign nan_mts_l0n1 = { wt_actv_data[31], wt_actv_data[28:19] };
  assign nan_mts_l0n10 = { wt_actv_data[175], wt_actv_data[172:163] };
  assign nan_mts_l0n100 = { dat_actv_data[591], dat_actv_data[588:579] };
  assign nan_mts_l0n101 = { dat_actv_data[607], dat_actv_data[604:595] };
  assign nan_mts_l0n102 = { dat_actv_data[623], dat_actv_data[620:611] };
  assign nan_mts_l0n103 = { dat_actv_data[639], dat_actv_data[636:627] };
  assign nan_mts_l0n104 = { dat_actv_data[655], dat_actv_data[652:643] };
  assign nan_mts_l0n105 = { dat_actv_data[671], dat_actv_data[668:659] };
  assign nan_mts_l0n106 = { dat_actv_data[687], dat_actv_data[684:675] };
  assign nan_mts_l0n107 = { dat_actv_data[703], dat_actv_data[700:691] };
  assign nan_mts_l0n108 = { dat_actv_data[719], dat_actv_data[716:707] };
  assign nan_mts_l0n109 = { dat_actv_data[735], dat_actv_data[732:723] };
  assign nan_mts_l0n11 = { wt_actv_data[191], wt_actv_data[188:179] };
  assign nan_mts_l0n110 = { dat_actv_data[751], dat_actv_data[748:739] };
  assign nan_mts_l0n111 = { dat_actv_data[767], dat_actv_data[764:755] };
  assign nan_mts_l0n112 = { dat_actv_data[783], dat_actv_data[780:771] };
  assign nan_mts_l0n113 = { dat_actv_data[799], dat_actv_data[796:787] };
  assign nan_mts_l0n114 = { dat_actv_data[815], dat_actv_data[812:803] };
  assign nan_mts_l0n115 = { dat_actv_data[831], dat_actv_data[828:819] };
  assign nan_mts_l0n116 = { dat_actv_data[847], dat_actv_data[844:835] };
  assign nan_mts_l0n117 = { dat_actv_data[863], dat_actv_data[860:851] };
  assign nan_mts_l0n118 = { dat_actv_data[879], dat_actv_data[876:867] };
  assign nan_mts_l0n119 = { dat_actv_data[895], dat_actv_data[892:883] };
  assign nan_mts_l0n12 = { wt_actv_data[207], wt_actv_data[204:195] };
  assign nan_mts_l0n120 = { dat_actv_data[911], dat_actv_data[908:899] };
  assign nan_mts_l0n121 = { dat_actv_data[927], dat_actv_data[924:915] };
  assign nan_mts_l0n122 = { dat_actv_data[943], dat_actv_data[940:931] };
  assign nan_mts_l0n123 = { dat_actv_data[959], dat_actv_data[956:947] };
  assign nan_mts_l0n124 = { dat_actv_data[975], dat_actv_data[972:963] };
  assign nan_mts_l0n125 = { dat_actv_data[991], dat_actv_data[988:979] };
  assign nan_mts_l0n126 = { dat_actv_data[1007], dat_actv_data[1004:995] };
  assign nan_mts_l0n127 = { dat_actv_data[1023], dat_actv_data[1020:1011] };
  assign nan_mts_l0n13 = { wt_actv_data[223], wt_actv_data[220:211] };
  assign nan_mts_l0n14 = { wt_actv_data[239], wt_actv_data[236:227] };
  assign nan_mts_l0n15 = { wt_actv_data[255], wt_actv_data[252:243] };
  assign nan_mts_l0n16 = { wt_actv_data[271], wt_actv_data[268:259] };
  assign nan_mts_l0n17 = { wt_actv_data[287], wt_actv_data[284:275] };
  assign nan_mts_l0n18 = { wt_actv_data[303], wt_actv_data[300:291] };
  assign nan_mts_l0n19 = { wt_actv_data[319], wt_actv_data[316:307] };
  assign nan_mts_l0n2 = { wt_actv_data[47], wt_actv_data[44:35] };
  assign nan_mts_l0n20 = { wt_actv_data[335], wt_actv_data[332:323] };
  assign nan_mts_l0n21 = { wt_actv_data[351], wt_actv_data[348:339] };
  assign nan_mts_l0n22 = { wt_actv_data[367], wt_actv_data[364:355] };
  assign nan_mts_l0n23 = { wt_actv_data[383], wt_actv_data[380:371] };
  assign nan_mts_l0n24 = { wt_actv_data[399], wt_actv_data[396:387] };
  assign nan_mts_l0n25 = { wt_actv_data[415], wt_actv_data[412:403] };
  assign nan_mts_l0n26 = { wt_actv_data[431], wt_actv_data[428:419] };
  assign nan_mts_l0n27 = { wt_actv_data[447], wt_actv_data[444:435] };
  assign nan_mts_l0n28 = { wt_actv_data[463], wt_actv_data[460:451] };
  assign nan_mts_l0n29 = { wt_actv_data[479], wt_actv_data[476:467] };
  assign nan_mts_l0n3 = { wt_actv_data[63], wt_actv_data[60:51] };
  assign nan_mts_l0n30 = { wt_actv_data[495], wt_actv_data[492:483] };
  assign nan_mts_l0n31 = { wt_actv_data[511], wt_actv_data[508:499] };
  assign nan_mts_l0n32 = { wt_actv_data[527], wt_actv_data[524:515] };
  assign nan_mts_l0n33 = { wt_actv_data[543], wt_actv_data[540:531] };
  assign nan_mts_l0n34 = { wt_actv_data[559], wt_actv_data[556:547] };
  assign nan_mts_l0n35 = { wt_actv_data[575], wt_actv_data[572:563] };
  assign nan_mts_l0n36 = { wt_actv_data[591], wt_actv_data[588:579] };
  assign nan_mts_l0n37 = { wt_actv_data[607], wt_actv_data[604:595] };
  assign nan_mts_l0n38 = { wt_actv_data[623], wt_actv_data[620:611] };
  assign nan_mts_l0n39 = { wt_actv_data[639], wt_actv_data[636:627] };
  assign nan_mts_l0n4 = { wt_actv_data[79], wt_actv_data[76:67] };
  assign nan_mts_l0n40 = { wt_actv_data[655], wt_actv_data[652:643] };
  assign nan_mts_l0n41 = { wt_actv_data[671], wt_actv_data[668:659] };
  assign nan_mts_l0n42 = { wt_actv_data[687], wt_actv_data[684:675] };
  assign nan_mts_l0n43 = { wt_actv_data[703], wt_actv_data[700:691] };
  assign nan_mts_l0n44 = { wt_actv_data[719], wt_actv_data[716:707] };
  assign nan_mts_l0n45 = { wt_actv_data[735], wt_actv_data[732:723] };
  assign nan_mts_l0n46 = { wt_actv_data[751], wt_actv_data[748:739] };
  assign nan_mts_l0n47 = { wt_actv_data[767], wt_actv_data[764:755] };
  assign nan_mts_l0n48 = { wt_actv_data[783], wt_actv_data[780:771] };
  assign nan_mts_l0n49 = { wt_actv_data[799], wt_actv_data[796:787] };
  assign nan_mts_l0n5 = { wt_actv_data[95], wt_actv_data[92:83] };
  assign nan_mts_l0n50 = { wt_actv_data[815], wt_actv_data[812:803] };
  assign nan_mts_l0n51 = { wt_actv_data[831], wt_actv_data[828:819] };
  assign nan_mts_l0n52 = { wt_actv_data[847], wt_actv_data[844:835] };
  assign nan_mts_l0n53 = { wt_actv_data[863], wt_actv_data[860:851] };
  assign nan_mts_l0n54 = { wt_actv_data[879], wt_actv_data[876:867] };
  assign nan_mts_l0n55 = { wt_actv_data[895], wt_actv_data[892:883] };
  assign nan_mts_l0n56 = { wt_actv_data[911], wt_actv_data[908:899] };
  assign nan_mts_l0n57 = { wt_actv_data[927], wt_actv_data[924:915] };
  assign nan_mts_l0n58 = { wt_actv_data[943], wt_actv_data[940:931] };
  assign nan_mts_l0n59 = { wt_actv_data[959], wt_actv_data[956:947] };
  assign nan_mts_l0n6 = { wt_actv_data[111], wt_actv_data[108:99] };
  assign nan_mts_l0n60 = { wt_actv_data[975], wt_actv_data[972:963] };
  assign nan_mts_l0n61 = { wt_actv_data[991], wt_actv_data[988:979] };
  assign nan_mts_l0n62 = { wt_actv_data[1007], wt_actv_data[1004:995] };
  assign nan_mts_l0n63 = { wt_actv_data[1023], wt_actv_data[1020:1011] };
  assign nan_mts_l0n64 = { dat_actv_data[15], dat_actv_data[12:3] };
  assign nan_mts_l0n65 = { dat_actv_data[31], dat_actv_data[28:19] };
  assign nan_mts_l0n66 = { dat_actv_data[47], dat_actv_data[44:35] };
  assign nan_mts_l0n67 = { dat_actv_data[63], dat_actv_data[60:51] };
  assign nan_mts_l0n68 = { dat_actv_data[79], dat_actv_data[76:67] };
  assign nan_mts_l0n69 = { dat_actv_data[95], dat_actv_data[92:83] };
  assign nan_mts_l0n7 = { wt_actv_data[127], wt_actv_data[124:115] };
  assign nan_mts_l0n70 = { dat_actv_data[111], dat_actv_data[108:99] };
  assign nan_mts_l0n71 = { dat_actv_data[127], dat_actv_data[124:115] };
  assign nan_mts_l0n72 = { dat_actv_data[143], dat_actv_data[140:131] };
  assign nan_mts_l0n73 = { dat_actv_data[159], dat_actv_data[156:147] };
  assign nan_mts_l0n74 = { dat_actv_data[175], dat_actv_data[172:163] };
  assign nan_mts_l0n75 = { dat_actv_data[191], dat_actv_data[188:179] };
  assign nan_mts_l0n76 = { dat_actv_data[207], dat_actv_data[204:195] };
  assign nan_mts_l0n77 = { dat_actv_data[223], dat_actv_data[220:211] };
  assign nan_mts_l0n78 = { dat_actv_data[239], dat_actv_data[236:227] };
  assign nan_mts_l0n79 = { dat_actv_data[255], dat_actv_data[252:243] };
  assign nan_mts_l0n8 = { wt_actv_data[143], wt_actv_data[140:131] };
  assign nan_mts_l0n80 = { dat_actv_data[271], dat_actv_data[268:259] };
  assign nan_mts_l0n81 = { dat_actv_data[287], dat_actv_data[284:275] };
  assign nan_mts_l0n82 = { dat_actv_data[303], dat_actv_data[300:291] };
  assign nan_mts_l0n83 = { dat_actv_data[319], dat_actv_data[316:307] };
  assign nan_mts_l0n84 = { dat_actv_data[335], dat_actv_data[332:323] };
  assign nan_mts_l0n85 = { dat_actv_data[351], dat_actv_data[348:339] };
  assign nan_mts_l0n86 = { dat_actv_data[367], dat_actv_data[364:355] };
  assign nan_mts_l0n87 = { dat_actv_data[383], dat_actv_data[380:371] };
  assign nan_mts_l0n88 = { dat_actv_data[399], dat_actv_data[396:387] };
  assign nan_mts_l0n89 = { dat_actv_data[415], dat_actv_data[412:403] };
  assign nan_mts_l0n9 = { wt_actv_data[159], wt_actv_data[156:147] };
  assign nan_mts_l0n90 = { dat_actv_data[431], dat_actv_data[428:419] };
  assign nan_mts_l0n91 = { dat_actv_data[447], dat_actv_data[444:435] };
  assign nan_mts_l0n92 = { dat_actv_data[463], dat_actv_data[460:451] };
  assign nan_mts_l0n93 = { dat_actv_data[479], dat_actv_data[476:467] };
  assign nan_mts_l0n94 = { dat_actv_data[495], dat_actv_data[492:483] };
  assign nan_mts_l0n95 = { dat_actv_data[511], dat_actv_data[508:499] };
  assign nan_mts_l0n96 = { dat_actv_data[527], dat_actv_data[524:515] };
  assign nan_mts_l0n97 = { dat_actv_data[543], dat_actv_data[540:531] };
  assign nan_mts_l0n98 = { dat_actv_data[559], dat_actv_data[556:547] };
  assign nan_mts_l0n99 = { dat_actv_data[575], dat_actv_data[572:563] };
endmodule
