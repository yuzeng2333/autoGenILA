module SDP_X_cfg_mul_shift_value_rsc_triosy_obj_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:2107" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:2108" *)
  output outsig;
  assign outsig = in_0;
endmodule
