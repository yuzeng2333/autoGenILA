module AesEncrypt(clock, reset, io_dataIn, io_ivIn, io_dataValid, io_keys_0_0_0, io_keys_0_0_1, io_keys_0_0_2, io_keys_0_0_3, io_keys_0_1_0, io_keys_0_1_1, io_keys_0_1_2, io_keys_0_1_3, io_keys_0_2_0, io_keys_0_2_1, io_keys_0_2_2, io_keys_0_2_3, io_keys_0_3_0, io_keys_0_3_1, io_keys_0_3_2, io_keys_0_3_3, io_aes256, io_shiftCyc, io_shift, io_ready, io_dataOut, io_ivOut, io_outputValid);
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0000_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0001_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0002_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0003_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0004_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0005_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0006_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0007_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0008_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0009_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0010_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0011_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0012_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0013_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0014_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [7:0] _0015_;
  (* src = "crypto_accelerator.v:2979" *)
  wire [5:0] _0016_;
  wire [7:0] _0017_;
  wire [7:0] _0018_;
  wire [7:0] _0019_;
  wire [7:0] _0020_;
  wire [7:0] _0021_;
  wire [7:0] _0022_;
  wire [7:0] _0023_;
  wire [7:0] _0024_;
  wire [7:0] _0025_;
  wire [7:0] _0026_;
  wire [7:0] _0027_;
  wire [7:0] _0028_;
  wire [7:0] _0029_;
  wire [7:0] _0030_;
  wire [7:0] _0031_;
  wire [7:0] _0032_;
  wire [7:0] _0033_;
  wire [7:0] _0034_;
  wire [7:0] _0035_;
  wire [7:0] _0036_;
  wire [7:0] _0037_;
  wire [7:0] _0038_;
  wire [7:0] _0039_;
  wire [7:0] _0040_;
  wire [7:0] _0041_;
  wire [7:0] _0042_;
  wire [7:0] _0043_;
  wire [7:0] _0044_;
  wire [7:0] _0045_;
  wire [7:0] _0046_;
  wire [7:0] _0047_;
  wire [7:0] _0048_;
  wire [7:0] _0049_;
  wire [7:0] _0050_;
  wire [7:0] _0051_;
  wire [7:0] _0052_;
  wire [7:0] _0053_;
  wire [7:0] _0054_;
  wire [7:0] _0055_;
  wire [7:0] _0056_;
  wire [7:0] _0057_;
  wire [7:0] _0058_;
  wire [7:0] _0059_;
  wire [7:0] _0060_;
  wire [7:0] _0061_;
  wire [7:0] _0062_;
  wire [7:0] _0063_;
  wire [7:0] _0064_;
  wire [5:0] _0065_;
  wire [5:0] _0066_;
  wire [5:0] _0067_;
  (* src = "crypto_accelerator.v:652" *)
  wire [7:0] MixColsModule_io_in_0_0;
  (* src = "crypto_accelerator.v:653" *)
  wire [7:0] MixColsModule_io_in_0_1;
  (* src = "crypto_accelerator.v:654" *)
  wire [7:0] MixColsModule_io_in_0_2;
  (* src = "crypto_accelerator.v:655" *)
  wire [7:0] MixColsModule_io_in_0_3;
  (* src = "crypto_accelerator.v:656" *)
  wire [7:0] MixColsModule_io_in_1_0;
  (* src = "crypto_accelerator.v:657" *)
  wire [7:0] MixColsModule_io_in_1_1;
  (* src = "crypto_accelerator.v:658" *)
  wire [7:0] MixColsModule_io_in_1_2;
  (* src = "crypto_accelerator.v:659" *)
  wire [7:0] MixColsModule_io_in_1_3;
  (* src = "crypto_accelerator.v:660" *)
  wire [7:0] MixColsModule_io_in_2_0;
  (* src = "crypto_accelerator.v:661" *)
  wire [7:0] MixColsModule_io_in_2_1;
  (* src = "crypto_accelerator.v:662" *)
  wire [7:0] MixColsModule_io_in_2_2;
  (* src = "crypto_accelerator.v:663" *)
  wire [7:0] MixColsModule_io_in_2_3;
  (* src = "crypto_accelerator.v:664" *)
  wire [7:0] MixColsModule_io_in_3_0;
  (* src = "crypto_accelerator.v:665" *)
  wire [7:0] MixColsModule_io_in_3_1;
  (* src = "crypto_accelerator.v:666" *)
  wire [7:0] MixColsModule_io_in_3_2;
  (* src = "crypto_accelerator.v:667" *)
  wire [7:0] MixColsModule_io_in_3_3;
  (* src = "crypto_accelerator.v:668" *)
  wire [7:0] MixColsModule_io_out_0_0;
  (* src = "crypto_accelerator.v:669" *)
  wire [7:0] MixColsModule_io_out_0_1;
  (* src = "crypto_accelerator.v:670" *)
  wire [7:0] MixColsModule_io_out_0_2;
  (* src = "crypto_accelerator.v:671" *)
  wire [7:0] MixColsModule_io_out_0_3;
  (* src = "crypto_accelerator.v:672" *)
  wire [7:0] MixColsModule_io_out_1_0;
  (* src = "crypto_accelerator.v:673" *)
  wire [7:0] MixColsModule_io_out_1_1;
  (* src = "crypto_accelerator.v:674" *)
  wire [7:0] MixColsModule_io_out_1_2;
  (* src = "crypto_accelerator.v:675" *)
  wire [7:0] MixColsModule_io_out_1_3;
  (* src = "crypto_accelerator.v:676" *)
  wire [7:0] MixColsModule_io_out_2_0;
  (* src = "crypto_accelerator.v:677" *)
  wire [7:0] MixColsModule_io_out_2_1;
  (* src = "crypto_accelerator.v:678" *)
  wire [7:0] MixColsModule_io_out_2_2;
  (* src = "crypto_accelerator.v:679" *)
  wire [7:0] MixColsModule_io_out_2_3;
  (* src = "crypto_accelerator.v:680" *)
  wire [7:0] MixColsModule_io_out_3_0;
  (* src = "crypto_accelerator.v:681" *)
  wire [7:0] MixColsModule_io_out_3_1;
  (* src = "crypto_accelerator.v:682" *)
  wire [7:0] MixColsModule_io_out_3_2;
  (* src = "crypto_accelerator.v:683" *)
  wire [7:0] MixColsModule_io_out_3_3;
  (* src = "crypto_accelerator.v:2845" *)
  wire _GEN_34;
  (* src = "crypto_accelerator.v:685" *)
  wire _T;
  (* src = "crypto_accelerator.v:686" *)
  wire _T_1;
  (* src = "crypto_accelerator.v:1175" *)
  wire _T_1000;
  (* src = "crypto_accelerator.v:1176" *)
  wire _T_1002;
  (* src = "crypto_accelerator.v:1177" *)
  wire _T_1004;
  (* src = "crypto_accelerator.v:1178" *)
  wire _T_1006;
  (* src = "crypto_accelerator.v:1179" *)
  wire _T_1008;
  (* src = "crypto_accelerator.v:739" *)
  wire _T_101;
  (* src = "crypto_accelerator.v:1180" *)
  wire _T_1010;
  (* src = "crypto_accelerator.v:1181" *)
  wire _T_1012;
  (* src = "crypto_accelerator.v:1182" *)
  wire _T_1014;
  (* src = "crypto_accelerator.v:1183" *)
  wire _T_1016;
  (* src = "crypto_accelerator.v:1184" *)
  wire _T_1018;
  (* src = "crypto_accelerator.v:1185" *)
  wire _T_1020;
  (* src = "crypto_accelerator.v:1186" *)
  wire _T_1022;
  (* src = "crypto_accelerator.v:1187" *)
  wire _T_1024;
  (* src = "crypto_accelerator.v:1188" *)
  wire _T_1026;
  (* src = "crypto_accelerator.v:1189" *)
  wire _T_1028;
  (* src = "crypto_accelerator.v:740" *)
  wire _T_103;
  (* src = "crypto_accelerator.v:1190" *)
  wire _T_1030;
  (* src = "crypto_accelerator.v:1191" *)
  wire _T_1032;
  (* src = "crypto_accelerator.v:1192" *)
  wire _T_1034;
  (* src = "crypto_accelerator.v:1193" *)
  wire _T_1036;
  (* src = "crypto_accelerator.v:1194" *)
  wire _T_1038;
  (* src = "crypto_accelerator.v:1195" *)
  wire _T_1040;
  (* src = "crypto_accelerator.v:1196" *)
  wire _T_1042;
  (* src = "crypto_accelerator.v:1197" *)
  wire _T_1044;
  (* src = "crypto_accelerator.v:1198" *)
  wire _T_1046;
  (* src = "crypto_accelerator.v:1199" *)
  wire _T_1048;
  (* src = "crypto_accelerator.v:741" *)
  wire _T_105;
  (* src = "crypto_accelerator.v:1200" *)
  wire _T_1050;
  (* src = "crypto_accelerator.v:1201" *)
  wire _T_1052;
  (* src = "crypto_accelerator.v:1202" *)
  wire _T_1054;
  (* src = "crypto_accelerator.v:1203" *)
  wire _T_1056;
  (* src = "crypto_accelerator.v:1204" *)
  wire _T_1058;
  (* src = "crypto_accelerator.v:1205" *)
  wire _T_1060;
  (* src = "crypto_accelerator.v:1206" *)
  wire _T_1062;
  (* src = "crypto_accelerator.v:1207" *)
  wire _T_1064;
  (* src = "crypto_accelerator.v:1208" *)
  wire _T_1066;
  (* src = "crypto_accelerator.v:1209" *)
  wire _T_1068;
  (* src = "crypto_accelerator.v:742" *)
  wire _T_107;
  (* src = "crypto_accelerator.v:1210" *)
  wire _T_1070;
  (* src = "crypto_accelerator.v:1211" *)
  wire _T_1072;
  (* src = "crypto_accelerator.v:1212" *)
  wire _T_1074;
  (* src = "crypto_accelerator.v:1213" *)
  wire _T_1076;
  (* src = "crypto_accelerator.v:1214" *)
  wire _T_1078;
  (* src = "crypto_accelerator.v:1215" *)
  wire _T_1080;
  (* src = "crypto_accelerator.v:1216" *)
  wire _T_1082;
  (* src = "crypto_accelerator.v:1217" *)
  wire _T_1084;
  (* src = "crypto_accelerator.v:1218" *)
  wire _T_1086;
  (* src = "crypto_accelerator.v:1219" *)
  wire _T_1088;
  (* src = "crypto_accelerator.v:743" *)
  wire _T_109;
  (* src = "crypto_accelerator.v:1220" *)
  wire _T_1090;
  (* src = "crypto_accelerator.v:1221" *)
  wire _T_1092;
  (* src = "crypto_accelerator.v:1222" *)
  wire _T_1094;
  (* src = "crypto_accelerator.v:1223" *)
  wire _T_1096;
  (* src = "crypto_accelerator.v:1224" *)
  wire _T_1098;
  (* src = "crypto_accelerator.v:1225" *)
  wire _T_1100;
  (* src = "crypto_accelerator.v:1226" *)
  wire _T_1102;
  (* src = "crypto_accelerator.v:1227" *)
  wire _T_1103;
  (* src = "crypto_accelerator.v:1228" *)
  wire _T_1104;
  (* src = "crypto_accelerator.v:1229" *)
  wire _T_1105;
  (* src = "crypto_accelerator.v:1230" *)
  wire _T_1107;
  (* src = "crypto_accelerator.v:1231" *)
  wire _T_1108;
  (* src = "crypto_accelerator.v:1232" *)
  wire _T_1109;
  (* src = "crypto_accelerator.v:744" *)
  wire _T_111;
  (* src = "crypto_accelerator.v:1233" *)
  wire _T_1111;
  (* src = "crypto_accelerator.v:1234" *)
  wire _T_1113;
  (* src = "crypto_accelerator.v:1235" *)
  wire _T_1114;
  (* src = "crypto_accelerator.v:1236" *)
  wire _T_1115;
  (* src = "crypto_accelerator.v:1237" *)
  wire _T_1117;
  (* src = "crypto_accelerator.v:1238" *)
  wire _T_1119;
  (* src = "crypto_accelerator.v:1239" *)
  wire _T_1121;
  (* src = "crypto_accelerator.v:1240" *)
  wire _T_1122;
  (* src = "crypto_accelerator.v:1241" *)
  wire _T_1123;
  (* src = "crypto_accelerator.v:1242" *)
  wire _T_1125;
  (* src = "crypto_accelerator.v:1243" *)
  wire _T_1126;
  (* src = "crypto_accelerator.v:1244" *)
  wire _T_1128;
  (* src = "crypto_accelerator.v:1245" *)
  wire _T_1129;
  (* src = "crypto_accelerator.v:745" *)
  wire _T_113;
  (* src = "crypto_accelerator.v:1246" *)
  wire _T_1130;
  (* src = "crypto_accelerator.v:746" *)
  wire _T_115;
  (* src = "crypto_accelerator.v:1248" *)
  wire _T_1156;
  (* src = "crypto_accelerator.v:1249" *)
  wire _T_1158;
  (* src = "crypto_accelerator.v:1250" *)
  wire _T_1160;
  (* src = "crypto_accelerator.v:1251" *)
  wire _T_1162;
  (* src = "crypto_accelerator.v:1252" *)
  wire _T_1164;
  (* src = "crypto_accelerator.v:1253" *)
  wire _T_1166;
  (* src = "crypto_accelerator.v:1254" *)
  wire _T_1168;
  (* src = "crypto_accelerator.v:747" *)
  wire _T_117;
  (* src = "crypto_accelerator.v:1255" *)
  wire _T_1170;
  (* src = "crypto_accelerator.v:1256" *)
  wire _T_1172;
  (* src = "crypto_accelerator.v:1257" *)
  wire _T_1174;
  (* src = "crypto_accelerator.v:1258" *)
  wire _T_1176;
  (* src = "crypto_accelerator.v:1259" *)
  wire _T_1178;
  (* src = "crypto_accelerator.v:1260" *)
  wire _T_1180;
  (* src = "crypto_accelerator.v:1261" *)
  wire _T_1182;
  (* src = "crypto_accelerator.v:1262" *)
  wire _T_1184;
  (* src = "crypto_accelerator.v:1263" *)
  wire _T_1186;
  (* src = "crypto_accelerator.v:1264" *)
  wire _T_1188;
  (* src = "crypto_accelerator.v:748" *)
  wire _T_119;
  (* src = "crypto_accelerator.v:1265" *)
  wire _T_1190;
  (* src = "crypto_accelerator.v:1266" *)
  wire _T_1192;
  (* src = "crypto_accelerator.v:1267" *)
  wire _T_1194;
  (* src = "crypto_accelerator.v:1268" *)
  wire _T_1196;
  (* src = "crypto_accelerator.v:1269" *)
  wire _T_1198;
  (* src = "crypto_accelerator.v:1270" *)
  wire _T_1200;
  (* src = "crypto_accelerator.v:1271" *)
  wire _T_1202;
  (* src = "crypto_accelerator.v:1272" *)
  wire _T_1204;
  (* src = "crypto_accelerator.v:1273" *)
  wire _T_1206;
  (* src = "crypto_accelerator.v:1274" *)
  wire _T_1208;
  (* src = "crypto_accelerator.v:749" *)
  wire _T_121;
  (* src = "crypto_accelerator.v:1275" *)
  wire _T_1210;
  (* src = "crypto_accelerator.v:1276" *)
  wire _T_1212;
  (* src = "crypto_accelerator.v:1277" *)
  wire _T_1214;
  (* src = "crypto_accelerator.v:1278" *)
  wire _T_1216;
  (* src = "crypto_accelerator.v:1279" *)
  wire _T_1218;
  (* src = "crypto_accelerator.v:1280" *)
  wire _T_1220;
  (* src = "crypto_accelerator.v:1281" *)
  wire _T_1222;
  (* src = "crypto_accelerator.v:1282" *)
  wire _T_1224;
  (* src = "crypto_accelerator.v:1283" *)
  wire _T_1226;
  (* src = "crypto_accelerator.v:1284" *)
  wire _T_1228;
  (* src = "crypto_accelerator.v:750" *)
  wire _T_123;
  (* src = "crypto_accelerator.v:1285" *)
  wire _T_1230;
  (* src = "crypto_accelerator.v:1286" *)
  wire _T_1232;
  (* src = "crypto_accelerator.v:1287" *)
  wire _T_1234;
  (* src = "crypto_accelerator.v:1288" *)
  wire _T_1236;
  (* src = "crypto_accelerator.v:1289" *)
  wire _T_1238;
  (* src = "crypto_accelerator.v:1290" *)
  wire _T_1240;
  (* src = "crypto_accelerator.v:1291" *)
  wire _T_1242;
  (* src = "crypto_accelerator.v:1292" *)
  wire _T_1244;
  (* src = "crypto_accelerator.v:1293" *)
  wire _T_1246;
  (* src = "crypto_accelerator.v:1294" *)
  wire _T_1248;
  (* src = "crypto_accelerator.v:751" *)
  wire _T_125;
  (* src = "crypto_accelerator.v:1295" *)
  wire _T_1250;
  (* src = "crypto_accelerator.v:1296" *)
  wire _T_1252;
  (* src = "crypto_accelerator.v:1297" *)
  wire _T_1254;
  (* src = "crypto_accelerator.v:1298" *)
  wire _T_1256;
  (* src = "crypto_accelerator.v:1299" *)
  wire _T_1258;
  (* src = "crypto_accelerator.v:1300" *)
  wire _T_1260;
  (* src = "crypto_accelerator.v:1301" *)
  wire _T_1262;
  (* src = "crypto_accelerator.v:1302" *)
  wire _T_1264;
  (* src = "crypto_accelerator.v:1303" *)
  wire _T_1266;
  (* src = "crypto_accelerator.v:1304" *)
  wire _T_1268;
  (* src = "crypto_accelerator.v:752" *)
  wire _T_127;
  (* src = "crypto_accelerator.v:1305" *)
  wire _T_1270;
  (* src = "crypto_accelerator.v:1306" *)
  wire _T_1272;
  (* src = "crypto_accelerator.v:1307" *)
  wire _T_1274;
  (* src = "crypto_accelerator.v:1308" *)
  wire _T_1276;
  (* src = "crypto_accelerator.v:1309" *)
  wire _T_1278;
  (* src = "crypto_accelerator.v:1310" *)
  wire _T_1280;
  (* src = "crypto_accelerator.v:1311" *)
  wire _T_1282;
  (* src = "crypto_accelerator.v:1312" *)
  wire _T_1284;
  (* src = "crypto_accelerator.v:1313" *)
  wire _T_1286;
  (* src = "crypto_accelerator.v:1314" *)
  wire _T_1288;
  (* src = "crypto_accelerator.v:753" *)
  wire _T_129;
  (* src = "crypto_accelerator.v:1315" *)
  wire _T_1290;
  (* src = "crypto_accelerator.v:1316" *)
  wire _T_1292;
  (* src = "crypto_accelerator.v:1317" *)
  wire _T_1294;
  (* src = "crypto_accelerator.v:1318" *)
  wire _T_1296;
  (* src = "crypto_accelerator.v:1319" *)
  wire _T_1298;
  (* src = "crypto_accelerator.v:1320" *)
  wire _T_1300;
  (* src = "crypto_accelerator.v:1321" *)
  wire _T_1302;
  (* src = "crypto_accelerator.v:1322" *)
  wire _T_1304;
  (* src = "crypto_accelerator.v:1323" *)
  wire _T_1306;
  (* src = "crypto_accelerator.v:1324" *)
  wire _T_1308;
  (* src = "crypto_accelerator.v:754" *)
  wire _T_131;
  (* src = "crypto_accelerator.v:1325" *)
  wire _T_1310;
  (* src = "crypto_accelerator.v:1326" *)
  wire _T_1312;
  (* src = "crypto_accelerator.v:1327" *)
  wire _T_1314;
  (* src = "crypto_accelerator.v:1328" *)
  wire _T_1316;
  (* src = "crypto_accelerator.v:1329" *)
  wire _T_1318;
  (* src = "crypto_accelerator.v:1330" *)
  wire _T_1320;
  (* src = "crypto_accelerator.v:1331" *)
  wire _T_1322;
  (* src = "crypto_accelerator.v:1332" *)
  wire _T_1324;
  (* src = "crypto_accelerator.v:1333" *)
  wire _T_1326;
  (* src = "crypto_accelerator.v:1334" *)
  wire _T_1328;
  (* src = "crypto_accelerator.v:755" *)
  wire _T_133;
  (* src = "crypto_accelerator.v:1335" *)
  wire _T_1330;
  (* src = "crypto_accelerator.v:1336" *)
  wire _T_1332;
  (* src = "crypto_accelerator.v:1337" *)
  wire _T_1334;
  (* src = "crypto_accelerator.v:1338" *)
  wire _T_1336;
  (* src = "crypto_accelerator.v:1339" *)
  wire _T_1338;
  (* src = "crypto_accelerator.v:1340" *)
  wire _T_1340;
  (* src = "crypto_accelerator.v:1341" *)
  wire _T_1342;
  (* src = "crypto_accelerator.v:1342" *)
  wire _T_1344;
  (* src = "crypto_accelerator.v:1343" *)
  wire _T_1346;
  (* src = "crypto_accelerator.v:1344" *)
  wire _T_1348;
  (* src = "crypto_accelerator.v:756" *)
  wire _T_135;
  (* src = "crypto_accelerator.v:1345" *)
  wire _T_1350;
  (* src = "crypto_accelerator.v:1346" *)
  wire _T_1352;
  (* src = "crypto_accelerator.v:1347" *)
  wire _T_1354;
  (* src = "crypto_accelerator.v:1348" *)
  wire _T_1356;
  (* src = "crypto_accelerator.v:1349" *)
  wire _T_1358;
  (* src = "crypto_accelerator.v:1350" *)
  wire _T_1360;
  (* src = "crypto_accelerator.v:1351" *)
  wire _T_1362;
  (* src = "crypto_accelerator.v:1352" *)
  wire _T_1364;
  (* src = "crypto_accelerator.v:1353" *)
  wire _T_1366;
  (* src = "crypto_accelerator.v:1354" *)
  wire _T_1368;
  (* src = "crypto_accelerator.v:757" *)
  wire _T_137;
  (* src = "crypto_accelerator.v:1355" *)
  wire _T_1370;
  (* src = "crypto_accelerator.v:1356" *)
  wire _T_1372;
  (* src = "crypto_accelerator.v:1357" *)
  wire _T_1373;
  (* src = "crypto_accelerator.v:1358" *)
  wire _T_1374;
  (* src = "crypto_accelerator.v:1359" *)
  wire _T_1375;
  (* src = "crypto_accelerator.v:1360" *)
  wire _T_1377;
  (* src = "crypto_accelerator.v:1361" *)
  wire _T_1378;
  (* src = "crypto_accelerator.v:1362" *)
  wire _T_1379;
  (* src = "crypto_accelerator.v:1363" *)
  wire _T_1381;
  (* src = "crypto_accelerator.v:1364" *)
  wire _T_1383;
  (* src = "crypto_accelerator.v:1365" *)
  wire _T_1384;
  (* src = "crypto_accelerator.v:1366" *)
  wire _T_1385;
  (* src = "crypto_accelerator.v:1367" *)
  wire _T_1387;
  (* src = "crypto_accelerator.v:1368" *)
  wire _T_1389;
  (* src = "crypto_accelerator.v:758" *)
  wire _T_139;
  (* src = "crypto_accelerator.v:1369" *)
  wire _T_1391;
  (* src = "crypto_accelerator.v:1370" *)
  wire _T_1392;
  (* src = "crypto_accelerator.v:1371" *)
  wire _T_1393;
  (* src = "crypto_accelerator.v:1372" *)
  wire _T_1395;
  (* src = "crypto_accelerator.v:1373" *)
  wire _T_1396;
  (* src = "crypto_accelerator.v:1374" *)
  wire _T_1398;
  (* src = "crypto_accelerator.v:1375" *)
  wire _T_1399;
  (* src = "crypto_accelerator.v:1376" *)
  wire _T_1400;
  (* src = "crypto_accelerator.v:759" *)
  wire _T_141;
  (* src = "crypto_accelerator.v:1378" *)
  wire _T_1425;
  (* src = "crypto_accelerator.v:1379" *)
  wire _T_1427;
  (* src = "crypto_accelerator.v:1380" *)
  wire _T_1429;
  (* src = "crypto_accelerator.v:760" *)
  wire _T_143;
  (* src = "crypto_accelerator.v:1381" *)
  wire _T_1431;
  (* src = "crypto_accelerator.v:1382" *)
  wire _T_1433;
  (* src = "crypto_accelerator.v:1383" *)
  wire _T_1435;
  (* src = "crypto_accelerator.v:1384" *)
  wire _T_1437;
  (* src = "crypto_accelerator.v:1385" *)
  wire _T_1439;
  (* src = "crypto_accelerator.v:1386" *)
  wire _T_1441;
  (* src = "crypto_accelerator.v:1387" *)
  wire _T_1443;
  (* src = "crypto_accelerator.v:1388" *)
  wire _T_1445;
  (* src = "crypto_accelerator.v:1389" *)
  wire _T_1447;
  (* src = "crypto_accelerator.v:1390" *)
  wire _T_1449;
  (* src = "crypto_accelerator.v:761" *)
  wire _T_145;
  (* src = "crypto_accelerator.v:1391" *)
  wire _T_1451;
  (* src = "crypto_accelerator.v:1392" *)
  wire _T_1453;
  (* src = "crypto_accelerator.v:1393" *)
  wire _T_1455;
  (* src = "crypto_accelerator.v:1394" *)
  wire _T_1457;
  (* src = "crypto_accelerator.v:1395" *)
  wire _T_1459;
  (* src = "crypto_accelerator.v:1396" *)
  wire _T_1461;
  (* src = "crypto_accelerator.v:1397" *)
  wire _T_1463;
  (* src = "crypto_accelerator.v:1398" *)
  wire _T_1465;
  (* src = "crypto_accelerator.v:1399" *)
  wire _T_1467;
  (* src = "crypto_accelerator.v:1400" *)
  wire _T_1469;
  (* src = "crypto_accelerator.v:762" *)
  wire _T_147;
  (* src = "crypto_accelerator.v:1401" *)
  wire _T_1471;
  (* src = "crypto_accelerator.v:1402" *)
  wire _T_1473;
  (* src = "crypto_accelerator.v:1403" *)
  wire _T_1475;
  (* src = "crypto_accelerator.v:1404" *)
  wire _T_1477;
  (* src = "crypto_accelerator.v:1405" *)
  wire _T_1479;
  (* src = "crypto_accelerator.v:1406" *)
  wire _T_1481;
  (* src = "crypto_accelerator.v:1407" *)
  wire _T_1483;
  (* src = "crypto_accelerator.v:1408" *)
  wire _T_1485;
  (* src = "crypto_accelerator.v:1409" *)
  wire _T_1487;
  (* src = "crypto_accelerator.v:1410" *)
  wire _T_1489;
  (* src = "crypto_accelerator.v:763" *)
  wire _T_149;
  (* src = "crypto_accelerator.v:1411" *)
  wire _T_1491;
  (* src = "crypto_accelerator.v:1412" *)
  wire _T_1493;
  (* src = "crypto_accelerator.v:1413" *)
  wire _T_1495;
  (* src = "crypto_accelerator.v:1414" *)
  wire _T_1497;
  (* src = "crypto_accelerator.v:1415" *)
  wire _T_1499;
  (* src = "crypto_accelerator.v:1416" *)
  wire _T_1501;
  (* src = "crypto_accelerator.v:1417" *)
  wire _T_1503;
  (* src = "crypto_accelerator.v:1418" *)
  wire _T_1505;
  (* src = "crypto_accelerator.v:1419" *)
  wire _T_1507;
  (* src = "crypto_accelerator.v:1420" *)
  wire _T_1509;
  (* src = "crypto_accelerator.v:764" *)
  wire _T_151;
  (* src = "crypto_accelerator.v:1421" *)
  wire _T_1511;
  (* src = "crypto_accelerator.v:1422" *)
  wire _T_1513;
  (* src = "crypto_accelerator.v:1423" *)
  wire _T_1515;
  (* src = "crypto_accelerator.v:1424" *)
  wire _T_1517;
  (* src = "crypto_accelerator.v:1425" *)
  wire _T_1519;
  (* src = "crypto_accelerator.v:1426" *)
  wire _T_1521;
  (* src = "crypto_accelerator.v:1427" *)
  wire _T_1523;
  (* src = "crypto_accelerator.v:1428" *)
  wire _T_1525;
  (* src = "crypto_accelerator.v:1429" *)
  wire _T_1527;
  (* src = "crypto_accelerator.v:1430" *)
  wire _T_1529;
  (* src = "crypto_accelerator.v:765" *)
  wire _T_153;
  (* src = "crypto_accelerator.v:1431" *)
  wire _T_1531;
  (* src = "crypto_accelerator.v:1432" *)
  wire _T_1533;
  (* src = "crypto_accelerator.v:1433" *)
  wire _T_1535;
  (* src = "crypto_accelerator.v:1434" *)
  wire _T_1537;
  (* src = "crypto_accelerator.v:1435" *)
  wire _T_1539;
  (* src = "crypto_accelerator.v:1436" *)
  wire _T_1541;
  (* src = "crypto_accelerator.v:1437" *)
  wire _T_1543;
  (* src = "crypto_accelerator.v:1438" *)
  wire _T_1545;
  (* src = "crypto_accelerator.v:1439" *)
  wire _T_1547;
  (* src = "crypto_accelerator.v:1440" *)
  wire _T_1549;
  (* src = "crypto_accelerator.v:766" *)
  wire _T_155;
  (* src = "crypto_accelerator.v:1441" *)
  wire _T_1551;
  (* src = "crypto_accelerator.v:1442" *)
  wire _T_1553;
  (* src = "crypto_accelerator.v:1443" *)
  wire _T_1555;
  (* src = "crypto_accelerator.v:1444" *)
  wire _T_1557;
  (* src = "crypto_accelerator.v:1445" *)
  wire _T_1559;
  (* src = "crypto_accelerator.v:1446" *)
  wire _T_1561;
  (* src = "crypto_accelerator.v:1447" *)
  wire _T_1563;
  (* src = "crypto_accelerator.v:1448" *)
  wire _T_1565;
  (* src = "crypto_accelerator.v:1449" *)
  wire _T_1567;
  (* src = "crypto_accelerator.v:1450" *)
  wire _T_1569;
  (* src = "crypto_accelerator.v:767" *)
  wire _T_157;
  (* src = "crypto_accelerator.v:1451" *)
  wire _T_1571;
  (* src = "crypto_accelerator.v:1452" *)
  wire _T_1573;
  (* src = "crypto_accelerator.v:1453" *)
  wire _T_1575;
  (* src = "crypto_accelerator.v:1454" *)
  wire _T_1577;
  (* src = "crypto_accelerator.v:1455" *)
  wire _T_1579;
  (* src = "crypto_accelerator.v:1456" *)
  wire _T_1581;
  (* src = "crypto_accelerator.v:1457" *)
  wire _T_1583;
  (* src = "crypto_accelerator.v:1458" *)
  wire _T_1585;
  (* src = "crypto_accelerator.v:1459" *)
  wire _T_1587;
  (* src = "crypto_accelerator.v:1460" *)
  wire _T_1589;
  (* src = "crypto_accelerator.v:768" *)
  wire _T_159;
  (* src = "crypto_accelerator.v:1461" *)
  wire _T_1591;
  (* src = "crypto_accelerator.v:1462" *)
  wire _T_1593;
  (* src = "crypto_accelerator.v:1463" *)
  wire _T_1595;
  (* src = "crypto_accelerator.v:1464" *)
  wire _T_1597;
  (* src = "crypto_accelerator.v:1465" *)
  wire _T_1599;
  (* src = "crypto_accelerator.v:706" *)
  wire [63:0] _T_16;
  (* src = "crypto_accelerator.v:1466" *)
  wire _T_1601;
  (* src = "crypto_accelerator.v:1467" *)
  wire _T_1603;
  (* src = "crypto_accelerator.v:1468" *)
  wire _T_1605;
  (* src = "crypto_accelerator.v:1469" *)
  wire _T_1607;
  (* src = "crypto_accelerator.v:1470" *)
  wire _T_1609;
  (* src = "crypto_accelerator.v:769" *)
  wire _T_161;
  (* src = "crypto_accelerator.v:1471" *)
  wire _T_1611;
  (* src = "crypto_accelerator.v:1472" *)
  wire _T_1613;
  (* src = "crypto_accelerator.v:1473" *)
  wire _T_1615;
  (* src = "crypto_accelerator.v:1474" *)
  wire _T_1617;
  (* src = "crypto_accelerator.v:1475" *)
  wire _T_1619;
  (* src = "crypto_accelerator.v:1476" *)
  wire _T_1621;
  (* src = "crypto_accelerator.v:1477" *)
  wire _T_1623;
  (* src = "crypto_accelerator.v:1478" *)
  wire _T_1625;
  (* src = "crypto_accelerator.v:1479" *)
  wire _T_1627;
  (* src = "crypto_accelerator.v:1480" *)
  wire _T_1629;
  (* src = "crypto_accelerator.v:770" *)
  wire _T_163;
  (* src = "crypto_accelerator.v:1481" *)
  wire _T_1631;
  (* src = "crypto_accelerator.v:1482" *)
  wire _T_1633;
  (* src = "crypto_accelerator.v:1483" *)
  wire _T_1635;
  (* src = "crypto_accelerator.v:1484" *)
  wire _T_1637;
  (* src = "crypto_accelerator.v:1485" *)
  wire _T_1639;
  (* src = "crypto_accelerator.v:1486" *)
  wire _T_1641;
  (* src = "crypto_accelerator.v:1487" *)
  wire _T_1642;
  (* src = "crypto_accelerator.v:1488" *)
  wire _T_1643;
  (* src = "crypto_accelerator.v:1489" *)
  wire _T_1644;
  (* src = "crypto_accelerator.v:1490" *)
  wire _T_1646;
  (* src = "crypto_accelerator.v:1491" *)
  wire _T_1647;
  (* src = "crypto_accelerator.v:1492" *)
  wire _T_1648;
  (* src = "crypto_accelerator.v:771" *)
  wire _T_165;
  (* src = "crypto_accelerator.v:1493" *)
  wire _T_1650;
  (* src = "crypto_accelerator.v:1494" *)
  wire _T_1652;
  (* src = "crypto_accelerator.v:1495" *)
  wire _T_1653;
  (* src = "crypto_accelerator.v:1496" *)
  wire _T_1654;
  (* src = "crypto_accelerator.v:1497" *)
  wire _T_1656;
  (* src = "crypto_accelerator.v:1498" *)
  wire _T_1658;
  (* src = "crypto_accelerator.v:1499" *)
  wire _T_1660;
  (* src = "crypto_accelerator.v:1500" *)
  wire _T_1661;
  (* src = "crypto_accelerator.v:1501" *)
  wire _T_1662;
  (* src = "crypto_accelerator.v:1502" *)
  wire _T_1664;
  (* src = "crypto_accelerator.v:1503" *)
  wire _T_1665;
  (* src = "crypto_accelerator.v:1504" *)
  wire _T_1667;
  (* src = "crypto_accelerator.v:1505" *)
  wire _T_1668;
  (* src = "crypto_accelerator.v:1506" *)
  wire _T_1669;
  (* src = "crypto_accelerator.v:772" *)
  wire _T_167;
  (* src = "crypto_accelerator.v:773" *)
  wire _T_169;
  (* src = "crypto_accelerator.v:1508" *)
  wire _T_1694;
  (* src = "crypto_accelerator.v:1509" *)
  wire _T_1696;
  (* src = "crypto_accelerator.v:1510" *)
  wire _T_1698;
  (* src = "crypto_accelerator.v:1511" *)
  wire _T_1700;
  (* src = "crypto_accelerator.v:1512" *)
  wire _T_1702;
  (* src = "crypto_accelerator.v:1513" *)
  wire _T_1704;
  (* src = "crypto_accelerator.v:1514" *)
  wire _T_1706;
  (* src = "crypto_accelerator.v:1515" *)
  wire _T_1708;
  (* src = "crypto_accelerator.v:774" *)
  wire _T_171;
  (* src = "crypto_accelerator.v:1516" *)
  wire _T_1710;
  (* src = "crypto_accelerator.v:1517" *)
  wire _T_1712;
  (* src = "crypto_accelerator.v:1518" *)
  wire _T_1714;
  (* src = "crypto_accelerator.v:1519" *)
  wire _T_1716;
  (* src = "crypto_accelerator.v:1520" *)
  wire _T_1718;
  (* src = "crypto_accelerator.v:1521" *)
  wire _T_1720;
  (* src = "crypto_accelerator.v:1522" *)
  wire _T_1722;
  (* src = "crypto_accelerator.v:1523" *)
  wire _T_1724;
  (* src = "crypto_accelerator.v:1524" *)
  wire _T_1726;
  (* src = "crypto_accelerator.v:1525" *)
  wire _T_1728;
  (* src = "crypto_accelerator.v:775" *)
  wire _T_173;
  (* src = "crypto_accelerator.v:1526" *)
  wire _T_1730;
  (* src = "crypto_accelerator.v:1527" *)
  wire _T_1732;
  (* src = "crypto_accelerator.v:1528" *)
  wire _T_1734;
  (* src = "crypto_accelerator.v:1529" *)
  wire _T_1736;
  (* src = "crypto_accelerator.v:1530" *)
  wire _T_1738;
  (* src = "crypto_accelerator.v:1531" *)
  wire _T_1740;
  (* src = "crypto_accelerator.v:1532" *)
  wire _T_1742;
  (* src = "crypto_accelerator.v:1533" *)
  wire _T_1744;
  (* src = "crypto_accelerator.v:1534" *)
  wire _T_1746;
  (* src = "crypto_accelerator.v:1535" *)
  wire _T_1748;
  (* src = "crypto_accelerator.v:776" *)
  wire _T_175;
  (* src = "crypto_accelerator.v:1536" *)
  wire _T_1750;
  (* src = "crypto_accelerator.v:1537" *)
  wire _T_1752;
  (* src = "crypto_accelerator.v:1538" *)
  wire _T_1754;
  (* src = "crypto_accelerator.v:1539" *)
  wire _T_1756;
  (* src = "crypto_accelerator.v:1540" *)
  wire _T_1758;
  (* src = "crypto_accelerator.v:1541" *)
  wire _T_1760;
  (* src = "crypto_accelerator.v:1542" *)
  wire _T_1762;
  (* src = "crypto_accelerator.v:1543" *)
  wire _T_1764;
  (* src = "crypto_accelerator.v:1544" *)
  wire _T_1766;
  (* src = "crypto_accelerator.v:1545" *)
  wire _T_1768;
  (* src = "crypto_accelerator.v:777" *)
  wire _T_177;
  (* src = "crypto_accelerator.v:1546" *)
  wire _T_1770;
  (* src = "crypto_accelerator.v:1547" *)
  wire _T_1772;
  (* src = "crypto_accelerator.v:1548" *)
  wire _T_1774;
  (* src = "crypto_accelerator.v:1549" *)
  wire _T_1776;
  (* src = "crypto_accelerator.v:1550" *)
  wire _T_1778;
  (* src = "crypto_accelerator.v:1551" *)
  wire _T_1780;
  (* src = "crypto_accelerator.v:1552" *)
  wire _T_1782;
  (* src = "crypto_accelerator.v:1553" *)
  wire _T_1784;
  (* src = "crypto_accelerator.v:1554" *)
  wire _T_1786;
  (* src = "crypto_accelerator.v:1555" *)
  wire _T_1788;
  (* src = "crypto_accelerator.v:778" *)
  wire _T_179;
  (* src = "crypto_accelerator.v:1556" *)
  wire _T_1790;
  (* src = "crypto_accelerator.v:1557" *)
  wire _T_1792;
  (* src = "crypto_accelerator.v:1558" *)
  wire _T_1794;
  (* src = "crypto_accelerator.v:1559" *)
  wire _T_1796;
  (* src = "crypto_accelerator.v:1560" *)
  wire _T_1798;
  (* src = "crypto_accelerator.v:1561" *)
  wire _T_1800;
  (* src = "crypto_accelerator.v:1562" *)
  wire _T_1802;
  (* src = "crypto_accelerator.v:1563" *)
  wire _T_1804;
  (* src = "crypto_accelerator.v:1564" *)
  wire _T_1806;
  (* src = "crypto_accelerator.v:1565" *)
  wire _T_1808;
  (* src = "crypto_accelerator.v:779" *)
  wire _T_181;
  (* src = "crypto_accelerator.v:1566" *)
  wire _T_1810;
  (* src = "crypto_accelerator.v:1567" *)
  wire _T_1812;
  (* src = "crypto_accelerator.v:1568" *)
  wire _T_1814;
  (* src = "crypto_accelerator.v:1569" *)
  wire _T_1816;
  (* src = "crypto_accelerator.v:1570" *)
  wire _T_1818;
  (* src = "crypto_accelerator.v:1571" *)
  wire _T_1820;
  (* src = "crypto_accelerator.v:1572" *)
  wire _T_1822;
  (* src = "crypto_accelerator.v:1573" *)
  wire _T_1824;
  (* src = "crypto_accelerator.v:1574" *)
  wire _T_1826;
  (* src = "crypto_accelerator.v:1575" *)
  wire _T_1828;
  (* src = "crypto_accelerator.v:780" *)
  wire _T_183;
  (* src = "crypto_accelerator.v:1576" *)
  wire _T_1830;
  (* src = "crypto_accelerator.v:1577" *)
  wire _T_1832;
  (* src = "crypto_accelerator.v:1578" *)
  wire _T_1834;
  (* src = "crypto_accelerator.v:1579" *)
  wire _T_1836;
  (* src = "crypto_accelerator.v:1580" *)
  wire _T_1838;
  (* src = "crypto_accelerator.v:1581" *)
  wire _T_1840;
  (* src = "crypto_accelerator.v:1582" *)
  wire _T_1842;
  (* src = "crypto_accelerator.v:1583" *)
  wire _T_1844;
  (* src = "crypto_accelerator.v:1584" *)
  wire _T_1846;
  (* src = "crypto_accelerator.v:1585" *)
  wire _T_1848;
  (* src = "crypto_accelerator.v:781" *)
  wire _T_185;
  (* src = "crypto_accelerator.v:1586" *)
  wire _T_1850;
  (* src = "crypto_accelerator.v:1587" *)
  wire _T_1852;
  (* src = "crypto_accelerator.v:1588" *)
  wire _T_1854;
  (* src = "crypto_accelerator.v:1589" *)
  wire _T_1856;
  (* src = "crypto_accelerator.v:1590" *)
  wire _T_1858;
  (* src = "crypto_accelerator.v:1591" *)
  wire _T_1860;
  (* src = "crypto_accelerator.v:1592" *)
  wire _T_1862;
  (* src = "crypto_accelerator.v:1593" *)
  wire _T_1864;
  (* src = "crypto_accelerator.v:1594" *)
  wire _T_1866;
  (* src = "crypto_accelerator.v:1595" *)
  wire _T_1868;
  (* src = "crypto_accelerator.v:782" *)
  wire _T_187;
  (* src = "crypto_accelerator.v:1596" *)
  wire _T_1870;
  (* src = "crypto_accelerator.v:1597" *)
  wire _T_1872;
  (* src = "crypto_accelerator.v:1598" *)
  wire _T_1874;
  (* src = "crypto_accelerator.v:1599" *)
  wire _T_1876;
  (* src = "crypto_accelerator.v:1600" *)
  wire _T_1878;
  (* src = "crypto_accelerator.v:1601" *)
  wire _T_1880;
  (* src = "crypto_accelerator.v:1602" *)
  wire _T_1882;
  (* src = "crypto_accelerator.v:1603" *)
  wire _T_1884;
  (* src = "crypto_accelerator.v:1604" *)
  wire _T_1886;
  (* src = "crypto_accelerator.v:1605" *)
  wire _T_1888;
  (* src = "crypto_accelerator.v:783" *)
  wire _T_189;
  (* src = "crypto_accelerator.v:1606" *)
  wire _T_1890;
  (* src = "crypto_accelerator.v:1607" *)
  wire _T_1892;
  (* src = "crypto_accelerator.v:1608" *)
  wire _T_1894;
  (* src = "crypto_accelerator.v:1609" *)
  wire _T_1896;
  (* src = "crypto_accelerator.v:1610" *)
  wire _T_1898;
  (* src = "crypto_accelerator.v:1611" *)
  wire _T_1900;
  (* src = "crypto_accelerator.v:1612" *)
  wire _T_1902;
  (* src = "crypto_accelerator.v:1613" *)
  wire _T_1904;
  (* src = "crypto_accelerator.v:1614" *)
  wire _T_1906;
  (* src = "crypto_accelerator.v:1615" *)
  wire _T_1908;
  (* src = "crypto_accelerator.v:784" *)
  wire _T_191;
  (* src = "crypto_accelerator.v:1616" *)
  wire _T_1910;
  (* src = "crypto_accelerator.v:1617" *)
  wire _T_1911;
  (* src = "crypto_accelerator.v:1618" *)
  wire _T_1912;
  (* src = "crypto_accelerator.v:1619" *)
  wire _T_1913;
  (* src = "crypto_accelerator.v:1620" *)
  wire _T_1915;
  (* src = "crypto_accelerator.v:1621" *)
  wire _T_1916;
  (* src = "crypto_accelerator.v:1622" *)
  wire _T_1917;
  (* src = "crypto_accelerator.v:1623" *)
  wire _T_1919;
  (* src = "crypto_accelerator.v:1624" *)
  wire _T_1921;
  (* src = "crypto_accelerator.v:1625" *)
  wire _T_1922;
  (* src = "crypto_accelerator.v:1626" *)
  wire _T_1923;
  (* src = "crypto_accelerator.v:1627" *)
  wire _T_1925;
  (* src = "crypto_accelerator.v:1628" *)
  wire _T_1927;
  (* src = "crypto_accelerator.v:1629" *)
  wire _T_1929;
  (* src = "crypto_accelerator.v:785" *)
  wire _T_193;
  (* src = "crypto_accelerator.v:1630" *)
  wire _T_1930;
  (* src = "crypto_accelerator.v:1631" *)
  wire _T_1931;
  (* src = "crypto_accelerator.v:1632" *)
  wire _T_1933;
  (* src = "crypto_accelerator.v:1633" *)
  wire _T_1934;
  (* src = "crypto_accelerator.v:1634" *)
  wire _T_1936;
  (* src = "crypto_accelerator.v:1635" *)
  wire _T_1937;
  (* src = "crypto_accelerator.v:1636" *)
  wire _T_1938;
  (* src = "crypto_accelerator.v:786" *)
  wire _T_195;
  (* src = "crypto_accelerator.v:1638" *)
  wire _T_1963;
  (* src = "crypto_accelerator.v:1639" *)
  wire _T_1965;
  (* src = "crypto_accelerator.v:1640" *)
  wire _T_1967;
  (* src = "crypto_accelerator.v:1641" *)
  wire _T_1969;
  (* src = "crypto_accelerator.v:787" *)
  wire _T_197;
  (* src = "crypto_accelerator.v:1642" *)
  wire _T_1971;
  (* src = "crypto_accelerator.v:1643" *)
  wire _T_1973;
  (* src = "crypto_accelerator.v:1644" *)
  wire _T_1975;
  (* src = "crypto_accelerator.v:1645" *)
  wire _T_1977;
  (* src = "crypto_accelerator.v:1646" *)
  wire _T_1979;
  (* src = "crypto_accelerator.v:1647" *)
  wire _T_1981;
  (* src = "crypto_accelerator.v:1648" *)
  wire _T_1983;
  (* src = "crypto_accelerator.v:1649" *)
  wire _T_1985;
  (* src = "crypto_accelerator.v:1650" *)
  wire _T_1987;
  (* src = "crypto_accelerator.v:1651" *)
  wire _T_1989;
  (* src = "crypto_accelerator.v:788" *)
  wire _T_199;
  (* src = "crypto_accelerator.v:1652" *)
  wire _T_1991;
  (* src = "crypto_accelerator.v:1653" *)
  wire _T_1993;
  (* src = "crypto_accelerator.v:1654" *)
  wire _T_1995;
  (* src = "crypto_accelerator.v:1655" *)
  wire _T_1997;
  (* src = "crypto_accelerator.v:1656" *)
  wire _T_1999;
  (* src = "crypto_accelerator.v:687" *)
  wire _T_2;
  (* src = "crypto_accelerator.v:1657" *)
  wire _T_2001;
  (* src = "crypto_accelerator.v:1658" *)
  wire _T_2003;
  (* src = "crypto_accelerator.v:1659" *)
  wire _T_2005;
  (* src = "crypto_accelerator.v:1660" *)
  wire _T_2007;
  (* src = "crypto_accelerator.v:1661" *)
  wire _T_2009;
  (* src = "crypto_accelerator.v:789" *)
  wire _T_201;
  (* src = "crypto_accelerator.v:1662" *)
  wire _T_2011;
  (* src = "crypto_accelerator.v:1663" *)
  wire _T_2013;
  (* src = "crypto_accelerator.v:1664" *)
  wire _T_2015;
  (* src = "crypto_accelerator.v:1665" *)
  wire _T_2017;
  (* src = "crypto_accelerator.v:1666" *)
  wire _T_2019;
  (* src = "crypto_accelerator.v:1667" *)
  wire _T_2021;
  (* src = "crypto_accelerator.v:1668" *)
  wire _T_2023;
  (* src = "crypto_accelerator.v:1669" *)
  wire _T_2025;
  (* src = "crypto_accelerator.v:1670" *)
  wire _T_2027;
  (* src = "crypto_accelerator.v:1671" *)
  wire _T_2029;
  (* src = "crypto_accelerator.v:790" *)
  wire _T_203;
  (* src = "crypto_accelerator.v:1672" *)
  wire _T_2031;
  (* src = "crypto_accelerator.v:1673" *)
  wire _T_2033;
  (* src = "crypto_accelerator.v:1674" *)
  wire _T_2035;
  (* src = "crypto_accelerator.v:1675" *)
  wire _T_2037;
  (* src = "crypto_accelerator.v:1676" *)
  wire _T_2039;
  (* src = "crypto_accelerator.v:1677" *)
  wire _T_2041;
  (* src = "crypto_accelerator.v:1678" *)
  wire _T_2043;
  (* src = "crypto_accelerator.v:1679" *)
  wire _T_2045;
  (* src = "crypto_accelerator.v:1680" *)
  wire _T_2047;
  (* src = "crypto_accelerator.v:1681" *)
  wire _T_2049;
  (* src = "crypto_accelerator.v:791" *)
  wire _T_205;
  (* src = "crypto_accelerator.v:1682" *)
  wire _T_2051;
  (* src = "crypto_accelerator.v:1683" *)
  wire _T_2053;
  (* src = "crypto_accelerator.v:1684" *)
  wire _T_2055;
  (* src = "crypto_accelerator.v:1685" *)
  wire _T_2057;
  (* src = "crypto_accelerator.v:1686" *)
  wire _T_2059;
  (* src = "crypto_accelerator.v:1687" *)
  wire _T_2061;
  (* src = "crypto_accelerator.v:1688" *)
  wire _T_2063;
  (* src = "crypto_accelerator.v:1689" *)
  wire _T_2065;
  (* src = "crypto_accelerator.v:1690" *)
  wire _T_2067;
  (* src = "crypto_accelerator.v:1691" *)
  wire _T_2069;
  (* src = "crypto_accelerator.v:792" *)
  wire _T_207;
  (* src = "crypto_accelerator.v:1692" *)
  wire _T_2071;
  (* src = "crypto_accelerator.v:1693" *)
  wire _T_2073;
  (* src = "crypto_accelerator.v:1694" *)
  wire _T_2075;
  (* src = "crypto_accelerator.v:1695" *)
  wire _T_2077;
  (* src = "crypto_accelerator.v:1696" *)
  wire _T_2079;
  (* src = "crypto_accelerator.v:1697" *)
  wire _T_2081;
  (* src = "crypto_accelerator.v:1698" *)
  wire _T_2083;
  (* src = "crypto_accelerator.v:1699" *)
  wire _T_2085;
  (* src = "crypto_accelerator.v:1700" *)
  wire _T_2087;
  (* src = "crypto_accelerator.v:1701" *)
  wire _T_2089;
  (* src = "crypto_accelerator.v:793" *)
  wire _T_209;
  (* src = "crypto_accelerator.v:1702" *)
  wire _T_2091;
  (* src = "crypto_accelerator.v:1703" *)
  wire _T_2093;
  (* src = "crypto_accelerator.v:1704" *)
  wire _T_2095;
  (* src = "crypto_accelerator.v:1705" *)
  wire _T_2097;
  (* src = "crypto_accelerator.v:1706" *)
  wire _T_2099;
  (* src = "crypto_accelerator.v:1707" *)
  wire _T_2101;
  (* src = "crypto_accelerator.v:1708" *)
  wire _T_2103;
  (* src = "crypto_accelerator.v:1709" *)
  wire _T_2105;
  (* src = "crypto_accelerator.v:1710" *)
  wire _T_2107;
  (* src = "crypto_accelerator.v:1711" *)
  wire _T_2109;
  (* src = "crypto_accelerator.v:794" *)
  wire _T_211;
  (* src = "crypto_accelerator.v:1712" *)
  wire _T_2111;
  (* src = "crypto_accelerator.v:1713" *)
  wire _T_2113;
  (* src = "crypto_accelerator.v:1714" *)
  wire _T_2115;
  (* src = "crypto_accelerator.v:1715" *)
  wire _T_2117;
  (* src = "crypto_accelerator.v:1716" *)
  wire _T_2119;
  (* src = "crypto_accelerator.v:1717" *)
  wire _T_2121;
  (* src = "crypto_accelerator.v:1718" *)
  wire _T_2123;
  (* src = "crypto_accelerator.v:1719" *)
  wire _T_2125;
  (* src = "crypto_accelerator.v:1720" *)
  wire _T_2127;
  (* src = "crypto_accelerator.v:1721" *)
  wire _T_2129;
  (* src = "crypto_accelerator.v:795" *)
  wire _T_213;
  (* src = "crypto_accelerator.v:1722" *)
  wire _T_2131;
  (* src = "crypto_accelerator.v:1723" *)
  wire _T_2133;
  (* src = "crypto_accelerator.v:1724" *)
  wire _T_2135;
  (* src = "crypto_accelerator.v:1725" *)
  wire _T_2137;
  (* src = "crypto_accelerator.v:1726" *)
  wire _T_2139;
  (* src = "crypto_accelerator.v:1727" *)
  wire _T_2141;
  (* src = "crypto_accelerator.v:1728" *)
  wire _T_2143;
  (* src = "crypto_accelerator.v:1729" *)
  wire _T_2145;
  (* src = "crypto_accelerator.v:1730" *)
  wire _T_2147;
  (* src = "crypto_accelerator.v:1731" *)
  wire _T_2149;
  (* src = "crypto_accelerator.v:796" *)
  wire _T_215;
  (* src = "crypto_accelerator.v:1732" *)
  wire _T_2151;
  (* src = "crypto_accelerator.v:1733" *)
  wire _T_2153;
  (* src = "crypto_accelerator.v:1734" *)
  wire _T_2155;
  (* src = "crypto_accelerator.v:1735" *)
  wire _T_2157;
  (* src = "crypto_accelerator.v:1736" *)
  wire _T_2159;
  (* src = "crypto_accelerator.v:1737" *)
  wire _T_2161;
  (* src = "crypto_accelerator.v:1738" *)
  wire _T_2163;
  (* src = "crypto_accelerator.v:1739" *)
  wire _T_2165;
  (* src = "crypto_accelerator.v:1740" *)
  wire _T_2167;
  (* src = "crypto_accelerator.v:1741" *)
  wire _T_2169;
  (* src = "crypto_accelerator.v:797" *)
  wire _T_217;
  (* src = "crypto_accelerator.v:1742" *)
  wire _T_2171;
  (* src = "crypto_accelerator.v:1743" *)
  wire _T_2173;
  (* src = "crypto_accelerator.v:1744" *)
  wire _T_2175;
  (* src = "crypto_accelerator.v:1745" *)
  wire _T_2177;
  (* src = "crypto_accelerator.v:1746" *)
  wire _T_2179;
  (* src = "crypto_accelerator.v:1747" *)
  wire _T_2180;
  (* src = "crypto_accelerator.v:1748" *)
  wire _T_2181;
  (* src = "crypto_accelerator.v:1749" *)
  wire _T_2182;
  (* src = "crypto_accelerator.v:1750" *)
  wire _T_2184;
  (* src = "crypto_accelerator.v:1751" *)
  wire _T_2185;
  (* src = "crypto_accelerator.v:1752" *)
  wire _T_2186;
  (* src = "crypto_accelerator.v:1753" *)
  wire _T_2188;
  (* src = "crypto_accelerator.v:798" *)
  wire _T_219;
  (* src = "crypto_accelerator.v:1754" *)
  wire _T_2190;
  (* src = "crypto_accelerator.v:1755" *)
  wire _T_2191;
  (* src = "crypto_accelerator.v:1756" *)
  wire _T_2192;
  (* src = "crypto_accelerator.v:1757" *)
  wire _T_2194;
  (* src = "crypto_accelerator.v:1758" *)
  wire _T_2196;
  (* src = "crypto_accelerator.v:1759" *)
  wire _T_2198;
  (* src = "crypto_accelerator.v:1760" *)
  wire _T_2199;
  (* src = "crypto_accelerator.v:1761" *)
  wire _T_2200;
  (* src = "crypto_accelerator.v:1762" *)
  wire _T_2202;
  (* src = "crypto_accelerator.v:1763" *)
  wire _T_2203;
  (* src = "crypto_accelerator.v:1764" *)
  wire _T_2205;
  (* src = "crypto_accelerator.v:1765" *)
  wire _T_2206;
  (* src = "crypto_accelerator.v:1766" *)
  wire _T_2207;
  (* src = "crypto_accelerator.v:799" *)
  wire _T_221;
  (* src = "crypto_accelerator.v:800" *)
  wire _T_223;
  (* src = "crypto_accelerator.v:1768" *)
  wire _T_2233;
  (* src = "crypto_accelerator.v:1769" *)
  wire _T_2235;
  (* src = "crypto_accelerator.v:1770" *)
  wire _T_2237;
  (* src = "crypto_accelerator.v:1771" *)
  wire _T_2239;
  (* src = "crypto_accelerator.v:1772" *)
  wire _T_2241;
  (* src = "crypto_accelerator.v:1773" *)
  wire _T_2243;
  (* src = "crypto_accelerator.v:1774" *)
  wire _T_2245;
  (* src = "crypto_accelerator.v:1775" *)
  wire _T_2247;
  (* src = "crypto_accelerator.v:1776" *)
  wire _T_2249;
  (* src = "crypto_accelerator.v:801" *)
  wire _T_225;
  (* src = "crypto_accelerator.v:1777" *)
  wire _T_2251;
  (* src = "crypto_accelerator.v:1778" *)
  wire _T_2253;
  (* src = "crypto_accelerator.v:1779" *)
  wire _T_2255;
  (* src = "crypto_accelerator.v:1780" *)
  wire _T_2257;
  (* src = "crypto_accelerator.v:1781" *)
  wire _T_2259;
  (* src = "crypto_accelerator.v:1782" *)
  wire _T_2261;
  (* src = "crypto_accelerator.v:1783" *)
  wire _T_2263;
  (* src = "crypto_accelerator.v:1784" *)
  wire _T_2265;
  (* src = "crypto_accelerator.v:1785" *)
  wire _T_2267;
  (* src = "crypto_accelerator.v:1786" *)
  wire _T_2269;
  (* src = "crypto_accelerator.v:802" *)
  wire _T_227;
  (* src = "crypto_accelerator.v:1787" *)
  wire _T_2271;
  (* src = "crypto_accelerator.v:1788" *)
  wire _T_2273;
  (* src = "crypto_accelerator.v:1789" *)
  wire _T_2275;
  (* src = "crypto_accelerator.v:1790" *)
  wire _T_2277;
  (* src = "crypto_accelerator.v:1791" *)
  wire _T_2279;
  (* src = "crypto_accelerator.v:1792" *)
  wire _T_2281;
  (* src = "crypto_accelerator.v:1793" *)
  wire _T_2283;
  (* src = "crypto_accelerator.v:1794" *)
  wire _T_2285;
  (* src = "crypto_accelerator.v:1795" *)
  wire _T_2287;
  (* src = "crypto_accelerator.v:1796" *)
  wire _T_2289;
  (* src = "crypto_accelerator.v:803" *)
  wire _T_229;
  (* src = "crypto_accelerator.v:1797" *)
  wire _T_2291;
  (* src = "crypto_accelerator.v:1798" *)
  wire _T_2293;
  (* src = "crypto_accelerator.v:1799" *)
  wire _T_2295;
  (* src = "crypto_accelerator.v:1800" *)
  wire _T_2297;
  (* src = "crypto_accelerator.v:1801" *)
  wire _T_2299;
  (* src = "crypto_accelerator.v:707" *)
  wire [63:0] _T_23;
  (* src = "crypto_accelerator.v:1802" *)
  wire _T_2301;
  (* src = "crypto_accelerator.v:1803" *)
  wire _T_2303;
  (* src = "crypto_accelerator.v:1804" *)
  wire _T_2305;
  (* src = "crypto_accelerator.v:1805" *)
  wire _T_2307;
  (* src = "crypto_accelerator.v:1806" *)
  wire _T_2309;
  (* src = "crypto_accelerator.v:804" *)
  wire _T_231;
  (* src = "crypto_accelerator.v:1807" *)
  wire _T_2311;
  (* src = "crypto_accelerator.v:1808" *)
  wire _T_2313;
  (* src = "crypto_accelerator.v:1809" *)
  wire _T_2315;
  (* src = "crypto_accelerator.v:1810" *)
  wire _T_2317;
  (* src = "crypto_accelerator.v:1811" *)
  wire _T_2319;
  (* src = "crypto_accelerator.v:1812" *)
  wire _T_2321;
  (* src = "crypto_accelerator.v:1813" *)
  wire _T_2323;
  (* src = "crypto_accelerator.v:1814" *)
  wire _T_2325;
  (* src = "crypto_accelerator.v:1815" *)
  wire _T_2327;
  (* src = "crypto_accelerator.v:1816" *)
  wire _T_2329;
  (* src = "crypto_accelerator.v:805" *)
  wire _T_233;
  (* src = "crypto_accelerator.v:1817" *)
  wire _T_2331;
  (* src = "crypto_accelerator.v:1818" *)
  wire _T_2333;
  (* src = "crypto_accelerator.v:1819" *)
  wire _T_2335;
  (* src = "crypto_accelerator.v:1820" *)
  wire _T_2337;
  (* src = "crypto_accelerator.v:1821" *)
  wire _T_2339;
  (* src = "crypto_accelerator.v:1822" *)
  wire _T_2341;
  (* src = "crypto_accelerator.v:1823" *)
  wire _T_2343;
  (* src = "crypto_accelerator.v:1824" *)
  wire _T_2345;
  (* src = "crypto_accelerator.v:1825" *)
  wire _T_2347;
  (* src = "crypto_accelerator.v:1826" *)
  wire _T_2349;
  (* src = "crypto_accelerator.v:806" *)
  wire _T_235;
  (* src = "crypto_accelerator.v:1827" *)
  wire _T_2351;
  (* src = "crypto_accelerator.v:1828" *)
  wire _T_2353;
  (* src = "crypto_accelerator.v:1829" *)
  wire _T_2355;
  (* src = "crypto_accelerator.v:1830" *)
  wire _T_2357;
  (* src = "crypto_accelerator.v:1831" *)
  wire _T_2359;
  (* src = "crypto_accelerator.v:1832" *)
  wire _T_2361;
  (* src = "crypto_accelerator.v:1833" *)
  wire _T_2363;
  (* src = "crypto_accelerator.v:1834" *)
  wire _T_2365;
  (* src = "crypto_accelerator.v:1835" *)
  wire _T_2367;
  (* src = "crypto_accelerator.v:1836" *)
  wire _T_2369;
  (* src = "crypto_accelerator.v:807" *)
  wire _T_237;
  (* src = "crypto_accelerator.v:1837" *)
  wire _T_2371;
  (* src = "crypto_accelerator.v:1838" *)
  wire _T_2373;
  (* src = "crypto_accelerator.v:1839" *)
  wire _T_2375;
  (* src = "crypto_accelerator.v:1840" *)
  wire _T_2377;
  (* src = "crypto_accelerator.v:1841" *)
  wire _T_2379;
  (* src = "crypto_accelerator.v:1842" *)
  wire _T_2381;
  (* src = "crypto_accelerator.v:1843" *)
  wire _T_2383;
  (* src = "crypto_accelerator.v:1844" *)
  wire _T_2385;
  (* src = "crypto_accelerator.v:1845" *)
  wire _T_2387;
  (* src = "crypto_accelerator.v:1846" *)
  wire _T_2389;
  (* src = "crypto_accelerator.v:808" *)
  wire _T_239;
  (* src = "crypto_accelerator.v:1847" *)
  wire _T_2391;
  (* src = "crypto_accelerator.v:1848" *)
  wire _T_2393;
  (* src = "crypto_accelerator.v:1849" *)
  wire _T_2395;
  (* src = "crypto_accelerator.v:1850" *)
  wire _T_2397;
  (* src = "crypto_accelerator.v:1851" *)
  wire _T_2399;
  (* src = "crypto_accelerator.v:1852" *)
  wire _T_2401;
  (* src = "crypto_accelerator.v:1853" *)
  wire _T_2403;
  (* src = "crypto_accelerator.v:1854" *)
  wire _T_2405;
  (* src = "crypto_accelerator.v:1855" *)
  wire _T_2407;
  (* src = "crypto_accelerator.v:1856" *)
  wire _T_2409;
  (* src = "crypto_accelerator.v:809" *)
  wire _T_241;
  (* src = "crypto_accelerator.v:1857" *)
  wire _T_2411;
  (* src = "crypto_accelerator.v:1858" *)
  wire _T_2413;
  (* src = "crypto_accelerator.v:1859" *)
  wire _T_2415;
  (* src = "crypto_accelerator.v:1860" *)
  wire _T_2417;
  (* src = "crypto_accelerator.v:1861" *)
  wire _T_2419;
  (* src = "crypto_accelerator.v:1862" *)
  wire _T_2421;
  (* src = "crypto_accelerator.v:1863" *)
  wire _T_2423;
  (* src = "crypto_accelerator.v:1864" *)
  wire _T_2425;
  (* src = "crypto_accelerator.v:1865" *)
  wire _T_2427;
  (* src = "crypto_accelerator.v:1866" *)
  wire _T_2429;
  (* src = "crypto_accelerator.v:810" *)
  wire _T_243;
  (* src = "crypto_accelerator.v:1867" *)
  wire _T_2431;
  (* src = "crypto_accelerator.v:1868" *)
  wire _T_2433;
  (* src = "crypto_accelerator.v:1869" *)
  wire _T_2435;
  (* src = "crypto_accelerator.v:1870" *)
  wire _T_2437;
  (* src = "crypto_accelerator.v:1871" *)
  wire _T_2439;
  (* src = "crypto_accelerator.v:1872" *)
  wire _T_2441;
  (* src = "crypto_accelerator.v:1873" *)
  wire _T_2443;
  (* src = "crypto_accelerator.v:1874" *)
  wire _T_2445;
  (* src = "crypto_accelerator.v:1875" *)
  wire _T_2447;
  (* src = "crypto_accelerator.v:1876" *)
  wire _T_2449;
  (* src = "crypto_accelerator.v:811" *)
  wire _T_245;
  (* src = "crypto_accelerator.v:1877" *)
  wire _T_2450;
  (* src = "crypto_accelerator.v:1878" *)
  wire _T_2451;
  (* src = "crypto_accelerator.v:1879" *)
  wire _T_2452;
  (* src = "crypto_accelerator.v:1880" *)
  wire _T_2454;
  (* src = "crypto_accelerator.v:1881" *)
  wire _T_2455;
  (* src = "crypto_accelerator.v:1882" *)
  wire _T_2456;
  (* src = "crypto_accelerator.v:1883" *)
  wire _T_2458;
  (* src = "crypto_accelerator.v:1884" *)
  wire _T_2460;
  (* src = "crypto_accelerator.v:1885" *)
  wire _T_2461;
  (* src = "crypto_accelerator.v:1886" *)
  wire _T_2462;
  (* src = "crypto_accelerator.v:1887" *)
  wire _T_2464;
  (* src = "crypto_accelerator.v:1888" *)
  wire _T_2466;
  (* src = "crypto_accelerator.v:1889" *)
  wire _T_2468;
  (* src = "crypto_accelerator.v:1890" *)
  wire _T_2469;
  (* src = "crypto_accelerator.v:812" *)
  wire _T_247;
  (* src = "crypto_accelerator.v:1891" *)
  wire _T_2470;
  (* src = "crypto_accelerator.v:1892" *)
  wire _T_2472;
  (* src = "crypto_accelerator.v:1893" *)
  wire _T_2473;
  (* src = "crypto_accelerator.v:1894" *)
  wire _T_2475;
  (* src = "crypto_accelerator.v:1895" *)
  wire _T_2476;
  (* src = "crypto_accelerator.v:1896" *)
  wire _T_2477;
  (* src = "crypto_accelerator.v:813" *)
  wire _T_249;
  (* src = "crypto_accelerator.v:708" *)
  wire [127:0] _T_25;
  (* src = "crypto_accelerator.v:1898" *)
  wire _T_2502;
  (* src = "crypto_accelerator.v:1899" *)
  wire _T_2504;
  (* src = "crypto_accelerator.v:1900" *)
  wire _T_2506;
  (* src = "crypto_accelerator.v:1901" *)
  wire _T_2508;
  (* src = "crypto_accelerator.v:814" *)
  wire _T_251;
  (* src = "crypto_accelerator.v:1902" *)
  wire _T_2510;
  (* src = "crypto_accelerator.v:1903" *)
  wire _T_2512;
  (* src = "crypto_accelerator.v:1904" *)
  wire _T_2514;
  (* src = "crypto_accelerator.v:1905" *)
  wire _T_2516;
  (* src = "crypto_accelerator.v:1906" *)
  wire _T_2518;
  (* src = "crypto_accelerator.v:1907" *)
  wire _T_2520;
  (* src = "crypto_accelerator.v:1908" *)
  wire _T_2522;
  (* src = "crypto_accelerator.v:1909" *)
  wire _T_2524;
  (* src = "crypto_accelerator.v:1910" *)
  wire _T_2526;
  (* src = "crypto_accelerator.v:1911" *)
  wire _T_2528;
  (* src = "crypto_accelerator.v:815" *)
  wire _T_253;
  (* src = "crypto_accelerator.v:1912" *)
  wire _T_2530;
  (* src = "crypto_accelerator.v:1913" *)
  wire _T_2532;
  (* src = "crypto_accelerator.v:1914" *)
  wire _T_2534;
  (* src = "crypto_accelerator.v:1915" *)
  wire _T_2536;
  (* src = "crypto_accelerator.v:1916" *)
  wire _T_2538;
  (* src = "crypto_accelerator.v:1917" *)
  wire _T_2540;
  (* src = "crypto_accelerator.v:1918" *)
  wire _T_2542;
  (* src = "crypto_accelerator.v:1919" *)
  wire _T_2544;
  (* src = "crypto_accelerator.v:1920" *)
  wire _T_2546;
  (* src = "crypto_accelerator.v:1921" *)
  wire _T_2548;
  (* src = "crypto_accelerator.v:816" *)
  wire _T_255;
  (* src = "crypto_accelerator.v:1922" *)
  wire _T_2550;
  (* src = "crypto_accelerator.v:1923" *)
  wire _T_2552;
  (* src = "crypto_accelerator.v:1924" *)
  wire _T_2554;
  (* src = "crypto_accelerator.v:1925" *)
  wire _T_2556;
  (* src = "crypto_accelerator.v:1926" *)
  wire _T_2558;
  (* src = "crypto_accelerator.v:1927" *)
  wire _T_2560;
  (* src = "crypto_accelerator.v:1928" *)
  wire _T_2562;
  (* src = "crypto_accelerator.v:1929" *)
  wire _T_2564;
  (* src = "crypto_accelerator.v:1930" *)
  wire _T_2566;
  (* src = "crypto_accelerator.v:1931" *)
  wire _T_2568;
  (* src = "crypto_accelerator.v:817" *)
  wire _T_257;
  (* src = "crypto_accelerator.v:1932" *)
  wire _T_2570;
  (* src = "crypto_accelerator.v:1933" *)
  wire _T_2572;
  (* src = "crypto_accelerator.v:1934" *)
  wire _T_2574;
  (* src = "crypto_accelerator.v:1935" *)
  wire _T_2576;
  (* src = "crypto_accelerator.v:1936" *)
  wire _T_2578;
  (* src = "crypto_accelerator.v:1937" *)
  wire _T_2580;
  (* src = "crypto_accelerator.v:1938" *)
  wire _T_2582;
  (* src = "crypto_accelerator.v:1939" *)
  wire _T_2584;
  (* src = "crypto_accelerator.v:1940" *)
  wire _T_2586;
  (* src = "crypto_accelerator.v:1941" *)
  wire _T_2588;
  (* src = "crypto_accelerator.v:818" *)
  wire _T_259;
  (* src = "crypto_accelerator.v:1942" *)
  wire _T_2590;
  (* src = "crypto_accelerator.v:1943" *)
  wire _T_2592;
  (* src = "crypto_accelerator.v:1944" *)
  wire _T_2594;
  (* src = "crypto_accelerator.v:1945" *)
  wire _T_2596;
  (* src = "crypto_accelerator.v:1946" *)
  wire _T_2598;
  (* src = "crypto_accelerator.v:1947" *)
  wire _T_2600;
  (* src = "crypto_accelerator.v:1948" *)
  wire _T_2602;
  (* src = "crypto_accelerator.v:1949" *)
  wire _T_2604;
  (* src = "crypto_accelerator.v:1950" *)
  wire _T_2606;
  (* src = "crypto_accelerator.v:1951" *)
  wire _T_2608;
  (* src = "crypto_accelerator.v:819" *)
  wire _T_261;
  (* src = "crypto_accelerator.v:1952" *)
  wire _T_2610;
  (* src = "crypto_accelerator.v:1953" *)
  wire _T_2612;
  (* src = "crypto_accelerator.v:1954" *)
  wire _T_2614;
  (* src = "crypto_accelerator.v:1955" *)
  wire _T_2616;
  (* src = "crypto_accelerator.v:1956" *)
  wire _T_2618;
  (* src = "crypto_accelerator.v:1957" *)
  wire _T_2620;
  (* src = "crypto_accelerator.v:1958" *)
  wire _T_2622;
  (* src = "crypto_accelerator.v:1959" *)
  wire _T_2624;
  (* src = "crypto_accelerator.v:1960" *)
  wire _T_2626;
  (* src = "crypto_accelerator.v:1961" *)
  wire _T_2628;
  (* src = "crypto_accelerator.v:820" *)
  wire _T_263;
  (* src = "crypto_accelerator.v:1962" *)
  wire _T_2630;
  (* src = "crypto_accelerator.v:1963" *)
  wire _T_2632;
  (* src = "crypto_accelerator.v:1964" *)
  wire _T_2634;
  (* src = "crypto_accelerator.v:1965" *)
  wire _T_2636;
  (* src = "crypto_accelerator.v:1966" *)
  wire _T_2638;
  (* src = "crypto_accelerator.v:1967" *)
  wire _T_2640;
  (* src = "crypto_accelerator.v:1968" *)
  wire _T_2642;
  (* src = "crypto_accelerator.v:1969" *)
  wire _T_2644;
  (* src = "crypto_accelerator.v:1970" *)
  wire _T_2646;
  (* src = "crypto_accelerator.v:1971" *)
  wire _T_2648;
  (* src = "crypto_accelerator.v:821" *)
  wire _T_265;
  (* src = "crypto_accelerator.v:1972" *)
  wire _T_2650;
  (* src = "crypto_accelerator.v:1973" *)
  wire _T_2652;
  (* src = "crypto_accelerator.v:1974" *)
  wire _T_2654;
  (* src = "crypto_accelerator.v:1975" *)
  wire _T_2656;
  (* src = "crypto_accelerator.v:1976" *)
  wire _T_2658;
  (* src = "crypto_accelerator.v:1977" *)
  wire _T_2660;
  (* src = "crypto_accelerator.v:1978" *)
  wire _T_2662;
  (* src = "crypto_accelerator.v:1979" *)
  wire _T_2664;
  (* src = "crypto_accelerator.v:1980" *)
  wire _T_2666;
  (* src = "crypto_accelerator.v:1981" *)
  wire _T_2668;
  (* src = "crypto_accelerator.v:822" *)
  wire _T_267;
  (* src = "crypto_accelerator.v:1982" *)
  wire _T_2670;
  (* src = "crypto_accelerator.v:1983" *)
  wire _T_2672;
  (* src = "crypto_accelerator.v:1984" *)
  wire _T_2674;
  (* src = "crypto_accelerator.v:1985" *)
  wire _T_2676;
  (* src = "crypto_accelerator.v:1986" *)
  wire _T_2678;
  (* src = "crypto_accelerator.v:1987" *)
  wire _T_2680;
  (* src = "crypto_accelerator.v:1988" *)
  wire _T_2682;
  (* src = "crypto_accelerator.v:1989" *)
  wire _T_2684;
  (* src = "crypto_accelerator.v:1990" *)
  wire _T_2686;
  (* src = "crypto_accelerator.v:1991" *)
  wire _T_2688;
  (* src = "crypto_accelerator.v:823" *)
  wire _T_269;
  (* src = "crypto_accelerator.v:1992" *)
  wire _T_2690;
  (* src = "crypto_accelerator.v:1993" *)
  wire _T_2692;
  (* src = "crypto_accelerator.v:1994" *)
  wire _T_2694;
  (* src = "crypto_accelerator.v:1995" *)
  wire _T_2696;
  (* src = "crypto_accelerator.v:1996" *)
  wire _T_2698;
  (* src = "crypto_accelerator.v:1997" *)
  wire _T_2700;
  (* src = "crypto_accelerator.v:1998" *)
  wire _T_2702;
  (* src = "crypto_accelerator.v:1999" *)
  wire _T_2704;
  (* src = "crypto_accelerator.v:2000" *)
  wire _T_2706;
  (* src = "crypto_accelerator.v:2001" *)
  wire _T_2708;
  (* src = "crypto_accelerator.v:824" *)
  wire _T_271;
  (* src = "crypto_accelerator.v:2002" *)
  wire _T_2710;
  (* src = "crypto_accelerator.v:2003" *)
  wire _T_2712;
  (* src = "crypto_accelerator.v:2004" *)
  wire _T_2714;
  (* src = "crypto_accelerator.v:2005" *)
  wire _T_2716;
  (* src = "crypto_accelerator.v:2006" *)
  wire _T_2718;
  (* src = "crypto_accelerator.v:2007" *)
  wire _T_2719;
  (* src = "crypto_accelerator.v:2008" *)
  wire _T_2720;
  (* src = "crypto_accelerator.v:2009" *)
  wire _T_2721;
  (* src = "crypto_accelerator.v:2010" *)
  wire _T_2723;
  (* src = "crypto_accelerator.v:2011" *)
  wire _T_2724;
  (* src = "crypto_accelerator.v:2012" *)
  wire _T_2725;
  (* src = "crypto_accelerator.v:2013" *)
  wire _T_2727;
  (* src = "crypto_accelerator.v:2014" *)
  wire _T_2729;
  (* src = "crypto_accelerator.v:825" *)
  wire _T_273;
  (* src = "crypto_accelerator.v:2015" *)
  wire _T_2730;
  (* src = "crypto_accelerator.v:2016" *)
  wire _T_2731;
  (* src = "crypto_accelerator.v:2017" *)
  wire _T_2733;
  (* src = "crypto_accelerator.v:2018" *)
  wire _T_2735;
  (* src = "crypto_accelerator.v:2019" *)
  wire _T_2737;
  (* src = "crypto_accelerator.v:2020" *)
  wire _T_2738;
  (* src = "crypto_accelerator.v:2021" *)
  wire _T_2739;
  (* src = "crypto_accelerator.v:2022" *)
  wire _T_2741;
  (* src = "crypto_accelerator.v:2023" *)
  wire _T_2742;
  (* src = "crypto_accelerator.v:2024" *)
  wire _T_2744;
  (* src = "crypto_accelerator.v:2025" *)
  wire _T_2745;
  (* src = "crypto_accelerator.v:2026" *)
  wire _T_2746;
  (* src = "crypto_accelerator.v:826" *)
  wire _T_275;
  (* src = "crypto_accelerator.v:827" *)
  wire _T_277;
  (* src = "crypto_accelerator.v:2028" *)
  wire _T_2771;
  (* src = "crypto_accelerator.v:2029" *)
  wire _T_2773;
  (* src = "crypto_accelerator.v:2030" *)
  wire _T_2775;
  (* src = "crypto_accelerator.v:2031" *)
  wire _T_2777;
  (* src = "crypto_accelerator.v:2032" *)
  wire _T_2779;
  (* src = "crypto_accelerator.v:2033" *)
  wire _T_2781;
  (* src = "crypto_accelerator.v:2034" *)
  wire _T_2783;
  (* src = "crypto_accelerator.v:2035" *)
  wire _T_2785;
  (* src = "crypto_accelerator.v:2036" *)
  wire _T_2787;
  (* src = "crypto_accelerator.v:2037" *)
  wire _T_2789;
  (* src = "crypto_accelerator.v:828" *)
  wire _T_279;
  (* src = "crypto_accelerator.v:2038" *)
  wire _T_2791;
  (* src = "crypto_accelerator.v:2039" *)
  wire _T_2793;
  (* src = "crypto_accelerator.v:2040" *)
  wire _T_2795;
  (* src = "crypto_accelerator.v:2041" *)
  wire _T_2797;
  (* src = "crypto_accelerator.v:2042" *)
  wire _T_2799;
  (* src = "crypto_accelerator.v:2043" *)
  wire _T_2801;
  (* src = "crypto_accelerator.v:2044" *)
  wire _T_2803;
  (* src = "crypto_accelerator.v:2045" *)
  wire _T_2805;
  (* src = "crypto_accelerator.v:2046" *)
  wire _T_2807;
  (* src = "crypto_accelerator.v:2047" *)
  wire _T_2809;
  (* src = "crypto_accelerator.v:829" *)
  wire _T_281;
  (* src = "crypto_accelerator.v:2048" *)
  wire _T_2811;
  (* src = "crypto_accelerator.v:2049" *)
  wire _T_2813;
  (* src = "crypto_accelerator.v:2050" *)
  wire _T_2815;
  (* src = "crypto_accelerator.v:2051" *)
  wire _T_2817;
  (* src = "crypto_accelerator.v:2052" *)
  wire _T_2819;
  (* src = "crypto_accelerator.v:2053" *)
  wire _T_2821;
  (* src = "crypto_accelerator.v:2054" *)
  wire _T_2823;
  (* src = "crypto_accelerator.v:2055" *)
  wire _T_2825;
  (* src = "crypto_accelerator.v:2056" *)
  wire _T_2827;
  (* src = "crypto_accelerator.v:2057" *)
  wire _T_2829;
  (* src = "crypto_accelerator.v:830" *)
  wire _T_283;
  (* src = "crypto_accelerator.v:2058" *)
  wire _T_2831;
  (* src = "crypto_accelerator.v:2059" *)
  wire _T_2833;
  (* src = "crypto_accelerator.v:2060" *)
  wire _T_2835;
  (* src = "crypto_accelerator.v:2061" *)
  wire _T_2837;
  (* src = "crypto_accelerator.v:2062" *)
  wire _T_2839;
  (* src = "crypto_accelerator.v:2063" *)
  wire _T_2841;
  (* src = "crypto_accelerator.v:2064" *)
  wire _T_2843;
  (* src = "crypto_accelerator.v:2065" *)
  wire _T_2845;
  (* src = "crypto_accelerator.v:2066" *)
  wire _T_2847;
  (* src = "crypto_accelerator.v:2067" *)
  wire _T_2849;
  (* src = "crypto_accelerator.v:831" *)
  wire _T_285;
  (* src = "crypto_accelerator.v:2068" *)
  wire _T_2851;
  (* src = "crypto_accelerator.v:2069" *)
  wire _T_2853;
  (* src = "crypto_accelerator.v:2070" *)
  wire _T_2855;
  (* src = "crypto_accelerator.v:2071" *)
  wire _T_2857;
  (* src = "crypto_accelerator.v:2072" *)
  wire _T_2859;
  (* src = "crypto_accelerator.v:2073" *)
  wire _T_2861;
  (* src = "crypto_accelerator.v:2074" *)
  wire _T_2863;
  (* src = "crypto_accelerator.v:2075" *)
  wire _T_2865;
  (* src = "crypto_accelerator.v:2076" *)
  wire _T_2867;
  (* src = "crypto_accelerator.v:2077" *)
  wire _T_2869;
  (* src = "crypto_accelerator.v:832" *)
  wire _T_287;
  (* src = "crypto_accelerator.v:2078" *)
  wire _T_2871;
  (* src = "crypto_accelerator.v:2079" *)
  wire _T_2873;
  (* src = "crypto_accelerator.v:2080" *)
  wire _T_2875;
  (* src = "crypto_accelerator.v:2081" *)
  wire _T_2877;
  (* src = "crypto_accelerator.v:2082" *)
  wire _T_2879;
  (* src = "crypto_accelerator.v:2083" *)
  wire _T_2881;
  (* src = "crypto_accelerator.v:2084" *)
  wire _T_2883;
  (* src = "crypto_accelerator.v:2085" *)
  wire _T_2885;
  (* src = "crypto_accelerator.v:2086" *)
  wire _T_2887;
  (* src = "crypto_accelerator.v:2087" *)
  wire _T_2889;
  (* src = "crypto_accelerator.v:833" *)
  wire _T_289;
  (* src = "crypto_accelerator.v:2088" *)
  wire _T_2891;
  (* src = "crypto_accelerator.v:2089" *)
  wire _T_2893;
  (* src = "crypto_accelerator.v:2090" *)
  wire _T_2895;
  (* src = "crypto_accelerator.v:2091" *)
  wire _T_2897;
  (* src = "crypto_accelerator.v:2092" *)
  wire _T_2899;
  (* src = "crypto_accelerator.v:2093" *)
  wire _T_2901;
  (* src = "crypto_accelerator.v:2094" *)
  wire _T_2903;
  (* src = "crypto_accelerator.v:2095" *)
  wire _T_2905;
  (* src = "crypto_accelerator.v:2096" *)
  wire _T_2907;
  (* src = "crypto_accelerator.v:2097" *)
  wire _T_2909;
  (* src = "crypto_accelerator.v:834" *)
  wire _T_291;
  (* src = "crypto_accelerator.v:2098" *)
  wire _T_2911;
  (* src = "crypto_accelerator.v:2099" *)
  wire _T_2913;
  (* src = "crypto_accelerator.v:2100" *)
  wire _T_2915;
  (* src = "crypto_accelerator.v:2101" *)
  wire _T_2917;
  (* src = "crypto_accelerator.v:2102" *)
  wire _T_2919;
  (* src = "crypto_accelerator.v:2103" *)
  wire _T_2921;
  (* src = "crypto_accelerator.v:2104" *)
  wire _T_2923;
  (* src = "crypto_accelerator.v:2105" *)
  wire _T_2925;
  (* src = "crypto_accelerator.v:2106" *)
  wire _T_2927;
  (* src = "crypto_accelerator.v:2107" *)
  wire _T_2929;
  (* src = "crypto_accelerator.v:835" *)
  wire _T_293;
  (* src = "crypto_accelerator.v:2108" *)
  wire _T_2931;
  (* src = "crypto_accelerator.v:2109" *)
  wire _T_2933;
  (* src = "crypto_accelerator.v:2110" *)
  wire _T_2935;
  (* src = "crypto_accelerator.v:2111" *)
  wire _T_2937;
  (* src = "crypto_accelerator.v:2112" *)
  wire _T_2939;
  (* src = "crypto_accelerator.v:2113" *)
  wire _T_2941;
  (* src = "crypto_accelerator.v:2114" *)
  wire _T_2943;
  (* src = "crypto_accelerator.v:2115" *)
  wire _T_2945;
  (* src = "crypto_accelerator.v:2116" *)
  wire _T_2947;
  (* src = "crypto_accelerator.v:2117" *)
  wire _T_2949;
  (* src = "crypto_accelerator.v:836" *)
  wire _T_295;
  (* src = "crypto_accelerator.v:2118" *)
  wire _T_2951;
  (* src = "crypto_accelerator.v:2119" *)
  wire _T_2953;
  (* src = "crypto_accelerator.v:2120" *)
  wire _T_2955;
  (* src = "crypto_accelerator.v:2121" *)
  wire _T_2957;
  (* src = "crypto_accelerator.v:2122" *)
  wire _T_2959;
  (* src = "crypto_accelerator.v:837" *)
  wire _T_296;
  (* src = "crypto_accelerator.v:2123" *)
  wire _T_2961;
  (* src = "crypto_accelerator.v:2124" *)
  wire _T_2963;
  (* src = "crypto_accelerator.v:2125" *)
  wire _T_2965;
  (* src = "crypto_accelerator.v:2126" *)
  wire _T_2967;
  (* src = "crypto_accelerator.v:2127" *)
  wire _T_2969;
  (* src = "crypto_accelerator.v:838" *)
  wire _T_297;
  (* src = "crypto_accelerator.v:2128" *)
  wire _T_2971;
  (* src = "crypto_accelerator.v:2129" *)
  wire _T_2973;
  (* src = "crypto_accelerator.v:2130" *)
  wire _T_2975;
  (* src = "crypto_accelerator.v:2131" *)
  wire _T_2977;
  (* src = "crypto_accelerator.v:2132" *)
  wire _T_2979;
  (* src = "crypto_accelerator.v:839" *)
  wire _T_298;
  (* src = "crypto_accelerator.v:2133" *)
  wire _T_2981;
  (* src = "crypto_accelerator.v:2134" *)
  wire _T_2983;
  (* src = "crypto_accelerator.v:2135" *)
  wire _T_2985;
  (* src = "crypto_accelerator.v:2136" *)
  wire _T_2987;
  (* src = "crypto_accelerator.v:2137" *)
  wire _T_2988;
  (* src = "crypto_accelerator.v:2138" *)
  wire _T_2989;
  (* src = "crypto_accelerator.v:2139" *)
  wire _T_2990;
  (* src = "crypto_accelerator.v:2140" *)
  wire _T_2992;
  (* src = "crypto_accelerator.v:2141" *)
  wire _T_2993;
  (* src = "crypto_accelerator.v:2142" *)
  wire _T_2994;
  (* src = "crypto_accelerator.v:2143" *)
  wire _T_2996;
  (* src = "crypto_accelerator.v:2144" *)
  wire _T_2998;
  (* src = "crypto_accelerator.v:2145" *)
  wire _T_2999;
  (* src = "crypto_accelerator.v:688" *)
  wire _T_3;
  (* src = "crypto_accelerator.v:840" *)
  wire _T_300;
  (* src = "crypto_accelerator.v:2146" *)
  wire _T_3000;
  (* src = "crypto_accelerator.v:2147" *)
  wire _T_3002;
  (* src = "crypto_accelerator.v:2148" *)
  wire _T_3004;
  (* src = "crypto_accelerator.v:2149" *)
  wire _T_3006;
  (* src = "crypto_accelerator.v:2150" *)
  wire _T_3007;
  (* src = "crypto_accelerator.v:2151" *)
  wire _T_3008;
  (* src = "crypto_accelerator.v:841" *)
  wire _T_301;
  (* src = "crypto_accelerator.v:2152" *)
  wire _T_3010;
  (* src = "crypto_accelerator.v:2153" *)
  wire _T_3011;
  (* src = "crypto_accelerator.v:2154" *)
  wire _T_3013;
  (* src = "crypto_accelerator.v:2155" *)
  wire _T_3014;
  (* src = "crypto_accelerator.v:2156" *)
  wire _T_3015;
  (* src = "crypto_accelerator.v:842" *)
  wire _T_302;
  (* src = "crypto_accelerator.v:843" *)
  wire _T_304;
  (* src = "crypto_accelerator.v:2158" *)
  wire _T_3040;
  (* src = "crypto_accelerator.v:2159" *)
  wire _T_3042;
  (* src = "crypto_accelerator.v:2160" *)
  wire _T_3044;
  (* src = "crypto_accelerator.v:2161" *)
  wire _T_3046;
  (* src = "crypto_accelerator.v:2162" *)
  wire _T_3048;
  (* src = "crypto_accelerator.v:2163" *)
  wire _T_3050;
  (* src = "crypto_accelerator.v:2164" *)
  wire _T_3052;
  (* src = "crypto_accelerator.v:2165" *)
  wire _T_3054;
  (* src = "crypto_accelerator.v:2166" *)
  wire _T_3056;
  (* src = "crypto_accelerator.v:2167" *)
  wire _T_3058;
  (* src = "crypto_accelerator.v:844" *)
  wire _T_306;
  (* src = "crypto_accelerator.v:2168" *)
  wire _T_3060;
  (* src = "crypto_accelerator.v:2169" *)
  wire _T_3062;
  (* src = "crypto_accelerator.v:2170" *)
  wire _T_3064;
  (* src = "crypto_accelerator.v:2171" *)
  wire _T_3066;
  (* src = "crypto_accelerator.v:2172" *)
  wire _T_3068;
  (* src = "crypto_accelerator.v:845" *)
  wire _T_307;
  (* src = "crypto_accelerator.v:2173" *)
  wire _T_3070;
  (* src = "crypto_accelerator.v:2174" *)
  wire _T_3072;
  (* src = "crypto_accelerator.v:2175" *)
  wire _T_3074;
  (* src = "crypto_accelerator.v:2176" *)
  wire _T_3076;
  (* src = "crypto_accelerator.v:2177" *)
  wire _T_3078;
  (* src = "crypto_accelerator.v:846" *)
  wire _T_308;
  (* src = "crypto_accelerator.v:2178" *)
  wire _T_3080;
  (* src = "crypto_accelerator.v:2179" *)
  wire _T_3082;
  (* src = "crypto_accelerator.v:2180" *)
  wire _T_3084;
  (* src = "crypto_accelerator.v:2181" *)
  wire _T_3086;
  (* src = "crypto_accelerator.v:2182" *)
  wire _T_3088;
  (* src = "crypto_accelerator.v:2183" *)
  wire _T_3090;
  (* src = "crypto_accelerator.v:2184" *)
  wire _T_3092;
  (* src = "crypto_accelerator.v:2185" *)
  wire _T_3094;
  (* src = "crypto_accelerator.v:2186" *)
  wire _T_3096;
  (* src = "crypto_accelerator.v:2187" *)
  wire _T_3098;
  (* src = "crypto_accelerator.v:847" *)
  wire _T_310;
  (* src = "crypto_accelerator.v:2188" *)
  wire _T_3100;
  (* src = "crypto_accelerator.v:2189" *)
  wire _T_3102;
  (* src = "crypto_accelerator.v:2190" *)
  wire _T_3104;
  (* src = "crypto_accelerator.v:2191" *)
  wire _T_3106;
  (* src = "crypto_accelerator.v:2192" *)
  wire _T_3108;
  (* src = "crypto_accelerator.v:2193" *)
  wire _T_3110;
  (* src = "crypto_accelerator.v:2194" *)
  wire _T_3112;
  (* src = "crypto_accelerator.v:2195" *)
  wire _T_3114;
  (* src = "crypto_accelerator.v:2196" *)
  wire _T_3116;
  (* src = "crypto_accelerator.v:2197" *)
  wire _T_3118;
  (* src = "crypto_accelerator.v:848" *)
  wire _T_312;
  (* src = "crypto_accelerator.v:2198" *)
  wire _T_3120;
  (* src = "crypto_accelerator.v:2199" *)
  wire _T_3122;
  (* src = "crypto_accelerator.v:2200" *)
  wire _T_3124;
  (* src = "crypto_accelerator.v:2201" *)
  wire _T_3126;
  (* src = "crypto_accelerator.v:2202" *)
  wire _T_3128;
  (* src = "crypto_accelerator.v:2203" *)
  wire _T_3130;
  (* src = "crypto_accelerator.v:2204" *)
  wire _T_3132;
  (* src = "crypto_accelerator.v:2205" *)
  wire _T_3134;
  (* src = "crypto_accelerator.v:2206" *)
  wire _T_3136;
  (* src = "crypto_accelerator.v:2207" *)
  wire _T_3138;
  (* src = "crypto_accelerator.v:849" *)
  wire _T_314;
  (* src = "crypto_accelerator.v:2208" *)
  wire _T_3140;
  (* src = "crypto_accelerator.v:2209" *)
  wire _T_3142;
  (* src = "crypto_accelerator.v:2210" *)
  wire _T_3144;
  (* src = "crypto_accelerator.v:2211" *)
  wire _T_3146;
  (* src = "crypto_accelerator.v:2212" *)
  wire _T_3148;
  (* src = "crypto_accelerator.v:850" *)
  wire _T_315;
  (* src = "crypto_accelerator.v:2213" *)
  wire _T_3150;
  (* src = "crypto_accelerator.v:2214" *)
  wire _T_3152;
  (* src = "crypto_accelerator.v:2215" *)
  wire _T_3154;
  (* src = "crypto_accelerator.v:2216" *)
  wire _T_3156;
  (* src = "crypto_accelerator.v:2217" *)
  wire _T_3158;
  (* src = "crypto_accelerator.v:851" *)
  wire _T_316;
  (* src = "crypto_accelerator.v:2218" *)
  wire _T_3160;
  (* src = "crypto_accelerator.v:2219" *)
  wire _T_3162;
  (* src = "crypto_accelerator.v:2220" *)
  wire _T_3164;
  (* src = "crypto_accelerator.v:2221" *)
  wire _T_3166;
  (* src = "crypto_accelerator.v:2222" *)
  wire _T_3168;
  (* src = "crypto_accelerator.v:2223" *)
  wire _T_3170;
  (* src = "crypto_accelerator.v:2224" *)
  wire _T_3172;
  (* src = "crypto_accelerator.v:2225" *)
  wire _T_3174;
  (* src = "crypto_accelerator.v:2226" *)
  wire _T_3176;
  (* src = "crypto_accelerator.v:2227" *)
  wire _T_3178;
  (* src = "crypto_accelerator.v:852" *)
  wire _T_318;
  (* src = "crypto_accelerator.v:2228" *)
  wire _T_3180;
  (* src = "crypto_accelerator.v:2229" *)
  wire _T_3182;
  (* src = "crypto_accelerator.v:2230" *)
  wire _T_3184;
  (* src = "crypto_accelerator.v:2231" *)
  wire _T_3186;
  (* src = "crypto_accelerator.v:2232" *)
  wire _T_3188;
  (* src = "crypto_accelerator.v:853" *)
  wire _T_319;
  (* src = "crypto_accelerator.v:2233" *)
  wire _T_3190;
  (* src = "crypto_accelerator.v:2234" *)
  wire _T_3192;
  (* src = "crypto_accelerator.v:2235" *)
  wire _T_3194;
  (* src = "crypto_accelerator.v:2236" *)
  wire _T_3196;
  (* src = "crypto_accelerator.v:2237" *)
  wire _T_3198;
  (* src = "crypto_accelerator.v:709" *)
  wire [63:0] _T_32;
  (* src = "crypto_accelerator.v:2238" *)
  wire _T_3200;
  (* src = "crypto_accelerator.v:2239" *)
  wire _T_3202;
  (* src = "crypto_accelerator.v:2240" *)
  wire _T_3204;
  (* src = "crypto_accelerator.v:2241" *)
  wire _T_3206;
  (* src = "crypto_accelerator.v:2242" *)
  wire _T_3208;
  (* src = "crypto_accelerator.v:854" *)
  wire _T_321;
  (* src = "crypto_accelerator.v:2243" *)
  wire _T_3210;
  (* src = "crypto_accelerator.v:2244" *)
  wire _T_3212;
  (* src = "crypto_accelerator.v:2245" *)
  wire _T_3214;
  (* src = "crypto_accelerator.v:2246" *)
  wire _T_3216;
  (* src = "crypto_accelerator.v:2247" *)
  wire _T_3218;
  (* src = "crypto_accelerator.v:855" *)
  wire _T_322;
  (* src = "crypto_accelerator.v:2248" *)
  wire _T_3220;
  (* src = "crypto_accelerator.v:2249" *)
  wire _T_3222;
  (* src = "crypto_accelerator.v:2250" *)
  wire _T_3224;
  (* src = "crypto_accelerator.v:2251" *)
  wire _T_3226;
  (* src = "crypto_accelerator.v:2252" *)
  wire _T_3228;
  (* src = "crypto_accelerator.v:856" *)
  wire _T_323;
  (* src = "crypto_accelerator.v:2253" *)
  wire _T_3230;
  (* src = "crypto_accelerator.v:2254" *)
  wire _T_3232;
  (* src = "crypto_accelerator.v:2255" *)
  wire _T_3234;
  (* src = "crypto_accelerator.v:2256" *)
  wire _T_3236;
  (* src = "crypto_accelerator.v:2257" *)
  wire _T_3238;
  (* src = "crypto_accelerator.v:2258" *)
  wire _T_3240;
  (* src = "crypto_accelerator.v:2259" *)
  wire _T_3242;
  (* src = "crypto_accelerator.v:2260" *)
  wire _T_3244;
  (* src = "crypto_accelerator.v:2261" *)
  wire _T_3246;
  (* src = "crypto_accelerator.v:2262" *)
  wire _T_3248;
  (* src = "crypto_accelerator.v:2263" *)
  wire _T_3250;
  (* src = "crypto_accelerator.v:2264" *)
  wire _T_3252;
  (* src = "crypto_accelerator.v:2265" *)
  wire _T_3254;
  (* src = "crypto_accelerator.v:2266" *)
  wire _T_3256;
  (* src = "crypto_accelerator.v:2267" *)
  wire _T_3257;
  (* src = "crypto_accelerator.v:2268" *)
  wire _T_3258;
  (* src = "crypto_accelerator.v:2269" *)
  wire _T_3259;
  (* src = "crypto_accelerator.v:2270" *)
  wire _T_3261;
  (* src = "crypto_accelerator.v:2271" *)
  wire _T_3262;
  (* src = "crypto_accelerator.v:2272" *)
  wire _T_3263;
  (* src = "crypto_accelerator.v:2273" *)
  wire _T_3265;
  (* src = "crypto_accelerator.v:2274" *)
  wire _T_3267;
  (* src = "crypto_accelerator.v:2275" *)
  wire _T_3268;
  (* src = "crypto_accelerator.v:2276" *)
  wire _T_3269;
  (* src = "crypto_accelerator.v:2277" *)
  wire _T_3271;
  (* src = "crypto_accelerator.v:2278" *)
  wire _T_3273;
  (* src = "crypto_accelerator.v:2279" *)
  wire _T_3275;
  (* src = "crypto_accelerator.v:2280" *)
  wire _T_3276;
  (* src = "crypto_accelerator.v:2281" *)
  wire _T_3277;
  (* src = "crypto_accelerator.v:2282" *)
  wire _T_3279;
  (* src = "crypto_accelerator.v:2283" *)
  wire _T_3280;
  (* src = "crypto_accelerator.v:2284" *)
  wire _T_3282;
  (* src = "crypto_accelerator.v:2285" *)
  wire _T_3283;
  (* src = "crypto_accelerator.v:2286" *)
  wire _T_3284;
  (* src = "crypto_accelerator.v:2288" *)
  wire _T_3310;
  (* src = "crypto_accelerator.v:2289" *)
  wire _T_3312;
  (* src = "crypto_accelerator.v:2290" *)
  wire _T_3314;
  (* src = "crypto_accelerator.v:2291" *)
  wire _T_3316;
  (* src = "crypto_accelerator.v:2292" *)
  wire _T_3318;
  (* src = "crypto_accelerator.v:2293" *)
  wire _T_3320;
  (* src = "crypto_accelerator.v:2294" *)
  wire _T_3322;
  (* src = "crypto_accelerator.v:2295" *)
  wire _T_3324;
  (* src = "crypto_accelerator.v:2296" *)
  wire _T_3326;
  (* src = "crypto_accelerator.v:2297" *)
  wire _T_3328;
  (* src = "crypto_accelerator.v:2298" *)
  wire _T_3330;
  (* src = "crypto_accelerator.v:2299" *)
  wire _T_3332;
  (* src = "crypto_accelerator.v:2300" *)
  wire _T_3334;
  (* src = "crypto_accelerator.v:2301" *)
  wire _T_3336;
  (* src = "crypto_accelerator.v:2302" *)
  wire _T_3338;
  (* src = "crypto_accelerator.v:2303" *)
  wire _T_3340;
  (* src = "crypto_accelerator.v:2304" *)
  wire _T_3342;
  (* src = "crypto_accelerator.v:2305" *)
  wire _T_3344;
  (* src = "crypto_accelerator.v:2306" *)
  wire _T_3346;
  (* src = "crypto_accelerator.v:2307" *)
  wire _T_3348;
  (* src = "crypto_accelerator.v:2308" *)
  wire _T_3350;
  (* src = "crypto_accelerator.v:2309" *)
  wire _T_3352;
  (* src = "crypto_accelerator.v:2310" *)
  wire _T_3354;
  (* src = "crypto_accelerator.v:2311" *)
  wire _T_3356;
  (* src = "crypto_accelerator.v:2312" *)
  wire _T_3358;
  (* src = "crypto_accelerator.v:2313" *)
  wire _T_3360;
  (* src = "crypto_accelerator.v:2314" *)
  wire _T_3362;
  (* src = "crypto_accelerator.v:2315" *)
  wire _T_3364;
  (* src = "crypto_accelerator.v:2316" *)
  wire _T_3366;
  (* src = "crypto_accelerator.v:2317" *)
  wire _T_3368;
  (* src = "crypto_accelerator.v:2318" *)
  wire _T_3370;
  (* src = "crypto_accelerator.v:2319" *)
  wire _T_3372;
  (* src = "crypto_accelerator.v:2320" *)
  wire _T_3374;
  (* src = "crypto_accelerator.v:2321" *)
  wire _T_3376;
  (* src = "crypto_accelerator.v:2322" *)
  wire _T_3378;
  (* src = "crypto_accelerator.v:2323" *)
  wire _T_3380;
  (* src = "crypto_accelerator.v:2324" *)
  wire _T_3382;
  (* src = "crypto_accelerator.v:2325" *)
  wire _T_3384;
  (* src = "crypto_accelerator.v:2326" *)
  wire _T_3386;
  (* src = "crypto_accelerator.v:2327" *)
  wire _T_3388;
  (* src = "crypto_accelerator.v:2328" *)
  wire _T_3390;
  (* src = "crypto_accelerator.v:2329" *)
  wire _T_3392;
  (* src = "crypto_accelerator.v:2330" *)
  wire _T_3394;
  (* src = "crypto_accelerator.v:2331" *)
  wire _T_3396;
  (* src = "crypto_accelerator.v:2332" *)
  wire _T_3398;
  (* src = "crypto_accelerator.v:2333" *)
  wire _T_3400;
  (* src = "crypto_accelerator.v:2334" *)
  wire _T_3402;
  (* src = "crypto_accelerator.v:2335" *)
  wire _T_3404;
  (* src = "crypto_accelerator.v:2336" *)
  wire _T_3406;
  (* src = "crypto_accelerator.v:2337" *)
  wire _T_3408;
  (* src = "crypto_accelerator.v:2338" *)
  wire _T_3410;
  (* src = "crypto_accelerator.v:2339" *)
  wire _T_3412;
  (* src = "crypto_accelerator.v:2340" *)
  wire _T_3414;
  (* src = "crypto_accelerator.v:2341" *)
  wire _T_3416;
  (* src = "crypto_accelerator.v:2342" *)
  wire _T_3418;
  (* src = "crypto_accelerator.v:2343" *)
  wire _T_3420;
  (* src = "crypto_accelerator.v:2344" *)
  wire _T_3422;
  (* src = "crypto_accelerator.v:2345" *)
  wire _T_3424;
  (* src = "crypto_accelerator.v:2346" *)
  wire _T_3426;
  (* src = "crypto_accelerator.v:2347" *)
  wire _T_3428;
  (* src = "crypto_accelerator.v:2348" *)
  wire _T_3430;
  (* src = "crypto_accelerator.v:2349" *)
  wire _T_3432;
  (* src = "crypto_accelerator.v:2350" *)
  wire _T_3434;
  (* src = "crypto_accelerator.v:2351" *)
  wire _T_3436;
  (* src = "crypto_accelerator.v:2352" *)
  wire _T_3438;
  (* src = "crypto_accelerator.v:2353" *)
  wire _T_3440;
  (* src = "crypto_accelerator.v:2354" *)
  wire _T_3442;
  (* src = "crypto_accelerator.v:2355" *)
  wire _T_3444;
  (* src = "crypto_accelerator.v:2356" *)
  wire _T_3446;
  (* src = "crypto_accelerator.v:2357" *)
  wire _T_3448;
  (* src = "crypto_accelerator.v:2358" *)
  wire _T_3450;
  (* src = "crypto_accelerator.v:2359" *)
  wire _T_3452;
  (* src = "crypto_accelerator.v:2360" *)
  wire _T_3454;
  (* src = "crypto_accelerator.v:2361" *)
  wire _T_3456;
  (* src = "crypto_accelerator.v:2362" *)
  wire _T_3458;
  (* src = "crypto_accelerator.v:2363" *)
  wire _T_3460;
  (* src = "crypto_accelerator.v:2364" *)
  wire _T_3462;
  (* src = "crypto_accelerator.v:2365" *)
  wire _T_3464;
  (* src = "crypto_accelerator.v:2366" *)
  wire _T_3466;
  (* src = "crypto_accelerator.v:2367" *)
  wire _T_3468;
  (* src = "crypto_accelerator.v:2368" *)
  wire _T_3470;
  (* src = "crypto_accelerator.v:2369" *)
  wire _T_3472;
  (* src = "crypto_accelerator.v:2370" *)
  wire _T_3474;
  (* src = "crypto_accelerator.v:2371" *)
  wire _T_3476;
  (* src = "crypto_accelerator.v:2372" *)
  wire _T_3478;
  (* src = "crypto_accelerator.v:858" *)
  wire _T_348;
  (* src = "crypto_accelerator.v:2373" *)
  wire _T_3480;
  (* src = "crypto_accelerator.v:2374" *)
  wire _T_3482;
  (* src = "crypto_accelerator.v:2375" *)
  wire _T_3484;
  (* src = "crypto_accelerator.v:2376" *)
  wire _T_3486;
  (* src = "crypto_accelerator.v:2377" *)
  wire _T_3488;
  (* src = "crypto_accelerator.v:2378" *)
  wire _T_3490;
  (* src = "crypto_accelerator.v:2379" *)
  wire _T_3492;
  (* src = "crypto_accelerator.v:2380" *)
  wire _T_3494;
  (* src = "crypto_accelerator.v:2381" *)
  wire _T_3496;
  (* src = "crypto_accelerator.v:2382" *)
  wire _T_3498;
  (* src = "crypto_accelerator.v:859" *)
  wire _T_350;
  (* src = "crypto_accelerator.v:2383" *)
  wire _T_3500;
  (* src = "crypto_accelerator.v:2384" *)
  wire _T_3502;
  (* src = "crypto_accelerator.v:2385" *)
  wire _T_3504;
  (* src = "crypto_accelerator.v:2386" *)
  wire _T_3506;
  (* src = "crypto_accelerator.v:2387" *)
  wire _T_3508;
  (* src = "crypto_accelerator.v:2388" *)
  wire _T_3510;
  (* src = "crypto_accelerator.v:2389" *)
  wire _T_3512;
  (* src = "crypto_accelerator.v:2390" *)
  wire _T_3514;
  (* src = "crypto_accelerator.v:2391" *)
  wire _T_3516;
  (* src = "crypto_accelerator.v:2392" *)
  wire _T_3518;
  (* src = "crypto_accelerator.v:860" *)
  wire _T_352;
  (* src = "crypto_accelerator.v:2393" *)
  wire _T_3520;
  (* src = "crypto_accelerator.v:2394" *)
  wire _T_3522;
  (* src = "crypto_accelerator.v:2395" *)
  wire _T_3524;
  (* src = "crypto_accelerator.v:2396" *)
  wire _T_3526;
  (* src = "crypto_accelerator.v:2397" *)
  wire _T_3527;
  (* src = "crypto_accelerator.v:2398" *)
  wire _T_3528;
  (* src = "crypto_accelerator.v:2399" *)
  wire _T_3529;
  (* src = "crypto_accelerator.v:2400" *)
  wire _T_3531;
  (* src = "crypto_accelerator.v:2401" *)
  wire _T_3532;
  (* src = "crypto_accelerator.v:2402" *)
  wire _T_3533;
  (* src = "crypto_accelerator.v:2403" *)
  wire _T_3535;
  (* src = "crypto_accelerator.v:2404" *)
  wire _T_3537;
  (* src = "crypto_accelerator.v:2405" *)
  wire _T_3538;
  (* src = "crypto_accelerator.v:2406" *)
  wire _T_3539;
  (* src = "crypto_accelerator.v:861" *)
  wire _T_354;
  (* src = "crypto_accelerator.v:2407" *)
  wire _T_3541;
  (* src = "crypto_accelerator.v:2408" *)
  wire _T_3543;
  (* src = "crypto_accelerator.v:2409" *)
  wire _T_3545;
  (* src = "crypto_accelerator.v:2410" *)
  wire _T_3546;
  (* src = "crypto_accelerator.v:2411" *)
  wire _T_3547;
  (* src = "crypto_accelerator.v:2412" *)
  wire _T_3549;
  (* src = "crypto_accelerator.v:2413" *)
  wire _T_3550;
  (* src = "crypto_accelerator.v:2414" *)
  wire _T_3552;
  (* src = "crypto_accelerator.v:2415" *)
  wire _T_3553;
  (* src = "crypto_accelerator.v:2416" *)
  wire _T_3554;
  (* src = "crypto_accelerator.v:862" *)
  wire _T_356;
  (* src = "crypto_accelerator.v:2418" *)
  wire _T_3579;
  (* src = "crypto_accelerator.v:863" *)
  wire _T_358;
  (* src = "crypto_accelerator.v:2419" *)
  wire _T_3581;
  (* src = "crypto_accelerator.v:2420" *)
  wire _T_3583;
  (* src = "crypto_accelerator.v:2421" *)
  wire _T_3585;
  (* src = "crypto_accelerator.v:2422" *)
  wire _T_3587;
  (* src = "crypto_accelerator.v:2423" *)
  wire _T_3589;
  (* src = "crypto_accelerator.v:2424" *)
  wire _T_3591;
  (* src = "crypto_accelerator.v:2425" *)
  wire _T_3593;
  (* src = "crypto_accelerator.v:2426" *)
  wire _T_3595;
  (* src = "crypto_accelerator.v:2427" *)
  wire _T_3597;
  (* src = "crypto_accelerator.v:2428" *)
  wire _T_3599;
  (* src = "crypto_accelerator.v:864" *)
  wire _T_360;
  (* src = "crypto_accelerator.v:2429" *)
  wire _T_3601;
  (* src = "crypto_accelerator.v:2430" *)
  wire _T_3603;
  (* src = "crypto_accelerator.v:2431" *)
  wire _T_3605;
  (* src = "crypto_accelerator.v:2432" *)
  wire _T_3607;
  (* src = "crypto_accelerator.v:2433" *)
  wire _T_3609;
  (* src = "crypto_accelerator.v:2434" *)
  wire _T_3611;
  (* src = "crypto_accelerator.v:2435" *)
  wire _T_3613;
  (* src = "crypto_accelerator.v:2436" *)
  wire _T_3615;
  (* src = "crypto_accelerator.v:2437" *)
  wire _T_3617;
  (* src = "crypto_accelerator.v:2438" *)
  wire _T_3619;
  (* src = "crypto_accelerator.v:865" *)
  wire _T_362;
  (* src = "crypto_accelerator.v:2439" *)
  wire _T_3621;
  (* src = "crypto_accelerator.v:2440" *)
  wire _T_3623;
  (* src = "crypto_accelerator.v:2441" *)
  wire _T_3625;
  (* src = "crypto_accelerator.v:2442" *)
  wire _T_3627;
  (* src = "crypto_accelerator.v:2443" *)
  wire _T_3629;
  (* src = "crypto_accelerator.v:2444" *)
  wire _T_3631;
  (* src = "crypto_accelerator.v:2445" *)
  wire _T_3633;
  (* src = "crypto_accelerator.v:2446" *)
  wire _T_3635;
  (* src = "crypto_accelerator.v:2447" *)
  wire _T_3637;
  (* src = "crypto_accelerator.v:2448" *)
  wire _T_3639;
  (* src = "crypto_accelerator.v:866" *)
  wire _T_364;
  (* src = "crypto_accelerator.v:2449" *)
  wire _T_3641;
  (* src = "crypto_accelerator.v:2450" *)
  wire _T_3643;
  (* src = "crypto_accelerator.v:2451" *)
  wire _T_3645;
  (* src = "crypto_accelerator.v:2452" *)
  wire _T_3647;
  (* src = "crypto_accelerator.v:2453" *)
  wire _T_3649;
  (* src = "crypto_accelerator.v:2454" *)
  wire _T_3651;
  (* src = "crypto_accelerator.v:2455" *)
  wire _T_3653;
  (* src = "crypto_accelerator.v:2456" *)
  wire _T_3655;
  (* src = "crypto_accelerator.v:2457" *)
  wire _T_3657;
  (* src = "crypto_accelerator.v:2458" *)
  wire _T_3659;
  (* src = "crypto_accelerator.v:867" *)
  wire _T_366;
  (* src = "crypto_accelerator.v:2459" *)
  wire _T_3661;
  (* src = "crypto_accelerator.v:2460" *)
  wire _T_3663;
  (* src = "crypto_accelerator.v:2461" *)
  wire _T_3665;
  (* src = "crypto_accelerator.v:2462" *)
  wire _T_3667;
  (* src = "crypto_accelerator.v:2463" *)
  wire _T_3669;
  (* src = "crypto_accelerator.v:2464" *)
  wire _T_3671;
  (* src = "crypto_accelerator.v:2465" *)
  wire _T_3673;
  (* src = "crypto_accelerator.v:2466" *)
  wire _T_3675;
  (* src = "crypto_accelerator.v:2467" *)
  wire _T_3677;
  (* src = "crypto_accelerator.v:2468" *)
  wire _T_3679;
  (* src = "crypto_accelerator.v:868" *)
  wire _T_368;
  (* src = "crypto_accelerator.v:2469" *)
  wire _T_3681;
  (* src = "crypto_accelerator.v:2470" *)
  wire _T_3683;
  (* src = "crypto_accelerator.v:2471" *)
  wire _T_3685;
  (* src = "crypto_accelerator.v:2472" *)
  wire _T_3687;
  (* src = "crypto_accelerator.v:2473" *)
  wire _T_3689;
  (* src = "crypto_accelerator.v:2474" *)
  wire _T_3691;
  (* src = "crypto_accelerator.v:2475" *)
  wire _T_3693;
  (* src = "crypto_accelerator.v:2476" *)
  wire _T_3695;
  (* src = "crypto_accelerator.v:2477" *)
  wire _T_3697;
  (* src = "crypto_accelerator.v:2478" *)
  wire _T_3699;
  (* src = "crypto_accelerator.v:869" *)
  wire _T_370;
  (* src = "crypto_accelerator.v:2479" *)
  wire _T_3701;
  (* src = "crypto_accelerator.v:2480" *)
  wire _T_3703;
  (* src = "crypto_accelerator.v:2481" *)
  wire _T_3705;
  (* src = "crypto_accelerator.v:2482" *)
  wire _T_3707;
  (* src = "crypto_accelerator.v:2483" *)
  wire _T_3709;
  (* src = "crypto_accelerator.v:2484" *)
  wire _T_3711;
  (* src = "crypto_accelerator.v:2485" *)
  wire _T_3713;
  (* src = "crypto_accelerator.v:2486" *)
  wire _T_3715;
  (* src = "crypto_accelerator.v:2487" *)
  wire _T_3717;
  (* src = "crypto_accelerator.v:2488" *)
  wire _T_3719;
  (* src = "crypto_accelerator.v:870" *)
  wire _T_372;
  (* src = "crypto_accelerator.v:2489" *)
  wire _T_3721;
  (* src = "crypto_accelerator.v:2490" *)
  wire _T_3723;
  (* src = "crypto_accelerator.v:2491" *)
  wire _T_3725;
  (* src = "crypto_accelerator.v:2492" *)
  wire _T_3727;
  (* src = "crypto_accelerator.v:2493" *)
  wire _T_3729;
  (* src = "crypto_accelerator.v:2494" *)
  wire _T_3731;
  (* src = "crypto_accelerator.v:2495" *)
  wire _T_3733;
  (* src = "crypto_accelerator.v:2496" *)
  wire _T_3735;
  (* src = "crypto_accelerator.v:2497" *)
  wire _T_3737;
  (* src = "crypto_accelerator.v:2498" *)
  wire _T_3739;
  (* src = "crypto_accelerator.v:871" *)
  wire _T_374;
  (* src = "crypto_accelerator.v:2499" *)
  wire _T_3741;
  (* src = "crypto_accelerator.v:2500" *)
  wire _T_3743;
  (* src = "crypto_accelerator.v:2501" *)
  wire _T_3745;
  (* src = "crypto_accelerator.v:2502" *)
  wire _T_3747;
  (* src = "crypto_accelerator.v:2503" *)
  wire _T_3749;
  (* src = "crypto_accelerator.v:2504" *)
  wire _T_3751;
  (* src = "crypto_accelerator.v:2505" *)
  wire _T_3753;
  (* src = "crypto_accelerator.v:2506" *)
  wire _T_3755;
  (* src = "crypto_accelerator.v:2507" *)
  wire _T_3757;
  (* src = "crypto_accelerator.v:2508" *)
  wire _T_3759;
  (* src = "crypto_accelerator.v:872" *)
  wire _T_376;
  (* src = "crypto_accelerator.v:2509" *)
  wire _T_3761;
  (* src = "crypto_accelerator.v:2510" *)
  wire _T_3763;
  (* src = "crypto_accelerator.v:2511" *)
  wire _T_3765;
  (* src = "crypto_accelerator.v:2512" *)
  wire _T_3767;
  (* src = "crypto_accelerator.v:2513" *)
  wire _T_3769;
  (* src = "crypto_accelerator.v:2514" *)
  wire _T_3771;
  (* src = "crypto_accelerator.v:2515" *)
  wire _T_3773;
  (* src = "crypto_accelerator.v:2516" *)
  wire _T_3775;
  (* src = "crypto_accelerator.v:2517" *)
  wire _T_3777;
  (* src = "crypto_accelerator.v:2518" *)
  wire _T_3779;
  (* src = "crypto_accelerator.v:873" *)
  wire _T_378;
  (* src = "crypto_accelerator.v:2519" *)
  wire _T_3781;
  (* src = "crypto_accelerator.v:2520" *)
  wire _T_3783;
  (* src = "crypto_accelerator.v:2521" *)
  wire _T_3785;
  (* src = "crypto_accelerator.v:2522" *)
  wire _T_3787;
  (* src = "crypto_accelerator.v:2523" *)
  wire _T_3789;
  (* src = "crypto_accelerator.v:2524" *)
  wire _T_3791;
  (* src = "crypto_accelerator.v:2525" *)
  wire _T_3793;
  (* src = "crypto_accelerator.v:2526" *)
  wire _T_3795;
  (* src = "crypto_accelerator.v:2527" *)
  wire _T_3796;
  (* src = "crypto_accelerator.v:2528" *)
  wire _T_3797;
  (* src = "crypto_accelerator.v:2529" *)
  wire _T_3798;
  (* src = "crypto_accelerator.v:874" *)
  wire _T_380;
  (* src = "crypto_accelerator.v:2530" *)
  wire _T_3800;
  (* src = "crypto_accelerator.v:2531" *)
  wire _T_3801;
  (* src = "crypto_accelerator.v:2532" *)
  wire _T_3802;
  (* src = "crypto_accelerator.v:2533" *)
  wire _T_3804;
  (* src = "crypto_accelerator.v:2534" *)
  wire _T_3806;
  (* src = "crypto_accelerator.v:2535" *)
  wire _T_3807;
  (* src = "crypto_accelerator.v:2536" *)
  wire _T_3808;
  (* src = "crypto_accelerator.v:2537" *)
  wire _T_3810;
  (* src = "crypto_accelerator.v:2538" *)
  wire _T_3812;
  (* src = "crypto_accelerator.v:2539" *)
  wire _T_3814;
  (* src = "crypto_accelerator.v:2540" *)
  wire _T_3815;
  (* src = "crypto_accelerator.v:2541" *)
  wire _T_3816;
  (* src = "crypto_accelerator.v:2542" *)
  wire _T_3818;
  (* src = "crypto_accelerator.v:2543" *)
  wire _T_3819;
  (* src = "crypto_accelerator.v:875" *)
  wire _T_382;
  (* src = "crypto_accelerator.v:2544" *)
  wire _T_3821;
  (* src = "crypto_accelerator.v:2545" *)
  wire _T_3822;
  (* src = "crypto_accelerator.v:2546" *)
  wire _T_3823;
  (* src = "crypto_accelerator.v:876" *)
  wire _T_384;
  (* src = "crypto_accelerator.v:2548" *)
  wire _T_3848;
  (* src = "crypto_accelerator.v:2549" *)
  wire _T_3850;
  (* src = "crypto_accelerator.v:2550" *)
  wire _T_3852;
  (* src = "crypto_accelerator.v:2551" *)
  wire _T_3854;
  (* src = "crypto_accelerator.v:2552" *)
  wire _T_3856;
  (* src = "crypto_accelerator.v:2553" *)
  wire _T_3858;
  (* src = "crypto_accelerator.v:877" *)
  wire _T_386;
  (* src = "crypto_accelerator.v:2554" *)
  wire _T_3860;
  (* src = "crypto_accelerator.v:2555" *)
  wire _T_3862;
  (* src = "crypto_accelerator.v:2556" *)
  wire _T_3864;
  (* src = "crypto_accelerator.v:2557" *)
  wire _T_3866;
  (* src = "crypto_accelerator.v:2558" *)
  wire _T_3868;
  (* src = "crypto_accelerator.v:2559" *)
  wire _T_3870;
  (* src = "crypto_accelerator.v:2560" *)
  wire _T_3872;
  (* src = "crypto_accelerator.v:2561" *)
  wire _T_3874;
  (* src = "crypto_accelerator.v:2562" *)
  wire _T_3876;
  (* src = "crypto_accelerator.v:2563" *)
  wire _T_3878;
  (* src = "crypto_accelerator.v:878" *)
  wire _T_388;
  (* src = "crypto_accelerator.v:2564" *)
  wire _T_3880;
  (* src = "crypto_accelerator.v:2565" *)
  wire _T_3882;
  (* src = "crypto_accelerator.v:2566" *)
  wire _T_3884;
  (* src = "crypto_accelerator.v:2567" *)
  wire _T_3886;
  (* src = "crypto_accelerator.v:2568" *)
  wire _T_3888;
  (* src = "crypto_accelerator.v:2569" *)
  wire _T_3890;
  (* src = "crypto_accelerator.v:2570" *)
  wire _T_3892;
  (* src = "crypto_accelerator.v:2571" *)
  wire _T_3894;
  (* src = "crypto_accelerator.v:2572" *)
  wire _T_3896;
  (* src = "crypto_accelerator.v:2573" *)
  wire _T_3898;
  (* src = "crypto_accelerator.v:879" *)
  wire _T_390;
  (* src = "crypto_accelerator.v:2574" *)
  wire _T_3900;
  (* src = "crypto_accelerator.v:2575" *)
  wire _T_3902;
  (* src = "crypto_accelerator.v:2576" *)
  wire _T_3904;
  (* src = "crypto_accelerator.v:2577" *)
  wire _T_3906;
  (* src = "crypto_accelerator.v:2578" *)
  wire _T_3908;
  (* src = "crypto_accelerator.v:2579" *)
  wire _T_3910;
  (* src = "crypto_accelerator.v:2580" *)
  wire _T_3912;
  (* src = "crypto_accelerator.v:2581" *)
  wire _T_3914;
  (* src = "crypto_accelerator.v:2582" *)
  wire _T_3916;
  (* src = "crypto_accelerator.v:2583" *)
  wire _T_3918;
  (* src = "crypto_accelerator.v:880" *)
  wire _T_392;
  (* src = "crypto_accelerator.v:2584" *)
  wire _T_3920;
  (* src = "crypto_accelerator.v:2585" *)
  wire _T_3922;
  (* src = "crypto_accelerator.v:2586" *)
  wire _T_3924;
  (* src = "crypto_accelerator.v:2587" *)
  wire _T_3926;
  (* src = "crypto_accelerator.v:2588" *)
  wire _T_3928;
  (* src = "crypto_accelerator.v:2589" *)
  wire _T_3930;
  (* src = "crypto_accelerator.v:2590" *)
  wire _T_3932;
  (* src = "crypto_accelerator.v:2591" *)
  wire _T_3934;
  (* src = "crypto_accelerator.v:2592" *)
  wire _T_3936;
  (* src = "crypto_accelerator.v:2593" *)
  wire _T_3938;
  (* src = "crypto_accelerator.v:881" *)
  wire _T_394;
  (* src = "crypto_accelerator.v:2594" *)
  wire _T_3940;
  (* src = "crypto_accelerator.v:2595" *)
  wire _T_3942;
  (* src = "crypto_accelerator.v:2596" *)
  wire _T_3944;
  (* src = "crypto_accelerator.v:2597" *)
  wire _T_3946;
  (* src = "crypto_accelerator.v:2598" *)
  wire _T_3948;
  (* src = "crypto_accelerator.v:2599" *)
  wire _T_3950;
  (* src = "crypto_accelerator.v:2600" *)
  wire _T_3952;
  (* src = "crypto_accelerator.v:2601" *)
  wire _T_3954;
  (* src = "crypto_accelerator.v:2602" *)
  wire _T_3956;
  (* src = "crypto_accelerator.v:2603" *)
  wire _T_3958;
  (* src = "crypto_accelerator.v:882" *)
  wire _T_396;
  (* src = "crypto_accelerator.v:2604" *)
  wire _T_3960;
  (* src = "crypto_accelerator.v:2605" *)
  wire _T_3962;
  (* src = "crypto_accelerator.v:2606" *)
  wire _T_3964;
  (* src = "crypto_accelerator.v:2607" *)
  wire _T_3966;
  (* src = "crypto_accelerator.v:2608" *)
  wire _T_3968;
  (* src = "crypto_accelerator.v:2609" *)
  wire _T_3970;
  (* src = "crypto_accelerator.v:2610" *)
  wire _T_3972;
  (* src = "crypto_accelerator.v:2611" *)
  wire _T_3974;
  (* src = "crypto_accelerator.v:2612" *)
  wire _T_3976;
  (* src = "crypto_accelerator.v:2613" *)
  wire _T_3978;
  (* src = "crypto_accelerator.v:883" *)
  wire _T_398;
  (* src = "crypto_accelerator.v:2614" *)
  wire _T_3980;
  (* src = "crypto_accelerator.v:2615" *)
  wire _T_3982;
  (* src = "crypto_accelerator.v:2616" *)
  wire _T_3984;
  (* src = "crypto_accelerator.v:2617" *)
  wire _T_3986;
  (* src = "crypto_accelerator.v:2618" *)
  wire _T_3988;
  (* src = "crypto_accelerator.v:2619" *)
  wire _T_3990;
  (* src = "crypto_accelerator.v:2620" *)
  wire _T_3992;
  (* src = "crypto_accelerator.v:2621" *)
  wire _T_3994;
  (* src = "crypto_accelerator.v:2622" *)
  wire _T_3996;
  (* src = "crypto_accelerator.v:2623" *)
  wire _T_3998;
  (* src = "crypto_accelerator.v:710" *)
  wire [127:0] _T_40;
  (* src = "crypto_accelerator.v:884" *)
  wire _T_400;
  (* src = "crypto_accelerator.v:2624" *)
  wire _T_4000;
  (* src = "crypto_accelerator.v:2625" *)
  wire _T_4002;
  (* src = "crypto_accelerator.v:2626" *)
  wire _T_4004;
  (* src = "crypto_accelerator.v:2627" *)
  wire _T_4006;
  (* src = "crypto_accelerator.v:2628" *)
  wire _T_4008;
  (* src = "crypto_accelerator.v:2629" *)
  wire _T_4010;
  (* src = "crypto_accelerator.v:2630" *)
  wire _T_4012;
  (* src = "crypto_accelerator.v:2631" *)
  wire _T_4014;
  (* src = "crypto_accelerator.v:2632" *)
  wire _T_4016;
  (* src = "crypto_accelerator.v:2633" *)
  wire _T_4018;
  (* src = "crypto_accelerator.v:885" *)
  wire _T_402;
  (* src = "crypto_accelerator.v:2634" *)
  wire _T_4020;
  (* src = "crypto_accelerator.v:2635" *)
  wire _T_4022;
  (* src = "crypto_accelerator.v:2636" *)
  wire _T_4024;
  (* src = "crypto_accelerator.v:2637" *)
  wire _T_4026;
  (* src = "crypto_accelerator.v:2638" *)
  wire _T_4028;
  (* src = "crypto_accelerator.v:2639" *)
  wire _T_4030;
  (* src = "crypto_accelerator.v:2640" *)
  wire _T_4032;
  (* src = "crypto_accelerator.v:2641" *)
  wire _T_4034;
  (* src = "crypto_accelerator.v:2642" *)
  wire _T_4036;
  (* src = "crypto_accelerator.v:2643" *)
  wire _T_4038;
  (* src = "crypto_accelerator.v:886" *)
  wire _T_404;
  (* src = "crypto_accelerator.v:2644" *)
  wire _T_4040;
  (* src = "crypto_accelerator.v:2645" *)
  wire _T_4042;
  (* src = "crypto_accelerator.v:2646" *)
  wire _T_4044;
  (* src = "crypto_accelerator.v:2647" *)
  wire _T_4046;
  (* src = "crypto_accelerator.v:2648" *)
  wire _T_4048;
  (* src = "crypto_accelerator.v:2649" *)
  wire _T_4050;
  (* src = "crypto_accelerator.v:2650" *)
  wire _T_4052;
  (* src = "crypto_accelerator.v:2651" *)
  wire _T_4054;
  (* src = "crypto_accelerator.v:2652" *)
  wire _T_4056;
  (* src = "crypto_accelerator.v:2653" *)
  wire _T_4058;
  (* src = "crypto_accelerator.v:887" *)
  wire _T_406;
  (* src = "crypto_accelerator.v:2654" *)
  wire _T_4060;
  (* src = "crypto_accelerator.v:2655" *)
  wire _T_4062;
  (* src = "crypto_accelerator.v:2656" *)
  wire _T_4064;
  (* src = "crypto_accelerator.v:2657" *)
  wire _T_4065;
  (* src = "crypto_accelerator.v:2658" *)
  wire _T_4066;
  (* src = "crypto_accelerator.v:2659" *)
  wire _T_4067;
  (* src = "crypto_accelerator.v:2660" *)
  wire _T_4069;
  (* src = "crypto_accelerator.v:2661" *)
  wire _T_4070;
  (* src = "crypto_accelerator.v:2662" *)
  wire _T_4071;
  (* src = "crypto_accelerator.v:2663" *)
  wire _T_4073;
  (* src = "crypto_accelerator.v:2664" *)
  wire _T_4075;
  (* src = "crypto_accelerator.v:2665" *)
  wire _T_4076;
  (* src = "crypto_accelerator.v:2666" *)
  wire _T_4077;
  (* src = "crypto_accelerator.v:2667" *)
  wire _T_4079;
  (* src = "crypto_accelerator.v:888" *)
  wire _T_408;
  (* src = "crypto_accelerator.v:2668" *)
  wire _T_4081;
  (* src = "crypto_accelerator.v:2669" *)
  wire _T_4083;
  (* src = "crypto_accelerator.v:2670" *)
  wire _T_4084;
  (* src = "crypto_accelerator.v:2671" *)
  wire _T_4085;
  (* src = "crypto_accelerator.v:2672" *)
  wire _T_4087;
  (* src = "crypto_accelerator.v:2673" *)
  wire _T_4088;
  (* src = "crypto_accelerator.v:2674" *)
  wire _T_4090;
  (* src = "crypto_accelerator.v:2675" *)
  wire _T_4091;
  (* src = "crypto_accelerator.v:2676" *)
  wire _T_4092;
  (* src = "crypto_accelerator.v:711" *)
  wire [127:0] _T_41;
  (* src = "crypto_accelerator.v:889" *)
  wire _T_410;
  (* src = "crypto_accelerator.v:2678" *)
  wire _T_4117;
  (* src = "crypto_accelerator.v:2679" *)
  wire _T_4119;
  (* src = "crypto_accelerator.v:890" *)
  wire _T_412;
  (* src = "crypto_accelerator.v:2680" *)
  wire _T_4121;
  (* src = "crypto_accelerator.v:2681" *)
  wire _T_4123;
  (* src = "crypto_accelerator.v:2682" *)
  wire _T_4125;
  (* src = "crypto_accelerator.v:2683" *)
  wire _T_4127;
  (* src = "crypto_accelerator.v:2684" *)
  wire _T_4129;
  (* src = "crypto_accelerator.v:2685" *)
  wire _T_4131;
  (* src = "crypto_accelerator.v:2686" *)
  wire _T_4133;
  (* src = "crypto_accelerator.v:2687" *)
  wire _T_4135;
  (* src = "crypto_accelerator.v:2688" *)
  wire _T_4137;
  (* src = "crypto_accelerator.v:2689" *)
  wire _T_4139;
  (* src = "crypto_accelerator.v:891" *)
  wire _T_414;
  (* src = "crypto_accelerator.v:2690" *)
  wire _T_4141;
  (* src = "crypto_accelerator.v:2691" *)
  wire _T_4143;
  (* src = "crypto_accelerator.v:2692" *)
  wire _T_4145;
  (* src = "crypto_accelerator.v:2693" *)
  wire _T_4147;
  (* src = "crypto_accelerator.v:2694" *)
  wire _T_4149;
  (* src = "crypto_accelerator.v:2695" *)
  wire _T_4151;
  (* src = "crypto_accelerator.v:2696" *)
  wire _T_4153;
  (* src = "crypto_accelerator.v:2697" *)
  wire _T_4155;
  (* src = "crypto_accelerator.v:2698" *)
  wire _T_4157;
  (* src = "crypto_accelerator.v:2699" *)
  wire _T_4159;
  (* src = "crypto_accelerator.v:892" *)
  wire _T_416;
  (* src = "crypto_accelerator.v:2700" *)
  wire _T_4161;
  (* src = "crypto_accelerator.v:2701" *)
  wire _T_4163;
  (* src = "crypto_accelerator.v:2702" *)
  wire _T_4165;
  (* src = "crypto_accelerator.v:2703" *)
  wire _T_4167;
  (* src = "crypto_accelerator.v:2704" *)
  wire _T_4169;
  (* src = "crypto_accelerator.v:2705" *)
  wire _T_4171;
  (* src = "crypto_accelerator.v:2706" *)
  wire _T_4173;
  (* src = "crypto_accelerator.v:2707" *)
  wire _T_4175;
  (* src = "crypto_accelerator.v:2708" *)
  wire _T_4177;
  (* src = "crypto_accelerator.v:2709" *)
  wire _T_4179;
  (* src = "crypto_accelerator.v:893" *)
  wire _T_418;
  (* src = "crypto_accelerator.v:2710" *)
  wire _T_4181;
  (* src = "crypto_accelerator.v:2711" *)
  wire _T_4183;
  (* src = "crypto_accelerator.v:2712" *)
  wire _T_4185;
  (* src = "crypto_accelerator.v:2713" *)
  wire _T_4187;
  (* src = "crypto_accelerator.v:2714" *)
  wire _T_4189;
  (* src = "crypto_accelerator.v:2715" *)
  wire _T_4191;
  (* src = "crypto_accelerator.v:2716" *)
  wire _T_4193;
  (* src = "crypto_accelerator.v:2717" *)
  wire _T_4195;
  (* src = "crypto_accelerator.v:2718" *)
  wire _T_4197;
  (* src = "crypto_accelerator.v:2719" *)
  wire _T_4199;
  (* src = "crypto_accelerator.v:894" *)
  wire _T_420;
  (* src = "crypto_accelerator.v:2720" *)
  wire _T_4201;
  (* src = "crypto_accelerator.v:2721" *)
  wire _T_4203;
  (* src = "crypto_accelerator.v:2722" *)
  wire _T_4205;
  (* src = "crypto_accelerator.v:2723" *)
  wire _T_4207;
  (* src = "crypto_accelerator.v:2724" *)
  wire _T_4209;
  (* src = "crypto_accelerator.v:2725" *)
  wire _T_4211;
  (* src = "crypto_accelerator.v:2726" *)
  wire _T_4213;
  (* src = "crypto_accelerator.v:2727" *)
  wire _T_4215;
  (* src = "crypto_accelerator.v:2728" *)
  wire _T_4217;
  (* src = "crypto_accelerator.v:2729" *)
  wire _T_4219;
  (* src = "crypto_accelerator.v:895" *)
  wire _T_422;
  (* src = "crypto_accelerator.v:2730" *)
  wire _T_4221;
  (* src = "crypto_accelerator.v:2731" *)
  wire _T_4223;
  (* src = "crypto_accelerator.v:2732" *)
  wire _T_4225;
  (* src = "crypto_accelerator.v:2733" *)
  wire _T_4227;
  (* src = "crypto_accelerator.v:2734" *)
  wire _T_4229;
  (* src = "crypto_accelerator.v:2735" *)
  wire _T_4231;
  (* src = "crypto_accelerator.v:2736" *)
  wire _T_4233;
  (* src = "crypto_accelerator.v:2737" *)
  wire _T_4235;
  (* src = "crypto_accelerator.v:2738" *)
  wire _T_4237;
  (* src = "crypto_accelerator.v:2739" *)
  wire _T_4239;
  (* src = "crypto_accelerator.v:896" *)
  wire _T_424;
  (* src = "crypto_accelerator.v:2740" *)
  wire _T_4241;
  (* src = "crypto_accelerator.v:2741" *)
  wire _T_4243;
  (* src = "crypto_accelerator.v:2742" *)
  wire _T_4245;
  (* src = "crypto_accelerator.v:2743" *)
  wire _T_4247;
  (* src = "crypto_accelerator.v:2744" *)
  wire _T_4249;
  (* src = "crypto_accelerator.v:2745" *)
  wire _T_4251;
  (* src = "crypto_accelerator.v:2746" *)
  wire _T_4253;
  (* src = "crypto_accelerator.v:2747" *)
  wire _T_4255;
  (* src = "crypto_accelerator.v:2748" *)
  wire _T_4257;
  (* src = "crypto_accelerator.v:2749" *)
  wire _T_4259;
  (* src = "crypto_accelerator.v:897" *)
  wire _T_426;
  (* src = "crypto_accelerator.v:2750" *)
  wire _T_4261;
  (* src = "crypto_accelerator.v:2751" *)
  wire _T_4263;
  (* src = "crypto_accelerator.v:2752" *)
  wire _T_4265;
  (* src = "crypto_accelerator.v:2753" *)
  wire _T_4267;
  (* src = "crypto_accelerator.v:2754" *)
  wire _T_4269;
  (* src = "crypto_accelerator.v:2755" *)
  wire _T_4271;
  (* src = "crypto_accelerator.v:2756" *)
  wire _T_4273;
  (* src = "crypto_accelerator.v:2757" *)
  wire _T_4275;
  (* src = "crypto_accelerator.v:2758" *)
  wire _T_4277;
  (* src = "crypto_accelerator.v:2759" *)
  wire _T_4279;
  (* src = "crypto_accelerator.v:898" *)
  wire _T_428;
  (* src = "crypto_accelerator.v:2760" *)
  wire _T_4281;
  (* src = "crypto_accelerator.v:2761" *)
  wire _T_4283;
  (* src = "crypto_accelerator.v:2762" *)
  wire _T_4285;
  (* src = "crypto_accelerator.v:2763" *)
  wire _T_4287;
  (* src = "crypto_accelerator.v:2764" *)
  wire _T_4289;
  (* src = "crypto_accelerator.v:2765" *)
  wire _T_4291;
  (* src = "crypto_accelerator.v:2766" *)
  wire _T_4293;
  (* src = "crypto_accelerator.v:2767" *)
  wire _T_4295;
  (* src = "crypto_accelerator.v:2768" *)
  wire _T_4297;
  (* src = "crypto_accelerator.v:2769" *)
  wire _T_4299;
  (* src = "crypto_accelerator.v:899" *)
  wire _T_430;
  (* src = "crypto_accelerator.v:2770" *)
  wire _T_4301;
  (* src = "crypto_accelerator.v:2771" *)
  wire _T_4303;
  (* src = "crypto_accelerator.v:2772" *)
  wire _T_4305;
  (* src = "crypto_accelerator.v:2773" *)
  wire _T_4307;
  (* src = "crypto_accelerator.v:2774" *)
  wire _T_4309;
  (* src = "crypto_accelerator.v:2775" *)
  wire _T_4311;
  (* src = "crypto_accelerator.v:2776" *)
  wire _T_4313;
  (* src = "crypto_accelerator.v:2777" *)
  wire _T_4315;
  (* src = "crypto_accelerator.v:2778" *)
  wire _T_4317;
  (* src = "crypto_accelerator.v:2779" *)
  wire _T_4319;
  (* src = "crypto_accelerator.v:900" *)
  wire _T_432;
  (* src = "crypto_accelerator.v:2780" *)
  wire _T_4321;
  (* src = "crypto_accelerator.v:2781" *)
  wire _T_4323;
  (* src = "crypto_accelerator.v:2782" *)
  wire _T_4325;
  (* src = "crypto_accelerator.v:2783" *)
  wire _T_4327;
  (* src = "crypto_accelerator.v:2784" *)
  wire _T_4329;
  (* src = "crypto_accelerator.v:2785" *)
  wire _T_4331;
  (* src = "crypto_accelerator.v:2786" *)
  wire _T_4333;
  (* src = "crypto_accelerator.v:2787" *)
  wire _T_4334;
  (* src = "crypto_accelerator.v:2788" *)
  wire _T_4335;
  (* src = "crypto_accelerator.v:2789" *)
  wire _T_4336;
  (* src = "crypto_accelerator.v:2790" *)
  wire _T_4338;
  (* src = "crypto_accelerator.v:2791" *)
  wire _T_4339;
  (* src = "crypto_accelerator.v:901" *)
  wire _T_434;
  (* src = "crypto_accelerator.v:2792" *)
  wire _T_4340;
  (* src = "crypto_accelerator.v:2793" *)
  wire _T_4342;
  (* src = "crypto_accelerator.v:2794" *)
  wire _T_4344;
  (* src = "crypto_accelerator.v:2795" *)
  wire _T_4345;
  (* src = "crypto_accelerator.v:2796" *)
  wire _T_4346;
  (* src = "crypto_accelerator.v:2797" *)
  wire _T_4348;
  (* src = "crypto_accelerator.v:2798" *)
  wire _T_4350;
  (* src = "crypto_accelerator.v:2799" *)
  wire _T_4352;
  (* src = "crypto_accelerator.v:2800" *)
  wire _T_4353;
  (* src = "crypto_accelerator.v:2801" *)
  wire _T_4354;
  (* src = "crypto_accelerator.v:2802" *)
  wire _T_4356;
  (* src = "crypto_accelerator.v:2803" *)
  wire _T_4357;
  (* src = "crypto_accelerator.v:2804" *)
  wire _T_4359;
  (* src = "crypto_accelerator.v:902" *)
  wire _T_436;
  (* src = "crypto_accelerator.v:2805" *)
  wire _T_4360;
  (* src = "crypto_accelerator.v:2806" *)
  wire _T_4361;
  (* src = "crypto_accelerator.v:903" *)
  wire _T_438;
  (* src = "crypto_accelerator.v:904" *)
  wire _T_440;
  (* src = "crypto_accelerator.v:2840" *)
  wire _T_4415;
  (* src = "crypto_accelerator.v:905" *)
  wire _T_442;
  (* src = "crypto_accelerator.v:2841" *)
  wire _T_4420;
  (* src = "crypto_accelerator.v:2842" *)
  wire _T_4421;
  (* src = "crypto_accelerator.v:2843" *)
  wire _T_4422;
  (* src = "crypto_accelerator.v:2846" *)
  wire [5:0] _T_4427;
  (* src = "crypto_accelerator.v:906" *)
  wire _T_444;
  (* src = "crypto_accelerator.v:907" *)
  wire _T_446;
  (* src = "crypto_accelerator.v:908" *)
  wire _T_448;
  (* src = "crypto_accelerator.v:909" *)
  wire _T_450;
  (* src = "crypto_accelerator.v:910" *)
  wire _T_452;
  (* src = "crypto_accelerator.v:911" *)
  wire _T_454;
  (* src = "crypto_accelerator.v:912" *)
  wire _T_456;
  (* src = "crypto_accelerator.v:913" *)
  wire _T_458;
  (* src = "crypto_accelerator.v:914" *)
  wire _T_460;
  (* src = "crypto_accelerator.v:915" *)
  wire _T_462;
  (* src = "crypto_accelerator.v:916" *)
  wire _T_464;
  (* src = "crypto_accelerator.v:917" *)
  wire _T_466;
  (* src = "crypto_accelerator.v:918" *)
  wire _T_468;
  (* src = "crypto_accelerator.v:919" *)
  wire _T_470;
  (* src = "crypto_accelerator.v:920" *)
  wire _T_472;
  (* src = "crypto_accelerator.v:921" *)
  wire _T_474;
  (* src = "crypto_accelerator.v:922" *)
  wire _T_476;
  (* src = "crypto_accelerator.v:923" *)
  wire _T_478;
  (* src = "crypto_accelerator.v:924" *)
  wire _T_480;
  (* src = "crypto_accelerator.v:925" *)
  wire _T_482;
  (* src = "crypto_accelerator.v:926" *)
  wire _T_484;
  (* src = "crypto_accelerator.v:927" *)
  wire _T_486;
  (* src = "crypto_accelerator.v:928" *)
  wire _T_488;
  (* src = "crypto_accelerator.v:929" *)
  wire _T_490;
  (* src = "crypto_accelerator.v:930" *)
  wire _T_492;
  (* src = "crypto_accelerator.v:931" *)
  wire _T_494;
  (* src = "crypto_accelerator.v:932" *)
  wire _T_496;
  (* src = "crypto_accelerator.v:933" *)
  wire _T_498;
  (* src = "crypto_accelerator.v:934" *)
  wire _T_500;
  (* src = "crypto_accelerator.v:935" *)
  wire _T_502;
  (* src = "crypto_accelerator.v:936" *)
  wire _T_504;
  (* src = "crypto_accelerator.v:937" *)
  wire _T_506;
  (* src = "crypto_accelerator.v:938" *)
  wire _T_508;
  (* src = "crypto_accelerator.v:939" *)
  wire _T_510;
  (* src = "crypto_accelerator.v:940" *)
  wire _T_512;
  (* src = "crypto_accelerator.v:941" *)
  wire _T_514;
  (* src = "crypto_accelerator.v:942" *)
  wire _T_516;
  (* src = "crypto_accelerator.v:943" *)
  wire _T_518;
  (* src = "crypto_accelerator.v:944" *)
  wire _T_520;
  (* src = "crypto_accelerator.v:945" *)
  wire _T_522;
  (* src = "crypto_accelerator.v:946" *)
  wire _T_524;
  (* src = "crypto_accelerator.v:947" *)
  wire _T_526;
  (* src = "crypto_accelerator.v:948" *)
  wire _T_528;
  (* src = "crypto_accelerator.v:949" *)
  wire _T_530;
  (* src = "crypto_accelerator.v:950" *)
  wire _T_532;
  (* src = "crypto_accelerator.v:951" *)
  wire _T_534;
  (* src = "crypto_accelerator.v:952" *)
  wire _T_536;
  (* src = "crypto_accelerator.v:953" *)
  wire _T_538;
  (* src = "crypto_accelerator.v:954" *)
  wire _T_540;
  (* src = "crypto_accelerator.v:955" *)
  wire _T_542;
  (* src = "crypto_accelerator.v:956" *)
  wire _T_544;
  (* src = "crypto_accelerator.v:957" *)
  wire _T_546;
  (* src = "crypto_accelerator.v:958" *)
  wire _T_548;
  (* src = "crypto_accelerator.v:959" *)
  wire _T_550;
  (* src = "crypto_accelerator.v:960" *)
  wire _T_552;
  (* src = "crypto_accelerator.v:961" *)
  wire _T_554;
  (* src = "crypto_accelerator.v:962" *)
  wire _T_556;
  (* src = "crypto_accelerator.v:963" *)
  wire _T_558;
  (* src = "crypto_accelerator.v:964" *)
  wire _T_560;
  (* src = "crypto_accelerator.v:965" *)
  wire _T_562;
  (* src = "crypto_accelerator.v:966" *)
  wire _T_564;
  (* src = "crypto_accelerator.v:967" *)
  wire _T_565;
  (* src = "crypto_accelerator.v:968" *)
  wire _T_566;
  (* src = "crypto_accelerator.v:969" *)
  wire _T_567;
  (* src = "crypto_accelerator.v:970" *)
  wire _T_569;
  (* src = "crypto_accelerator.v:971" *)
  wire _T_570;
  (* src = "crypto_accelerator.v:972" *)
  wire _T_571;
  (* src = "crypto_accelerator.v:973" *)
  wire _T_573;
  (* src = "crypto_accelerator.v:974" *)
  wire _T_575;
  (* src = "crypto_accelerator.v:975" *)
  wire _T_576;
  (* src = "crypto_accelerator.v:976" *)
  wire _T_577;
  (* src = "crypto_accelerator.v:977" *)
  wire _T_579;
  (* src = "crypto_accelerator.v:978" *)
  wire _T_581;
  (* src = "crypto_accelerator.v:979" *)
  wire _T_583;
  (* src = "crypto_accelerator.v:980" *)
  wire _T_584;
  (* src = "crypto_accelerator.v:981" *)
  wire _T_585;
  (* src = "crypto_accelerator.v:982" *)
  wire _T_587;
  (* src = "crypto_accelerator.v:983" *)
  wire _T_588;
  (* src = "crypto_accelerator.v:984" *)
  wire _T_590;
  (* src = "crypto_accelerator.v:985" *)
  wire _T_591;
  (* src = "crypto_accelerator.v:986" *)
  wire _T_592;
  (* src = "crypto_accelerator.v:689" *)
  wire _T_6;
  (* src = "crypto_accelerator.v:988" *)
  wire _T_617;
  (* src = "crypto_accelerator.v:989" *)
  wire _T_619;
  (* src = "crypto_accelerator.v:990" *)
  wire _T_621;
  (* src = "crypto_accelerator.v:991" *)
  wire _T_623;
  (* src = "crypto_accelerator.v:992" *)
  wire _T_625;
  (* src = "crypto_accelerator.v:993" *)
  wire _T_627;
  (* src = "crypto_accelerator.v:994" *)
  wire _T_629;
  (* src = "crypto_accelerator.v:995" *)
  wire _T_631;
  (* src = "crypto_accelerator.v:996" *)
  wire _T_633;
  (* src = "crypto_accelerator.v:997" *)
  wire _T_635;
  (* src = "crypto_accelerator.v:998" *)
  wire _T_637;
  (* src = "crypto_accelerator.v:999" *)
  wire _T_639;
  (* src = "crypto_accelerator.v:1000" *)
  wire _T_641;
  (* src = "crypto_accelerator.v:1001" *)
  wire _T_643;
  (* src = "crypto_accelerator.v:1002" *)
  wire _T_645;
  (* src = "crypto_accelerator.v:1003" *)
  wire _T_647;
  (* src = "crypto_accelerator.v:1004" *)
  wire _T_649;
  (* src = "crypto_accelerator.v:1005" *)
  wire _T_651;
  (* src = "crypto_accelerator.v:1006" *)
  wire _T_653;
  (* src = "crypto_accelerator.v:1007" *)
  wire _T_655;
  (* src = "crypto_accelerator.v:1008" *)
  wire _T_657;
  (* src = "crypto_accelerator.v:1009" *)
  wire _T_659;
  (* src = "crypto_accelerator.v:1010" *)
  wire _T_661;
  (* src = "crypto_accelerator.v:1011" *)
  wire _T_663;
  (* src = "crypto_accelerator.v:1012" *)
  wire _T_665;
  (* src = "crypto_accelerator.v:1013" *)
  wire _T_667;
  (* src = "crypto_accelerator.v:1014" *)
  wire _T_669;
  (* src = "crypto_accelerator.v:1015" *)
  wire _T_671;
  (* src = "crypto_accelerator.v:1016" *)
  wire _T_673;
  (* src = "crypto_accelerator.v:1017" *)
  wire _T_675;
  (* src = "crypto_accelerator.v:1018" *)
  wire _T_677;
  (* src = "crypto_accelerator.v:1019" *)
  wire _T_679;
  (* src = "crypto_accelerator.v:1020" *)
  wire _T_681;
  (* src = "crypto_accelerator.v:1021" *)
  wire _T_683;
  (* src = "crypto_accelerator.v:1022" *)
  wire _T_685;
  (* src = "crypto_accelerator.v:1023" *)
  wire _T_687;
  (* src = "crypto_accelerator.v:1024" *)
  wire _T_689;
  (* src = "crypto_accelerator.v:1025" *)
  wire _T_691;
  (* src = "crypto_accelerator.v:1026" *)
  wire _T_693;
  (* src = "crypto_accelerator.v:1027" *)
  wire _T_695;
  (* src = "crypto_accelerator.v:1028" *)
  wire _T_697;
  (* src = "crypto_accelerator.v:1029" *)
  wire _T_699;
  (* src = "crypto_accelerator.v:1030" *)
  wire _T_701;
  (* src = "crypto_accelerator.v:1031" *)
  wire _T_703;
  (* src = "crypto_accelerator.v:1032" *)
  wire _T_705;
  (* src = "crypto_accelerator.v:1033" *)
  wire _T_707;
  (* src = "crypto_accelerator.v:1034" *)
  wire _T_709;
  (* src = "crypto_accelerator.v:1035" *)
  wire _T_711;
  (* src = "crypto_accelerator.v:1036" *)
  wire _T_713;
  (* src = "crypto_accelerator.v:1037" *)
  wire _T_715;
  (* src = "crypto_accelerator.v:1038" *)
  wire _T_717;
  (* src = "crypto_accelerator.v:1039" *)
  wire _T_719;
  (* src = "crypto_accelerator.v:1040" *)
  wire _T_721;
  (* src = "crypto_accelerator.v:1041" *)
  wire _T_723;
  (* src = "crypto_accelerator.v:1042" *)
  wire _T_725;
  (* src = "crypto_accelerator.v:1043" *)
  wire _T_727;
  (* src = "crypto_accelerator.v:1044" *)
  wire _T_729;
  (* src = "crypto_accelerator.v:1045" *)
  wire _T_731;
  (* src = "crypto_accelerator.v:1046" *)
  wire _T_733;
  (* src = "crypto_accelerator.v:1047" *)
  wire _T_735;
  (* src = "crypto_accelerator.v:1048" *)
  wire _T_737;
  (* src = "crypto_accelerator.v:1049" *)
  wire _T_739;
  (* src = "crypto_accelerator.v:1050" *)
  wire _T_741;
  (* src = "crypto_accelerator.v:1051" *)
  wire _T_743;
  (* src = "crypto_accelerator.v:1052" *)
  wire _T_745;
  (* src = "crypto_accelerator.v:1053" *)
  wire _T_747;
  (* src = "crypto_accelerator.v:1054" *)
  wire _T_749;
  (* src = "crypto_accelerator.v:1055" *)
  wire _T_751;
  (* src = "crypto_accelerator.v:1056" *)
  wire _T_753;
  (* src = "crypto_accelerator.v:1057" *)
  wire _T_755;
  (* src = "crypto_accelerator.v:1058" *)
  wire _T_757;
  (* src = "crypto_accelerator.v:1059" *)
  wire _T_759;
  (* src = "crypto_accelerator.v:1060" *)
  wire _T_761;
  (* src = "crypto_accelerator.v:1061" *)
  wire _T_763;
  (* src = "crypto_accelerator.v:1062" *)
  wire _T_765;
  (* src = "crypto_accelerator.v:1063" *)
  wire _T_767;
  (* src = "crypto_accelerator.v:1064" *)
  wire _T_769;
  (* src = "crypto_accelerator.v:1065" *)
  wire _T_771;
  (* src = "crypto_accelerator.v:1066" *)
  wire _T_773;
  (* src = "crypto_accelerator.v:1067" *)
  wire _T_775;
  (* src = "crypto_accelerator.v:1068" *)
  wire _T_777;
  (* src = "crypto_accelerator.v:1069" *)
  wire _T_779;
  (* src = "crypto_accelerator.v:1070" *)
  wire _T_781;
  (* src = "crypto_accelerator.v:1071" *)
  wire _T_783;
  (* src = "crypto_accelerator.v:1072" *)
  wire _T_785;
  (* src = "crypto_accelerator.v:1073" *)
  wire _T_787;
  (* src = "crypto_accelerator.v:1074" *)
  wire _T_789;
  (* src = "crypto_accelerator.v:728" *)
  wire _T_79;
  (* src = "crypto_accelerator.v:1075" *)
  wire _T_791;
  (* src = "crypto_accelerator.v:1076" *)
  wire _T_793;
  (* src = "crypto_accelerator.v:1077" *)
  wire _T_795;
  (* src = "crypto_accelerator.v:1078" *)
  wire _T_797;
  (* src = "crypto_accelerator.v:1079" *)
  wire _T_799;
  (* src = "crypto_accelerator.v:1080" *)
  wire _T_801;
  (* src = "crypto_accelerator.v:1081" *)
  wire _T_803;
  (* src = "crypto_accelerator.v:1082" *)
  wire _T_805;
  (* src = "crypto_accelerator.v:1083" *)
  wire _T_807;
  (* src = "crypto_accelerator.v:1084" *)
  wire _T_809;
  (* src = "crypto_accelerator.v:729" *)
  wire _T_81;
  (* src = "crypto_accelerator.v:1085" *)
  wire _T_811;
  (* src = "crypto_accelerator.v:1086" *)
  wire _T_813;
  (* src = "crypto_accelerator.v:1087" *)
  wire _T_815;
  (* src = "crypto_accelerator.v:1088" *)
  wire _T_817;
  (* src = "crypto_accelerator.v:1089" *)
  wire _T_819;
  (* src = "crypto_accelerator.v:1090" *)
  wire _T_821;
  (* src = "crypto_accelerator.v:1091" *)
  wire _T_823;
  (* src = "crypto_accelerator.v:1092" *)
  wire _T_825;
  (* src = "crypto_accelerator.v:1093" *)
  wire _T_827;
  (* src = "crypto_accelerator.v:1094" *)
  wire _T_829;
  (* src = "crypto_accelerator.v:730" *)
  wire _T_83;
  (* src = "crypto_accelerator.v:1095" *)
  wire _T_831;
  (* src = "crypto_accelerator.v:1096" *)
  wire _T_833;
  (* src = "crypto_accelerator.v:1097" *)
  wire _T_834;
  (* src = "crypto_accelerator.v:1098" *)
  wire _T_835;
  (* src = "crypto_accelerator.v:1099" *)
  wire _T_836;
  (* src = "crypto_accelerator.v:1100" *)
  wire _T_838;
  (* src = "crypto_accelerator.v:1101" *)
  wire _T_839;
  (* src = "crypto_accelerator.v:1102" *)
  wire _T_840;
  (* src = "crypto_accelerator.v:1103" *)
  wire _T_842;
  (* src = "crypto_accelerator.v:1104" *)
  wire _T_844;
  (* src = "crypto_accelerator.v:1105" *)
  wire _T_845;
  (* src = "crypto_accelerator.v:1106" *)
  wire _T_846;
  (* src = "crypto_accelerator.v:1107" *)
  wire _T_848;
  (* src = "crypto_accelerator.v:731" *)
  wire _T_85;
  (* src = "crypto_accelerator.v:1108" *)
  wire _T_850;
  (* src = "crypto_accelerator.v:1109" *)
  wire _T_852;
  (* src = "crypto_accelerator.v:1110" *)
  wire _T_853;
  (* src = "crypto_accelerator.v:1111" *)
  wire _T_854;
  (* src = "crypto_accelerator.v:1112" *)
  wire _T_856;
  (* src = "crypto_accelerator.v:1113" *)
  wire _T_857;
  (* src = "crypto_accelerator.v:1114" *)
  wire _T_859;
  (* src = "crypto_accelerator.v:1115" *)
  wire _T_860;
  (* src = "crypto_accelerator.v:1116" *)
  wire _T_861;
  (* src = "crypto_accelerator.v:732" *)
  wire _T_87;
  (* src = "crypto_accelerator.v:1118" *)
  wire _T_886;
  (* src = "crypto_accelerator.v:1119" *)
  wire _T_888;
  (* src = "crypto_accelerator.v:733" *)
  wire _T_89;
  (* src = "crypto_accelerator.v:1120" *)
  wire _T_890;
  (* src = "crypto_accelerator.v:1121" *)
  wire _T_892;
  (* src = "crypto_accelerator.v:1122" *)
  wire _T_894;
  (* src = "crypto_accelerator.v:1123" *)
  wire _T_896;
  (* src = "crypto_accelerator.v:1124" *)
  wire _T_898;
  (* src = "crypto_accelerator.v:1125" *)
  wire _T_900;
  (* src = "crypto_accelerator.v:1126" *)
  wire _T_902;
  (* src = "crypto_accelerator.v:1127" *)
  wire _T_904;
  (* src = "crypto_accelerator.v:1128" *)
  wire _T_906;
  (* src = "crypto_accelerator.v:1129" *)
  wire _T_908;
  (* src = "crypto_accelerator.v:734" *)
  wire _T_91;
  (* src = "crypto_accelerator.v:1130" *)
  wire _T_910;
  (* src = "crypto_accelerator.v:1131" *)
  wire _T_912;
  (* src = "crypto_accelerator.v:1132" *)
  wire _T_914;
  (* src = "crypto_accelerator.v:1133" *)
  wire _T_916;
  (* src = "crypto_accelerator.v:1134" *)
  wire _T_918;
  (* src = "crypto_accelerator.v:1135" *)
  wire _T_920;
  (* src = "crypto_accelerator.v:1136" *)
  wire _T_922;
  (* src = "crypto_accelerator.v:1137" *)
  wire _T_924;
  (* src = "crypto_accelerator.v:1138" *)
  wire _T_926;
  (* src = "crypto_accelerator.v:1139" *)
  wire _T_928;
  (* src = "crypto_accelerator.v:735" *)
  wire _T_93;
  (* src = "crypto_accelerator.v:1140" *)
  wire _T_930;
  (* src = "crypto_accelerator.v:1141" *)
  wire _T_932;
  (* src = "crypto_accelerator.v:1142" *)
  wire _T_934;
  (* src = "crypto_accelerator.v:1143" *)
  wire _T_936;
  (* src = "crypto_accelerator.v:1144" *)
  wire _T_938;
  (* src = "crypto_accelerator.v:1145" *)
  wire _T_940;
  (* src = "crypto_accelerator.v:1146" *)
  wire _T_942;
  (* src = "crypto_accelerator.v:1147" *)
  wire _T_944;
  (* src = "crypto_accelerator.v:1148" *)
  wire _T_946;
  (* src = "crypto_accelerator.v:1149" *)
  wire _T_948;
  (* src = "crypto_accelerator.v:736" *)
  wire _T_95;
  (* src = "crypto_accelerator.v:1150" *)
  wire _T_950;
  (* src = "crypto_accelerator.v:1151" *)
  wire _T_952;
  (* src = "crypto_accelerator.v:1152" *)
  wire _T_954;
  (* src = "crypto_accelerator.v:1153" *)
  wire _T_956;
  (* src = "crypto_accelerator.v:1154" *)
  wire _T_958;
  (* src = "crypto_accelerator.v:1155" *)
  wire _T_960;
  (* src = "crypto_accelerator.v:1156" *)
  wire _T_962;
  (* src = "crypto_accelerator.v:1157" *)
  wire _T_964;
  (* src = "crypto_accelerator.v:1158" *)
  wire _T_966;
  (* src = "crypto_accelerator.v:1159" *)
  wire _T_968;
  (* src = "crypto_accelerator.v:737" *)
  wire _T_97;
  (* src = "crypto_accelerator.v:1160" *)
  wire _T_970;
  (* src = "crypto_accelerator.v:1161" *)
  wire _T_972;
  (* src = "crypto_accelerator.v:1162" *)
  wire _T_974;
  (* src = "crypto_accelerator.v:1163" *)
  wire _T_976;
  (* src = "crypto_accelerator.v:1164" *)
  wire _T_978;
  (* src = "crypto_accelerator.v:1165" *)
  wire _T_980;
  (* src = "crypto_accelerator.v:1166" *)
  wire _T_982;
  (* src = "crypto_accelerator.v:1167" *)
  wire _T_984;
  (* src = "crypto_accelerator.v:1168" *)
  wire _T_986;
  (* src = "crypto_accelerator.v:1169" *)
  wire _T_988;
  (* src = "crypto_accelerator.v:738" *)
  wire _T_99;
  (* src = "crypto_accelerator.v:1170" *)
  wire _T_990;
  (* src = "crypto_accelerator.v:1171" *)
  wire _T_992;
  (* src = "crypto_accelerator.v:1172" *)
  wire _T_994;
  (* src = "crypto_accelerator.v:1173" *)
  wire _T_996;
  (* src = "crypto_accelerator.v:1174" *)
  wire _T_998;
  (* src = "crypto_accelerator.v:604" *)
  input clock;
  (* src = "crypto_accelerator.v:712" *)
  wire [7:0] initOut_0_0;
  (* src = "crypto_accelerator.v:713" *)
  wire [7:0] initOut_0_1;
  (* src = "crypto_accelerator.v:714" *)
  wire [7:0] initOut_0_2;
  (* src = "crypto_accelerator.v:715" *)
  wire [7:0] initOut_0_3;
  (* src = "crypto_accelerator.v:716" *)
  wire [7:0] initOut_1_0;
  (* src = "crypto_accelerator.v:717" *)
  wire [7:0] initOut_1_1;
  (* src = "crypto_accelerator.v:718" *)
  wire [7:0] initOut_1_2;
  (* src = "crypto_accelerator.v:719" *)
  wire [7:0] initOut_1_3;
  (* src = "crypto_accelerator.v:720" *)
  wire [7:0] initOut_2_0;
  (* src = "crypto_accelerator.v:721" *)
  wire [7:0] initOut_2_1;
  (* src = "crypto_accelerator.v:722" *)
  wire [7:0] initOut_2_2;
  (* src = "crypto_accelerator.v:723" *)
  wire [7:0] initOut_2_3;
  (* src = "crypto_accelerator.v:724" *)
  wire [7:0] initOut_3_0;
  (* src = "crypto_accelerator.v:725" *)
  wire [7:0] initOut_3_1;
  (* src = "crypto_accelerator.v:726" *)
  wire [7:0] initOut_3_2;
  (* src = "crypto_accelerator.v:727" *)
  wire [7:0] initOut_3_3;
  (* src = "crypto_accelerator.v:625" *)
  input io_aes256;
  (* src = "crypto_accelerator.v:606" *)
  input [127:0] io_dataIn;
  (* src = "crypto_accelerator.v:629" *)
  output [127:0] io_dataOut;
  (* src = "crypto_accelerator.v:608" *)
  input io_dataValid;
  (* src = "crypto_accelerator.v:607" *)
  input [127:0] io_ivIn;
  (* src = "crypto_accelerator.v:630" *)
  output [127:0] io_ivOut;
  (* src = "crypto_accelerator.v:609" *)
  input [7:0] io_keys_0_0_0;
  (* src = "crypto_accelerator.v:610" *)
  input [7:0] io_keys_0_0_1;
  (* src = "crypto_accelerator.v:611" *)
  input [7:0] io_keys_0_0_2;
  (* src = "crypto_accelerator.v:612" *)
  input [7:0] io_keys_0_0_3;
  (* src = "crypto_accelerator.v:613" *)
  input [7:0] io_keys_0_1_0;
  (* src = "crypto_accelerator.v:614" *)
  input [7:0] io_keys_0_1_1;
  (* src = "crypto_accelerator.v:615" *)
  input [7:0] io_keys_0_1_2;
  (* src = "crypto_accelerator.v:616" *)
  input [7:0] io_keys_0_1_3;
  (* src = "crypto_accelerator.v:617" *)
  input [7:0] io_keys_0_2_0;
  (* src = "crypto_accelerator.v:618" *)
  input [7:0] io_keys_0_2_1;
  (* src = "crypto_accelerator.v:619" *)
  input [7:0] io_keys_0_2_2;
  (* src = "crypto_accelerator.v:620" *)
  input [7:0] io_keys_0_2_3;
  (* src = "crypto_accelerator.v:621" *)
  input [7:0] io_keys_0_3_0;
  (* src = "crypto_accelerator.v:622" *)
  input [7:0] io_keys_0_3_1;
  (* src = "crypto_accelerator.v:623" *)
  input [7:0] io_keys_0_3_2;
  (* src = "crypto_accelerator.v:624" *)
  input [7:0] io_keys_0_3_3;
  (* src = "crypto_accelerator.v:631" *)
  output io_outputValid;
  (* src = "crypto_accelerator.v:628" *)
  output io_ready;
  (* src = "crypto_accelerator.v:627" *)
  output io_shift;
  (* src = "crypto_accelerator.v:626" *)
  output io_shiftCyc;
  (* src = "crypto_accelerator.v:690" *)
  reg [7:0] matrix_0_0;
  (* src = "crypto_accelerator.v:691" *)
  reg [7:0] matrix_0_1;
  (* src = "crypto_accelerator.v:692" *)
  reg [7:0] matrix_0_2;
  (* src = "crypto_accelerator.v:693" *)
  reg [7:0] matrix_0_3;
  (* src = "crypto_accelerator.v:694" *)
  reg [7:0] matrix_1_0;
  (* src = "crypto_accelerator.v:695" *)
  reg [7:0] matrix_1_1;
  (* src = "crypto_accelerator.v:696" *)
  reg [7:0] matrix_1_2;
  (* src = "crypto_accelerator.v:697" *)
  reg [7:0] matrix_1_3;
  (* src = "crypto_accelerator.v:698" *)
  reg [7:0] matrix_2_0;
  (* src = "crypto_accelerator.v:699" *)
  reg [7:0] matrix_2_1;
  (* src = "crypto_accelerator.v:700" *)
  reg [7:0] matrix_2_2;
  (* src = "crypto_accelerator.v:701" *)
  reg [7:0] matrix_2_3;
  (* src = "crypto_accelerator.v:702" *)
  reg [7:0] matrix_3_0;
  (* src = "crypto_accelerator.v:703" *)
  reg [7:0] matrix_3_1;
  (* src = "crypto_accelerator.v:704" *)
  reg [7:0] matrix_3_2;
  (* src = "crypto_accelerator.v:705" *)
  reg [7:0] matrix_3_3;
  (* src = "crypto_accelerator.v:605" *)
  input reset;
  (* src = "crypto_accelerator.v:857" *)
  wire [7:0] roundPart1_0_0;
  (* src = "crypto_accelerator.v:1507" *)
  wire [7:0] roundPart1_0_1;
  (* src = "crypto_accelerator.v:2157" *)
  wire [7:0] roundPart1_0_2;
  (* src = "crypto_accelerator.v:2807" *)
  wire [7:0] roundPart1_0_3;
  (* src = "crypto_accelerator.v:1377" *)
  wire [7:0] roundPart1_1_0;
  (* src = "crypto_accelerator.v:2027" *)
  wire [7:0] roundPart1_1_1;
  (* src = "crypto_accelerator.v:2677" *)
  wire [7:0] roundPart1_1_2;
  (* src = "crypto_accelerator.v:1247" *)
  wire [7:0] roundPart1_1_3;
  (* src = "crypto_accelerator.v:1897" *)
  wire [7:0] roundPart1_2_0;
  (* src = "crypto_accelerator.v:2547" *)
  wire [7:0] roundPart1_2_1;
  (* src = "crypto_accelerator.v:1117" *)
  wire [7:0] roundPart1_2_2;
  (* src = "crypto_accelerator.v:1767" *)
  wire [7:0] roundPart1_2_3;
  (* src = "crypto_accelerator.v:2417" *)
  wire [7:0] roundPart1_3_0;
  (* src = "crypto_accelerator.v:987" *)
  wire [7:0] roundPart1_3_1;
  (* src = "crypto_accelerator.v:1637" *)
  wire [7:0] roundPart1_3_2;
  (* src = "crypto_accelerator.v:2287" *)
  wire [7:0] roundPart1_3_3;
  (* src = "crypto_accelerator.v:2808" *)
  wire [7:0] roundPart2_0_0;
  (* src = "crypto_accelerator.v:2809" *)
  wire [7:0] roundPart2_0_1;
  (* src = "crypto_accelerator.v:2810" *)
  wire [7:0] roundPart2_0_2;
  (* src = "crypto_accelerator.v:2811" *)
  wire [7:0] roundPart2_0_3;
  (* src = "crypto_accelerator.v:2812" *)
  wire [7:0] roundPart2_1_0;
  (* src = "crypto_accelerator.v:2813" *)
  wire [7:0] roundPart2_1_1;
  (* src = "crypto_accelerator.v:2814" *)
  wire [7:0] roundPart2_1_2;
  (* src = "crypto_accelerator.v:2815" *)
  wire [7:0] roundPart2_1_3;
  (* src = "crypto_accelerator.v:2816" *)
  wire [7:0] roundPart2_2_0;
  (* src = "crypto_accelerator.v:2817" *)
  wire [7:0] roundPart2_2_1;
  (* src = "crypto_accelerator.v:2818" *)
  wire [7:0] roundPart2_2_2;
  (* src = "crypto_accelerator.v:2819" *)
  wire [7:0] roundPart2_2_3;
  (* src = "crypto_accelerator.v:2820" *)
  wire [7:0] roundPart2_3_0;
  (* src = "crypto_accelerator.v:2821" *)
  wire [7:0] roundPart2_3_1;
  (* src = "crypto_accelerator.v:2822" *)
  wire [7:0] roundPart2_3_2;
  (* src = "crypto_accelerator.v:2823" *)
  wire [7:0] roundPart2_3_3;
  (* src = "crypto_accelerator.v:2824" *)
  wire [7:0] roundPart2_last_0_0;
  (* src = "crypto_accelerator.v:2825" *)
  wire [7:0] roundPart2_last_0_1;
  (* src = "crypto_accelerator.v:2826" *)
  wire [7:0] roundPart2_last_0_2;
  (* src = "crypto_accelerator.v:2827" *)
  wire [7:0] roundPart2_last_0_3;
  (* src = "crypto_accelerator.v:2828" *)
  wire [7:0] roundPart2_last_1_0;
  (* src = "crypto_accelerator.v:2829" *)
  wire [7:0] roundPart2_last_1_1;
  (* src = "crypto_accelerator.v:2830" *)
  wire [7:0] roundPart2_last_1_2;
  (* src = "crypto_accelerator.v:2831" *)
  wire [7:0] roundPart2_last_1_3;
  (* src = "crypto_accelerator.v:2832" *)
  wire [7:0] roundPart2_last_2_0;
  (* src = "crypto_accelerator.v:2833" *)
  wire [7:0] roundPart2_last_2_1;
  (* src = "crypto_accelerator.v:2834" *)
  wire [7:0] roundPart2_last_2_2;
  (* src = "crypto_accelerator.v:2835" *)
  wire [7:0] roundPart2_last_2_3;
  (* src = "crypto_accelerator.v:2836" *)
  wire [7:0] roundPart2_last_3_0;
  (* src = "crypto_accelerator.v:2837" *)
  wire [7:0] roundPart2_last_3_1;
  (* src = "crypto_accelerator.v:2838" *)
  wire [7:0] roundPart2_last_3_2;
  (* src = "crypto_accelerator.v:2839" *)
  wire [7:0] roundPart2_last_3_3;
  (* src = "crypto_accelerator.v:684" *)
  reg [5:0] state;
  assign _T_4427 = state + (* src = "crypto_accelerator.v:2846" *) 1'b1;
  assign _T_671 = _T_653 & (* src = "crypto_accelerator.v:1015" *) _T_625;
  assign _T_673 = _T_655 & (* src = "crypto_accelerator.v:1016" *) _T_637;
  assign _T_677 = _T_635 & (* src = "crypto_accelerator.v:1018" *) matrix_0_2[0];
  assign _T_681 = _T_629 & (* src = "crypto_accelerator.v:1020" *) _T_657;
  assign _T_683 = _T_633 & (* src = "crypto_accelerator.v:1021" *) _T_623;
  assign _T_687 = _T_659 & (* src = "crypto_accelerator.v:1023" *) _T_649;
  assign _T_691 = _T_619 & (* src = "crypto_accelerator.v:1025" *) _T_631;
  assign _T_693 = _T_665 & (* src = "crypto_accelerator.v:1026" *) _T_661;
  assign _T_697 = _T_647 & (* src = "crypto_accelerator.v:1028" *) _T_643;
  assign _T_719 = _T_713 & (* src = "crypto_accelerator.v:1039" *) _T_709;
  assign _T_727 = _T_725 & (* src = "crypto_accelerator.v:1043" *) _T_723;
  assign _T_729 = _T_721 & (* src = "crypto_accelerator.v:1044" *) _T_717;
  assign _T_731 = _T_709 & (* src = "crypto_accelerator.v:1045" *) _T_715;
  assign _T_733 = _T_723 & (* src = "crypto_accelerator.v:1046" *) _T_731;
  assign _T_737 = _T_711 & (* src = "crypto_accelerator.v:1048" *) _T_713;
  assign _T_739 = _T_717 & (* src = "crypto_accelerator.v:1049" *) _T_737;
  assign _T_761 = _T_757 & (* src = "crypto_accelerator.v:1060" *) _T_625;
  assign _T_763 = _T_749 & (* src = "crypto_accelerator.v:1061" *) _T_637;
  assign _T_765 = _T_747 & (* src = "crypto_accelerator.v:1062" *) matrix_0_2[0];
  assign _T_767 = _T_755 & (* src = "crypto_accelerator.v:1063" *) _T_657;
  assign _T_769 = _T_745 & (* src = "crypto_accelerator.v:1064" *) _T_623;
  assign _T_771 = _T_743 & (* src = "crypto_accelerator.v:1065" *) _T_649;
  assign _T_773 = _T_753 & (* src = "crypto_accelerator.v:1066" *) _T_631;
  assign _T_775 = _T_759 & (* src = "crypto_accelerator.v:1067" *) _T_661;
  assign _T_777 = _T_751 & (* src = "crypto_accelerator.v:1068" *) _T_643;
  assign _T_779 = _T_757 & (* src = "crypto_accelerator.v:1069" *) _T_653;
  assign _T_781 = _T_749 & (* src = "crypto_accelerator.v:1070" *) _T_655;
  assign _T_783 = _T_747 & (* src = "crypto_accelerator.v:1071" *) _T_635;
  assign _T_785 = _T_755 & (* src = "crypto_accelerator.v:1072" *) _T_629;
  assign _T_787 = _T_745 & (* src = "crypto_accelerator.v:1073" *) _T_633;
  assign _T_789 = _T_743 & (* src = "crypto_accelerator.v:1074" *) _T_659;
  assign _T_791 = _T_753 & (* src = "crypto_accelerator.v:1075" *) _T_619;
  assign _T_793 = _T_759 & (* src = "crypto_accelerator.v:1076" *) _T_665;
  assign _T_795 = _T_751 & (* src = "crypto_accelerator.v:1077" *) _T_647;
  assign _T_940 = _T_922 & (* src = "crypto_accelerator.v:1145" *) _T_894;
  assign _T_942 = _T_924 & (* src = "crypto_accelerator.v:1146" *) _T_906;
  assign _T_946 = _T_904 & (* src = "crypto_accelerator.v:1148" *) matrix_0_3[0];
  assign _T_950 = _T_898 & (* src = "crypto_accelerator.v:1150" *) _T_926;
  assign _T_952 = _T_902 & (* src = "crypto_accelerator.v:1151" *) _T_892;
  assign _T_956 = _T_928 & (* src = "crypto_accelerator.v:1153" *) _T_918;
  assign _T_960 = _T_888 & (* src = "crypto_accelerator.v:1155" *) _T_900;
  assign _T_962 = _T_934 & (* src = "crypto_accelerator.v:1156" *) _T_930;
  assign _T_966 = _T_916 & (* src = "crypto_accelerator.v:1158" *) _T_912;
  assign _T_988 = _T_982 & (* src = "crypto_accelerator.v:1169" *) _T_978;
  assign _T_996 = _T_994 & (* src = "crypto_accelerator.v:1173" *) _T_992;
  assign _T_998 = _T_990 & (* src = "crypto_accelerator.v:1174" *) _T_986;
  assign _T_1000 = _T_978 & (* src = "crypto_accelerator.v:1175" *) _T_984;
  assign _T_1002 = _T_992 & (* src = "crypto_accelerator.v:1176" *) _T_1000;
  assign _T_1006 = _T_980 & (* src = "crypto_accelerator.v:1178" *) _T_982;
  assign _T_1008 = _T_986 & (* src = "crypto_accelerator.v:1179" *) _T_1006;
  assign _T_1030 = _T_1026 & (* src = "crypto_accelerator.v:1190" *) _T_894;
  assign _T_1032 = _T_1018 & (* src = "crypto_accelerator.v:1191" *) _T_906;
  assign _T_1034 = _T_1016 & (* src = "crypto_accelerator.v:1192" *) matrix_0_3[0];
  assign _T_1036 = _T_1024 & (* src = "crypto_accelerator.v:1193" *) _T_926;
  assign _T_1038 = _T_1014 & (* src = "crypto_accelerator.v:1194" *) _T_892;
  assign _T_1040 = _T_1012 & (* src = "crypto_accelerator.v:1195" *) _T_918;
  assign _T_1042 = _T_1022 & (* src = "crypto_accelerator.v:1196" *) _T_900;
  assign _T_1044 = _T_1028 & (* src = "crypto_accelerator.v:1197" *) _T_930;
  assign _T_1046 = _T_1020 & (* src = "crypto_accelerator.v:1198" *) _T_912;
  assign _T_1048 = _T_1026 & (* src = "crypto_accelerator.v:1199" *) _T_922;
  assign _T_1050 = _T_1018 & (* src = "crypto_accelerator.v:1200" *) _T_924;
  assign _T_1052 = _T_1016 & (* src = "crypto_accelerator.v:1201" *) _T_904;
  assign _T_1054 = _T_1024 & (* src = "crypto_accelerator.v:1202" *) _T_898;
  assign _T_1056 = _T_1014 & (* src = "crypto_accelerator.v:1203" *) _T_902;
  assign _T_1058 = _T_1012 & (* src = "crypto_accelerator.v:1204" *) _T_928;
  assign _T_1060 = _T_1022 & (* src = "crypto_accelerator.v:1205" *) _T_888;
  assign _T_1062 = _T_1028 & (* src = "crypto_accelerator.v:1206" *) _T_934;
  assign _T_1064 = _T_1020 & (* src = "crypto_accelerator.v:1207" *) _T_916;
  assign _T_1210 = _T_1192 & (* src = "crypto_accelerator.v:1275" *) _T_1164;
  assign _T_1212 = _T_1194 & (* src = "crypto_accelerator.v:1276" *) _T_1176;
  assign _T_1216 = _T_1174 & (* src = "crypto_accelerator.v:1278" *) matrix_1_0[0];
  assign _T_1220 = _T_1168 & (* src = "crypto_accelerator.v:1280" *) _T_1196;
  assign _T_1222 = _T_1172 & (* src = "crypto_accelerator.v:1281" *) _T_1162;
  assign _T_1226 = _T_1198 & (* src = "crypto_accelerator.v:1283" *) _T_1188;
  assign _T_1230 = _T_1158 & (* src = "crypto_accelerator.v:1285" *) _T_1170;
  assign _T_1232 = _T_1204 & (* src = "crypto_accelerator.v:1286" *) _T_1200;
  assign _T_1236 = _T_1186 & (* src = "crypto_accelerator.v:1288" *) _T_1182;
  assign _T_1258 = _T_1252 & (* src = "crypto_accelerator.v:1299" *) _T_1248;
  assign _T_1266 = _T_1264 & (* src = "crypto_accelerator.v:1303" *) _T_1262;
  assign _T_1268 = _T_1260 & (* src = "crypto_accelerator.v:1304" *) _T_1256;
  assign _T_1270 = _T_1248 & (* src = "crypto_accelerator.v:1305" *) _T_1254;
  assign _T_1272 = _T_1262 & (* src = "crypto_accelerator.v:1306" *) _T_1270;
  assign _T_1276 = _T_1250 & (* src = "crypto_accelerator.v:1308" *) _T_1252;
  assign _T_1278 = _T_1256 & (* src = "crypto_accelerator.v:1309" *) _T_1276;
  assign _T_1300 = _T_1296 & (* src = "crypto_accelerator.v:1320" *) _T_1164;
  assign _T_1302 = _T_1288 & (* src = "crypto_accelerator.v:1321" *) _T_1176;
  assign _T_1304 = _T_1286 & (* src = "crypto_accelerator.v:1322" *) matrix_1_0[0];
  assign _T_1306 = _T_1294 & (* src = "crypto_accelerator.v:1323" *) _T_1196;
  assign _T_1308 = _T_1284 & (* src = "crypto_accelerator.v:1324" *) _T_1162;
  assign _T_1310 = _T_1282 & (* src = "crypto_accelerator.v:1325" *) _T_1188;
  assign _T_1312 = _T_1292 & (* src = "crypto_accelerator.v:1326" *) _T_1170;
  assign _T_1314 = _T_1298 & (* src = "crypto_accelerator.v:1327" *) _T_1200;
  assign _T_1316 = _T_1290 & (* src = "crypto_accelerator.v:1328" *) _T_1182;
  assign _T_1318 = _T_1296 & (* src = "crypto_accelerator.v:1329" *) _T_1192;
  assign _T_1320 = _T_1288 & (* src = "crypto_accelerator.v:1330" *) _T_1194;
  assign _T_1322 = _T_1286 & (* src = "crypto_accelerator.v:1331" *) _T_1174;
  assign _T_1324 = _T_1294 & (* src = "crypto_accelerator.v:1332" *) _T_1168;
  assign _T_1326 = _T_1284 & (* src = "crypto_accelerator.v:1333" *) _T_1172;
  assign _T_1328 = _T_1282 & (* src = "crypto_accelerator.v:1334" *) _T_1198;
  assign _T_1330 = _T_1292 & (* src = "crypto_accelerator.v:1335" *) _T_1158;
  assign _T_1332 = _T_1298 & (* src = "crypto_accelerator.v:1336" *) _T_1204;
  assign _T_1334 = _T_1290 & (* src = "crypto_accelerator.v:1337" *) _T_1186;
  assign _T_1479 = _T_1461 & (* src = "crypto_accelerator.v:1405" *) _T_1433;
  assign _T_1481 = _T_1463 & (* src = "crypto_accelerator.v:1406" *) _T_1445;
  assign _T_1485 = _T_1443 & (* src = "crypto_accelerator.v:1408" *) matrix_1_1[0];
  assign _T_1489 = _T_1437 & (* src = "crypto_accelerator.v:1410" *) _T_1465;
  assign _T_1491 = _T_1441 & (* src = "crypto_accelerator.v:1411" *) _T_1431;
  assign _T_1495 = _T_1467 & (* src = "crypto_accelerator.v:1413" *) _T_1457;
  assign _T_1499 = _T_1427 & (* src = "crypto_accelerator.v:1415" *) _T_1439;
  assign _T_1501 = _T_1473 & (* src = "crypto_accelerator.v:1416" *) _T_1469;
  assign _T_1505 = _T_1455 & (* src = "crypto_accelerator.v:1418" *) _T_1451;
  assign _T_1527 = _T_1521 & (* src = "crypto_accelerator.v:1429" *) _T_1517;
  assign _T_1535 = _T_1533 & (* src = "crypto_accelerator.v:1433" *) _T_1531;
  assign _T_1537 = _T_1529 & (* src = "crypto_accelerator.v:1434" *) _T_1525;
  assign _T_1539 = _T_1517 & (* src = "crypto_accelerator.v:1435" *) _T_1523;
  assign _T_1541 = _T_1531 & (* src = "crypto_accelerator.v:1436" *) _T_1539;
  assign _T_1545 = _T_1519 & (* src = "crypto_accelerator.v:1438" *) _T_1521;
  assign _T_1547 = _T_1525 & (* src = "crypto_accelerator.v:1439" *) _T_1545;
  assign _T_1569 = _T_1565 & (* src = "crypto_accelerator.v:1450" *) _T_1433;
  assign _T_1571 = _T_1557 & (* src = "crypto_accelerator.v:1451" *) _T_1445;
  assign _T_1573 = _T_1555 & (* src = "crypto_accelerator.v:1452" *) matrix_1_1[0];
  assign _T_1575 = _T_1563 & (* src = "crypto_accelerator.v:1453" *) _T_1465;
  assign _T_1577 = _T_1553 & (* src = "crypto_accelerator.v:1454" *) _T_1431;
  assign _T_1579 = _T_1551 & (* src = "crypto_accelerator.v:1455" *) _T_1457;
  assign _T_1581 = _T_1561 & (* src = "crypto_accelerator.v:1456" *) _T_1439;
  assign _T_1583 = _T_1567 & (* src = "crypto_accelerator.v:1457" *) _T_1469;
  assign _T_1585 = _T_1559 & (* src = "crypto_accelerator.v:1458" *) _T_1451;
  assign _T_1587 = _T_1565 & (* src = "crypto_accelerator.v:1459" *) _T_1461;
  assign _T_1589 = _T_1557 & (* src = "crypto_accelerator.v:1460" *) _T_1463;
  assign _T_1591 = _T_1555 & (* src = "crypto_accelerator.v:1461" *) _T_1443;
  assign _T_1593 = _T_1563 & (* src = "crypto_accelerator.v:1462" *) _T_1437;
  assign _T_1595 = _T_1553 & (* src = "crypto_accelerator.v:1463" *) _T_1441;
  assign _T_1597 = _T_1551 & (* src = "crypto_accelerator.v:1464" *) _T_1467;
  assign _T_1599 = _T_1561 & (* src = "crypto_accelerator.v:1465" *) _T_1427;
  assign _T_1601 = _T_1567 & (* src = "crypto_accelerator.v:1466" *) _T_1473;
  assign _T_1603 = _T_1559 & (* src = "crypto_accelerator.v:1467" *) _T_1455;
  assign _T_1748 = _T_1730 & (* src = "crypto_accelerator.v:1535" *) _T_1702;
  assign _T_1750 = _T_1732 & (* src = "crypto_accelerator.v:1536" *) _T_1714;
  assign _T_1754 = _T_1712 & (* src = "crypto_accelerator.v:1538" *) matrix_1_2[0];
  assign _T_1758 = _T_1706 & (* src = "crypto_accelerator.v:1540" *) _T_1734;
  assign _T_1760 = _T_1710 & (* src = "crypto_accelerator.v:1541" *) _T_1700;
  assign _T_1764 = _T_1736 & (* src = "crypto_accelerator.v:1543" *) _T_1726;
  assign _T_1768 = _T_1696 & (* src = "crypto_accelerator.v:1545" *) _T_1708;
  assign _T_1770 = _T_1742 & (* src = "crypto_accelerator.v:1546" *) _T_1738;
  assign _T_1774 = _T_1724 & (* src = "crypto_accelerator.v:1548" *) _T_1720;
  assign _T_1796 = _T_1790 & (* src = "crypto_accelerator.v:1559" *) _T_1786;
  assign _T_1804 = _T_1802 & (* src = "crypto_accelerator.v:1563" *) _T_1800;
  assign _T_1806 = _T_1798 & (* src = "crypto_accelerator.v:1564" *) _T_1794;
  assign _T_1808 = _T_1786 & (* src = "crypto_accelerator.v:1565" *) _T_1792;
  assign _T_1810 = _T_1800 & (* src = "crypto_accelerator.v:1566" *) _T_1808;
  assign _T_1814 = _T_1788 & (* src = "crypto_accelerator.v:1568" *) _T_1790;
  assign _T_1816 = _T_1794 & (* src = "crypto_accelerator.v:1569" *) _T_1814;
  assign _T_1838 = _T_1834 & (* src = "crypto_accelerator.v:1580" *) _T_1702;
  assign _T_1840 = _T_1826 & (* src = "crypto_accelerator.v:1581" *) _T_1714;
  assign _T_1842 = _T_1824 & (* src = "crypto_accelerator.v:1582" *) matrix_1_2[0];
  assign _T_1844 = _T_1832 & (* src = "crypto_accelerator.v:1583" *) _T_1734;
  assign _T_1846 = _T_1822 & (* src = "crypto_accelerator.v:1584" *) _T_1700;
  assign _T_1848 = _T_1820 & (* src = "crypto_accelerator.v:1585" *) _T_1726;
  assign _T_1850 = _T_1830 & (* src = "crypto_accelerator.v:1586" *) _T_1708;
  assign _T_1852 = _T_1836 & (* src = "crypto_accelerator.v:1587" *) _T_1738;
  assign _T_1854 = _T_1828 & (* src = "crypto_accelerator.v:1588" *) _T_1720;
  assign _T_1856 = _T_1834 & (* src = "crypto_accelerator.v:1589" *) _T_1730;
  assign _T_1858 = _T_1826 & (* src = "crypto_accelerator.v:1590" *) _T_1732;
  assign _T_1860 = _T_1824 & (* src = "crypto_accelerator.v:1591" *) _T_1712;
  assign _T_1862 = _T_1832 & (* src = "crypto_accelerator.v:1592" *) _T_1706;
  assign _T_1864 = _T_1822 & (* src = "crypto_accelerator.v:1593" *) _T_1710;
  assign _T_1866 = _T_1820 & (* src = "crypto_accelerator.v:1594" *) _T_1736;
  assign _T_1868 = _T_1830 & (* src = "crypto_accelerator.v:1595" *) _T_1696;
  assign _T_1870 = _T_1836 & (* src = "crypto_accelerator.v:1596" *) _T_1742;
  assign _T_1872 = _T_1828 & (* src = "crypto_accelerator.v:1597" *) _T_1724;
  assign _T_2017 = _T_1999 & (* src = "crypto_accelerator.v:1665" *) _T_1971;
  assign _T_2019 = _T_2001 & (* src = "crypto_accelerator.v:1666" *) _T_1983;
  assign _T_2023 = _T_1981 & (* src = "crypto_accelerator.v:1668" *) matrix_1_3[0];
  assign _T_2027 = _T_1975 & (* src = "crypto_accelerator.v:1670" *) _T_2003;
  assign _T_2029 = _T_1979 & (* src = "crypto_accelerator.v:1671" *) _T_1969;
  assign _T_2033 = _T_2005 & (* src = "crypto_accelerator.v:1673" *) _T_1995;
  assign _T_2037 = _T_1965 & (* src = "crypto_accelerator.v:1675" *) _T_1977;
  assign _T_2039 = _T_2011 & (* src = "crypto_accelerator.v:1676" *) _T_2007;
  assign _T_2043 = _T_1993 & (* src = "crypto_accelerator.v:1678" *) _T_1989;
  assign _T_2065 = _T_2059 & (* src = "crypto_accelerator.v:1689" *) _T_2055;
  assign _T_2073 = _T_2071 & (* src = "crypto_accelerator.v:1693" *) _T_2069;
  assign _T_2075 = _T_2067 & (* src = "crypto_accelerator.v:1694" *) _T_2063;
  assign _T_2077 = _T_2055 & (* src = "crypto_accelerator.v:1695" *) _T_2061;
  assign _T_2079 = _T_2069 & (* src = "crypto_accelerator.v:1696" *) _T_2077;
  assign _T_2083 = _T_2057 & (* src = "crypto_accelerator.v:1698" *) _T_2059;
  assign _T_2085 = _T_2063 & (* src = "crypto_accelerator.v:1699" *) _T_2083;
  assign _T_2107 = _T_2103 & (* src = "crypto_accelerator.v:1710" *) _T_1971;
  assign _T_2109 = _T_2095 & (* src = "crypto_accelerator.v:1711" *) _T_1983;
  assign _T_2111 = _T_2093 & (* src = "crypto_accelerator.v:1712" *) matrix_1_3[0];
  assign _T_2113 = _T_2101 & (* src = "crypto_accelerator.v:1713" *) _T_2003;
  assign _T_2115 = _T_2091 & (* src = "crypto_accelerator.v:1714" *) _T_1969;
  assign _T_2117 = _T_2089 & (* src = "crypto_accelerator.v:1715" *) _T_1995;
  assign _T_2119 = _T_2099 & (* src = "crypto_accelerator.v:1716" *) _T_1977;
  assign _T_2121 = _T_2105 & (* src = "crypto_accelerator.v:1717" *) _T_2007;
  assign _T_2123 = _T_2097 & (* src = "crypto_accelerator.v:1718" *) _T_1989;
  assign _T_2125 = _T_2103 & (* src = "crypto_accelerator.v:1719" *) _T_1999;
  assign _T_2127 = _T_2095 & (* src = "crypto_accelerator.v:1720" *) _T_2001;
  assign _T_2129 = _T_2093 & (* src = "crypto_accelerator.v:1721" *) _T_1981;
  assign _T_2131 = _T_2101 & (* src = "crypto_accelerator.v:1722" *) _T_1975;
  assign _T_2133 = _T_2091 & (* src = "crypto_accelerator.v:1723" *) _T_1979;
  assign _T_2135 = _T_2089 & (* src = "crypto_accelerator.v:1724" *) _T_2005;
  assign _T_2137 = _T_2099 & (* src = "crypto_accelerator.v:1725" *) _T_1965;
  assign _T_2139 = _T_2105 & (* src = "crypto_accelerator.v:1726" *) _T_2011;
  assign _T_2141 = _T_2097 & (* src = "crypto_accelerator.v:1727" *) _T_1993;
  assign _T_2287 = _T_2269 & (* src = "crypto_accelerator.v:1795" *) _T_2241;
  assign _T_2289 = _T_2271 & (* src = "crypto_accelerator.v:1796" *) _T_2253;
  assign _T_2293 = _T_2251 & (* src = "crypto_accelerator.v:1798" *) matrix_2_0[0];
  assign _T_2297 = _T_2245 & (* src = "crypto_accelerator.v:1800" *) _T_2273;
  assign _T_2299 = _T_2249 & (* src = "crypto_accelerator.v:1801" *) _T_2239;
  assign _T_2303 = _T_2275 & (* src = "crypto_accelerator.v:1803" *) _T_2265;
  assign _T_2307 = _T_2235 & (* src = "crypto_accelerator.v:1805" *) _T_2247;
  assign _T_2309 = _T_2281 & (* src = "crypto_accelerator.v:1806" *) _T_2277;
  assign _T_2313 = _T_2263 & (* src = "crypto_accelerator.v:1808" *) _T_2259;
  assign _T_2335 = _T_2329 & (* src = "crypto_accelerator.v:1819" *) _T_2325;
  assign _T_2343 = _T_2341 & (* src = "crypto_accelerator.v:1823" *) _T_2339;
  assign _T_2345 = _T_2337 & (* src = "crypto_accelerator.v:1824" *) _T_2333;
  assign _T_2347 = _T_2325 & (* src = "crypto_accelerator.v:1825" *) _T_2331;
  assign _T_2349 = _T_2339 & (* src = "crypto_accelerator.v:1826" *) _T_2347;
  assign _T_2353 = _T_2327 & (* src = "crypto_accelerator.v:1828" *) _T_2329;
  assign _T_2355 = _T_2333 & (* src = "crypto_accelerator.v:1829" *) _T_2353;
  assign _T_2377 = _T_2373 & (* src = "crypto_accelerator.v:1840" *) _T_2241;
  assign _T_2379 = _T_2365 & (* src = "crypto_accelerator.v:1841" *) _T_2253;
  assign _T_2381 = _T_2363 & (* src = "crypto_accelerator.v:1842" *) matrix_2_0[0];
  assign _T_2383 = _T_2371 & (* src = "crypto_accelerator.v:1843" *) _T_2273;
  assign _T_2385 = _T_2361 & (* src = "crypto_accelerator.v:1844" *) _T_2239;
  assign _T_2387 = _T_2359 & (* src = "crypto_accelerator.v:1845" *) _T_2265;
  assign _T_2389 = _T_2369 & (* src = "crypto_accelerator.v:1846" *) _T_2247;
  assign _T_2391 = _T_2375 & (* src = "crypto_accelerator.v:1847" *) _T_2277;
  assign _T_2393 = _T_2367 & (* src = "crypto_accelerator.v:1848" *) _T_2259;
  assign _T_2395 = _T_2373 & (* src = "crypto_accelerator.v:1849" *) _T_2269;
  assign _T_2397 = _T_2365 & (* src = "crypto_accelerator.v:1850" *) _T_2271;
  assign _T_2399 = _T_2363 & (* src = "crypto_accelerator.v:1851" *) _T_2251;
  assign _T_2401 = _T_2371 & (* src = "crypto_accelerator.v:1852" *) _T_2245;
  assign _T_2403 = _T_2361 & (* src = "crypto_accelerator.v:1853" *) _T_2249;
  assign _T_2405 = _T_2359 & (* src = "crypto_accelerator.v:1854" *) _T_2275;
  assign _T_2407 = _T_2369 & (* src = "crypto_accelerator.v:1855" *) _T_2235;
  assign _T_2409 = _T_2375 & (* src = "crypto_accelerator.v:1856" *) _T_2281;
  assign _T_2411 = _T_2367 & (* src = "crypto_accelerator.v:1857" *) _T_2263;
  assign _T_2556 = _T_2538 & (* src = "crypto_accelerator.v:1925" *) _T_2510;
  assign _T_2558 = _T_2540 & (* src = "crypto_accelerator.v:1926" *) _T_2522;
  assign _T_2562 = _T_2520 & (* src = "crypto_accelerator.v:1928" *) matrix_2_1[0];
  assign _T_2566 = _T_2514 & (* src = "crypto_accelerator.v:1930" *) _T_2542;
  assign _T_2568 = _T_2518 & (* src = "crypto_accelerator.v:1931" *) _T_2508;
  assign _T_2572 = _T_2544 & (* src = "crypto_accelerator.v:1933" *) _T_2534;
  assign _T_2576 = _T_2504 & (* src = "crypto_accelerator.v:1935" *) _T_2516;
  assign _T_2578 = _T_2550 & (* src = "crypto_accelerator.v:1936" *) _T_2546;
  assign _T_2582 = _T_2532 & (* src = "crypto_accelerator.v:1938" *) _T_2528;
  assign _T_2604 = _T_2598 & (* src = "crypto_accelerator.v:1949" *) _T_2594;
  assign _T_2612 = _T_2610 & (* src = "crypto_accelerator.v:1953" *) _T_2608;
  assign _T_2614 = _T_2606 & (* src = "crypto_accelerator.v:1954" *) _T_2602;
  assign _T_2616 = _T_2594 & (* src = "crypto_accelerator.v:1955" *) _T_2600;
  assign _T_2618 = _T_2608 & (* src = "crypto_accelerator.v:1956" *) _T_2616;
  assign _T_2622 = _T_2596 & (* src = "crypto_accelerator.v:1958" *) _T_2598;
  assign _T_2624 = _T_2602 & (* src = "crypto_accelerator.v:1959" *) _T_2622;
  assign _T_2646 = _T_2642 & (* src = "crypto_accelerator.v:1970" *) _T_2510;
  assign _T_2648 = _T_2634 & (* src = "crypto_accelerator.v:1971" *) _T_2522;
  assign _T_2650 = _T_2632 & (* src = "crypto_accelerator.v:1972" *) matrix_2_1[0];
  assign _T_2652 = _T_2640 & (* src = "crypto_accelerator.v:1973" *) _T_2542;
  assign _T_2654 = _T_2630 & (* src = "crypto_accelerator.v:1974" *) _T_2508;
  assign _T_2656 = _T_2628 & (* src = "crypto_accelerator.v:1975" *) _T_2534;
  assign _T_2658 = _T_2638 & (* src = "crypto_accelerator.v:1976" *) _T_2516;
  assign _T_2660 = _T_2644 & (* src = "crypto_accelerator.v:1977" *) _T_2546;
  assign _T_2662 = _T_2636 & (* src = "crypto_accelerator.v:1978" *) _T_2528;
  assign _T_2664 = _T_2642 & (* src = "crypto_accelerator.v:1979" *) _T_2538;
  assign _T_2666 = _T_2634 & (* src = "crypto_accelerator.v:1980" *) _T_2540;
  assign _T_2668 = _T_2632 & (* src = "crypto_accelerator.v:1981" *) _T_2520;
  assign _T_2670 = _T_2640 & (* src = "crypto_accelerator.v:1982" *) _T_2514;
  assign _T_2672 = _T_2630 & (* src = "crypto_accelerator.v:1983" *) _T_2518;
  assign _T_2674 = _T_2628 & (* src = "crypto_accelerator.v:1984" *) _T_2544;
  assign _T_2676 = _T_2638 & (* src = "crypto_accelerator.v:1985" *) _T_2504;
  assign _T_2678 = _T_2644 & (* src = "crypto_accelerator.v:1986" *) _T_2550;
  assign _T_2680 = _T_2636 & (* src = "crypto_accelerator.v:1987" *) _T_2532;
  assign _T_2825 = _T_2807 & (* src = "crypto_accelerator.v:2055" *) _T_2779;
  assign _T_2827 = _T_2809 & (* src = "crypto_accelerator.v:2056" *) _T_2791;
  assign _T_2831 = _T_2789 & (* src = "crypto_accelerator.v:2058" *) matrix_2_2[0];
  assign _T_2835 = _T_2783 & (* src = "crypto_accelerator.v:2060" *) _T_2811;
  assign _T_2837 = _T_2787 & (* src = "crypto_accelerator.v:2061" *) _T_2777;
  assign _T_2841 = _T_2813 & (* src = "crypto_accelerator.v:2063" *) _T_2803;
  assign _T_2845 = _T_2773 & (* src = "crypto_accelerator.v:2065" *) _T_2785;
  assign _T_2847 = _T_2819 & (* src = "crypto_accelerator.v:2066" *) _T_2815;
  assign _T_2851 = _T_2801 & (* src = "crypto_accelerator.v:2068" *) _T_2797;
  assign _T_2873 = _T_2867 & (* src = "crypto_accelerator.v:2079" *) _T_2863;
  assign _T_2881 = _T_2879 & (* src = "crypto_accelerator.v:2083" *) _T_2877;
  assign _T_2883 = _T_2875 & (* src = "crypto_accelerator.v:2084" *) _T_2871;
  assign _T_2885 = _T_2863 & (* src = "crypto_accelerator.v:2085" *) _T_2869;
  assign _T_2887 = _T_2877 & (* src = "crypto_accelerator.v:2086" *) _T_2885;
  assign _T_2891 = _T_2865 & (* src = "crypto_accelerator.v:2088" *) _T_2867;
  assign _T_2893 = _T_2871 & (* src = "crypto_accelerator.v:2089" *) _T_2891;
  assign _T_2915 = _T_2911 & (* src = "crypto_accelerator.v:2100" *) _T_2779;
  assign _T_2917 = _T_2903 & (* src = "crypto_accelerator.v:2101" *) _T_2791;
  assign _T_2919 = _T_2901 & (* src = "crypto_accelerator.v:2102" *) matrix_2_2[0];
  assign _T_2921 = _T_2909 & (* src = "crypto_accelerator.v:2103" *) _T_2811;
  assign _T_2923 = _T_2899 & (* src = "crypto_accelerator.v:2104" *) _T_2777;
  assign _T_2925 = _T_2897 & (* src = "crypto_accelerator.v:2105" *) _T_2803;
  assign _T_2927 = _T_2907 & (* src = "crypto_accelerator.v:2106" *) _T_2785;
  assign _T_2929 = _T_2913 & (* src = "crypto_accelerator.v:2107" *) _T_2815;
  assign _T_2931 = _T_2905 & (* src = "crypto_accelerator.v:2108" *) _T_2797;
  assign _T_2933 = _T_2911 & (* src = "crypto_accelerator.v:2109" *) _T_2807;
  assign _T_2935 = _T_2903 & (* src = "crypto_accelerator.v:2110" *) _T_2809;
  assign _T_2937 = _T_2901 & (* src = "crypto_accelerator.v:2111" *) _T_2789;
  assign _T_2939 = _T_2909 & (* src = "crypto_accelerator.v:2112" *) _T_2783;
  assign _T_2941 = _T_2899 & (* src = "crypto_accelerator.v:2113" *) _T_2787;
  assign _T_2943 = _T_2897 & (* src = "crypto_accelerator.v:2114" *) _T_2813;
  assign _T_2945 = _T_2907 & (* src = "crypto_accelerator.v:2115" *) _T_2773;
  assign _T_2947 = _T_2913 & (* src = "crypto_accelerator.v:2116" *) _T_2819;
  assign _T_2949 = _T_2905 & (* src = "crypto_accelerator.v:2117" *) _T_2801;
  assign _T_3094 = _T_3076 & (* src = "crypto_accelerator.v:2185" *) _T_3048;
  assign _T_3096 = _T_3078 & (* src = "crypto_accelerator.v:2186" *) _T_3060;
  assign _T_3100 = _T_3058 & (* src = "crypto_accelerator.v:2188" *) matrix_2_3[0];
  assign _T_3104 = _T_3052 & (* src = "crypto_accelerator.v:2190" *) _T_3080;
  assign _T_3106 = _T_3056 & (* src = "crypto_accelerator.v:2191" *) _T_3046;
  assign _T_3110 = _T_3082 & (* src = "crypto_accelerator.v:2193" *) _T_3072;
  assign _T_3114 = _T_3042 & (* src = "crypto_accelerator.v:2195" *) _T_3054;
  assign _T_3116 = _T_3088 & (* src = "crypto_accelerator.v:2196" *) _T_3084;
  assign _T_3120 = _T_3070 & (* src = "crypto_accelerator.v:2198" *) _T_3066;
  assign _T_3142 = _T_3136 & (* src = "crypto_accelerator.v:2209" *) _T_3132;
  assign _T_3150 = _T_3148 & (* src = "crypto_accelerator.v:2213" *) _T_3146;
  assign _T_3152 = _T_3144 & (* src = "crypto_accelerator.v:2214" *) _T_3140;
  assign _T_3154 = _T_3132 & (* src = "crypto_accelerator.v:2215" *) _T_3138;
  assign _T_3156 = _T_3146 & (* src = "crypto_accelerator.v:2216" *) _T_3154;
  assign _T_3160 = _T_3134 & (* src = "crypto_accelerator.v:2218" *) _T_3136;
  assign _T_3162 = _T_3140 & (* src = "crypto_accelerator.v:2219" *) _T_3160;
  assign _T_3184 = _T_3180 & (* src = "crypto_accelerator.v:2230" *) _T_3048;
  assign _T_3186 = _T_3172 & (* src = "crypto_accelerator.v:2231" *) _T_3060;
  assign _T_3188 = _T_3170 & (* src = "crypto_accelerator.v:2232" *) matrix_2_3[0];
  assign _T_3190 = _T_3178 & (* src = "crypto_accelerator.v:2233" *) _T_3080;
  assign _T_3192 = _T_3168 & (* src = "crypto_accelerator.v:2234" *) _T_3046;
  assign _T_3194 = _T_3166 & (* src = "crypto_accelerator.v:2235" *) _T_3072;
  assign _T_3196 = _T_3176 & (* src = "crypto_accelerator.v:2236" *) _T_3054;
  assign _T_3198 = _T_3182 & (* src = "crypto_accelerator.v:2237" *) _T_3084;
  assign _T_3200 = _T_3174 & (* src = "crypto_accelerator.v:2238" *) _T_3066;
  assign _T_3202 = _T_3180 & (* src = "crypto_accelerator.v:2239" *) _T_3076;
  assign _T_3204 = _T_3172 & (* src = "crypto_accelerator.v:2240" *) _T_3078;
  assign _T_3206 = _T_3170 & (* src = "crypto_accelerator.v:2241" *) _T_3058;
  assign _T_3208 = _T_3178 & (* src = "crypto_accelerator.v:2242" *) _T_3052;
  assign _T_3210 = _T_3168 & (* src = "crypto_accelerator.v:2243" *) _T_3056;
  assign _T_3212 = _T_3166 & (* src = "crypto_accelerator.v:2244" *) _T_3082;
  assign _T_3214 = _T_3176 & (* src = "crypto_accelerator.v:2245" *) _T_3042;
  assign _T_3216 = _T_3182 & (* src = "crypto_accelerator.v:2246" *) _T_3088;
  assign _T_3218 = _T_3174 & (* src = "crypto_accelerator.v:2247" *) _T_3070;
  assign _T_3364 = _T_3346 & (* src = "crypto_accelerator.v:2315" *) _T_3318;
  assign _T_3366 = _T_3348 & (* src = "crypto_accelerator.v:2316" *) _T_3330;
  assign _T_3370 = _T_3328 & (* src = "crypto_accelerator.v:2318" *) matrix_3_0[0];
  assign _T_3374 = _T_3322 & (* src = "crypto_accelerator.v:2320" *) _T_3350;
  assign _T_3376 = _T_3326 & (* src = "crypto_accelerator.v:2321" *) _T_3316;
  assign _T_3380 = _T_3352 & (* src = "crypto_accelerator.v:2323" *) _T_3342;
  assign _T_3384 = _T_3312 & (* src = "crypto_accelerator.v:2325" *) _T_3324;
  assign _T_3386 = _T_3358 & (* src = "crypto_accelerator.v:2326" *) _T_3354;
  assign _T_3390 = _T_3340 & (* src = "crypto_accelerator.v:2328" *) _T_3336;
  assign _T_3412 = _T_3406 & (* src = "crypto_accelerator.v:2339" *) _T_3402;
  assign _T_3420 = _T_3418 & (* src = "crypto_accelerator.v:2343" *) _T_3416;
  assign _T_3422 = _T_3414 & (* src = "crypto_accelerator.v:2344" *) _T_3410;
  assign _T_3424 = _T_3402 & (* src = "crypto_accelerator.v:2345" *) _T_3408;
  assign _T_3426 = _T_3416 & (* src = "crypto_accelerator.v:2346" *) _T_3424;
  assign _T_3430 = _T_3404 & (* src = "crypto_accelerator.v:2348" *) _T_3406;
  assign _T_3432 = _T_3410 & (* src = "crypto_accelerator.v:2349" *) _T_3430;
  assign _T_3454 = _T_3450 & (* src = "crypto_accelerator.v:2360" *) _T_3318;
  assign _T_3456 = _T_3442 & (* src = "crypto_accelerator.v:2361" *) _T_3330;
  assign _T_3458 = _T_3440 & (* src = "crypto_accelerator.v:2362" *) matrix_3_0[0];
  assign _T_3460 = _T_3448 & (* src = "crypto_accelerator.v:2363" *) _T_3350;
  assign _T_3462 = _T_3438 & (* src = "crypto_accelerator.v:2364" *) _T_3316;
  assign _T_3464 = _T_3436 & (* src = "crypto_accelerator.v:2365" *) _T_3342;
  assign _T_3466 = _T_3446 & (* src = "crypto_accelerator.v:2366" *) _T_3324;
  assign _T_3468 = _T_3452 & (* src = "crypto_accelerator.v:2367" *) _T_3354;
  assign _T_3470 = _T_3444 & (* src = "crypto_accelerator.v:2368" *) _T_3336;
  assign _T_3472 = _T_3450 & (* src = "crypto_accelerator.v:2369" *) _T_3346;
  assign _T_3474 = _T_3442 & (* src = "crypto_accelerator.v:2370" *) _T_3348;
  assign _T_3476 = _T_3440 & (* src = "crypto_accelerator.v:2371" *) _T_3328;
  assign _T_3478 = _T_3448 & (* src = "crypto_accelerator.v:2372" *) _T_3322;
  assign _T_3480 = _T_3438 & (* src = "crypto_accelerator.v:2373" *) _T_3326;
  assign _T_3482 = _T_3436 & (* src = "crypto_accelerator.v:2374" *) _T_3352;
  assign _T_3484 = _T_3446 & (* src = "crypto_accelerator.v:2375" *) _T_3312;
  assign _T_3486 = _T_3452 & (* src = "crypto_accelerator.v:2376" *) _T_3358;
  assign _T_3488 = _T_3444 & (* src = "crypto_accelerator.v:2377" *) _T_3340;
  assign _T_3633 = _T_3615 & (* src = "crypto_accelerator.v:2445" *) _T_3587;
  assign _T_3635 = _T_3617 & (* src = "crypto_accelerator.v:2446" *) _T_3599;
  assign _T_3639 = _T_3597 & (* src = "crypto_accelerator.v:2448" *) matrix_3_1[0];
  assign _T_3643 = _T_3591 & (* src = "crypto_accelerator.v:2450" *) _T_3619;
  assign _T_3645 = _T_3595 & (* src = "crypto_accelerator.v:2451" *) _T_3585;
  assign _T_3649 = _T_3621 & (* src = "crypto_accelerator.v:2453" *) _T_3611;
  assign _T_3653 = _T_3581 & (* src = "crypto_accelerator.v:2455" *) _T_3593;
  assign _T_3655 = _T_3627 & (* src = "crypto_accelerator.v:2456" *) _T_3623;
  assign _T_3659 = _T_3609 & (* src = "crypto_accelerator.v:2458" *) _T_3605;
  assign _T_3681 = _T_3675 & (* src = "crypto_accelerator.v:2469" *) _T_3671;
  assign _T_3689 = _T_3687 & (* src = "crypto_accelerator.v:2473" *) _T_3685;
  assign _T_3691 = _T_3683 & (* src = "crypto_accelerator.v:2474" *) _T_3679;
  assign _T_3693 = _T_3671 & (* src = "crypto_accelerator.v:2475" *) _T_3677;
  assign _T_3695 = _T_3685 & (* src = "crypto_accelerator.v:2476" *) _T_3693;
  assign _T_3699 = _T_3673 & (* src = "crypto_accelerator.v:2478" *) _T_3675;
  assign _T_3701 = _T_3679 & (* src = "crypto_accelerator.v:2479" *) _T_3699;
  assign _T_3723 = _T_3719 & (* src = "crypto_accelerator.v:2490" *) _T_3587;
  assign _T_3725 = _T_3711 & (* src = "crypto_accelerator.v:2491" *) _T_3599;
  assign _T_3727 = _T_3709 & (* src = "crypto_accelerator.v:2492" *) matrix_3_1[0];
  assign _T_3729 = _T_3717 & (* src = "crypto_accelerator.v:2493" *) _T_3619;
  assign _T_3731 = _T_3707 & (* src = "crypto_accelerator.v:2494" *) _T_3585;
  assign _T_3733 = _T_3705 & (* src = "crypto_accelerator.v:2495" *) _T_3611;
  assign _T_3735 = _T_3715 & (* src = "crypto_accelerator.v:2496" *) _T_3593;
  assign _T_3737 = _T_3721 & (* src = "crypto_accelerator.v:2497" *) _T_3623;
  assign _T_3739 = _T_3713 & (* src = "crypto_accelerator.v:2498" *) _T_3605;
  assign _T_3741 = _T_3719 & (* src = "crypto_accelerator.v:2499" *) _T_3615;
  assign _T_3743 = _T_3711 & (* src = "crypto_accelerator.v:2500" *) _T_3617;
  assign _T_3745 = _T_3709 & (* src = "crypto_accelerator.v:2501" *) _T_3597;
  assign _T_3747 = _T_3717 & (* src = "crypto_accelerator.v:2502" *) _T_3591;
  assign _T_3749 = _T_3707 & (* src = "crypto_accelerator.v:2503" *) _T_3595;
  assign _T_3751 = _T_3705 & (* src = "crypto_accelerator.v:2504" *) _T_3621;
  assign _T_3753 = _T_3715 & (* src = "crypto_accelerator.v:2505" *) _T_3581;
  assign _T_3755 = _T_3721 & (* src = "crypto_accelerator.v:2506" *) _T_3627;
  assign _T_3757 = _T_3713 & (* src = "crypto_accelerator.v:2507" *) _T_3609;
  assign _T_3902 = _T_3884 & (* src = "crypto_accelerator.v:2575" *) _T_3856;
  assign _T_3904 = _T_3886 & (* src = "crypto_accelerator.v:2576" *) _T_3868;
  assign _T_3908 = _T_3866 & (* src = "crypto_accelerator.v:2578" *) matrix_3_2[0];
  assign _T_3912 = _T_3860 & (* src = "crypto_accelerator.v:2580" *) _T_3888;
  assign _T_3914 = _T_3864 & (* src = "crypto_accelerator.v:2581" *) _T_3854;
  assign _T_3918 = _T_3890 & (* src = "crypto_accelerator.v:2583" *) _T_3880;
  assign _T_3922 = _T_3850 & (* src = "crypto_accelerator.v:2585" *) _T_3862;
  assign _T_3924 = _T_3896 & (* src = "crypto_accelerator.v:2586" *) _T_3892;
  assign _T_3928 = _T_3878 & (* src = "crypto_accelerator.v:2588" *) _T_3874;
  assign _T_3950 = _T_3944 & (* src = "crypto_accelerator.v:2599" *) _T_3940;
  assign _T_3958 = _T_3956 & (* src = "crypto_accelerator.v:2603" *) _T_3954;
  assign _T_3960 = _T_3952 & (* src = "crypto_accelerator.v:2604" *) _T_3948;
  assign _T_3962 = _T_3940 & (* src = "crypto_accelerator.v:2605" *) _T_3946;
  assign _T_3964 = _T_3954 & (* src = "crypto_accelerator.v:2606" *) _T_3962;
  assign _T_3968 = _T_3942 & (* src = "crypto_accelerator.v:2608" *) _T_3944;
  assign _T_3970 = _T_3948 & (* src = "crypto_accelerator.v:2609" *) _T_3968;
  assign _T_3992 = _T_3988 & (* src = "crypto_accelerator.v:2620" *) _T_3856;
  assign _T_3994 = _T_3980 & (* src = "crypto_accelerator.v:2621" *) _T_3868;
  assign _T_3996 = _T_3978 & (* src = "crypto_accelerator.v:2622" *) matrix_3_2[0];
  assign _T_3998 = _T_3986 & (* src = "crypto_accelerator.v:2623" *) _T_3888;
  assign _T_4000 = _T_3976 & (* src = "crypto_accelerator.v:2624" *) _T_3854;
  assign _T_4002 = _T_3974 & (* src = "crypto_accelerator.v:2625" *) _T_3880;
  assign _T_4004 = _T_3984 & (* src = "crypto_accelerator.v:2626" *) _T_3862;
  assign _T_4006 = _T_3990 & (* src = "crypto_accelerator.v:2627" *) _T_3892;
  assign _T_4008 = _T_3982 & (* src = "crypto_accelerator.v:2628" *) _T_3874;
  assign _T_4010 = _T_3988 & (* src = "crypto_accelerator.v:2629" *) _T_3884;
  assign _T_4012 = _T_3980 & (* src = "crypto_accelerator.v:2630" *) _T_3886;
  assign _T_4014 = _T_3978 & (* src = "crypto_accelerator.v:2631" *) _T_3866;
  assign _T_4016 = _T_3986 & (* src = "crypto_accelerator.v:2632" *) _T_3860;
  assign _T_4018 = _T_3976 & (* src = "crypto_accelerator.v:2633" *) _T_3864;
  assign _T_4020 = _T_3974 & (* src = "crypto_accelerator.v:2634" *) _T_3890;
  assign _T_4022 = _T_3984 & (* src = "crypto_accelerator.v:2635" *) _T_3850;
  assign _T_4024 = _T_3990 & (* src = "crypto_accelerator.v:2636" *) _T_3896;
  assign _T_4026 = _T_3982 & (* src = "crypto_accelerator.v:2637" *) _T_3878;
  assign _T_4171 = _T_4153 & (* src = "crypto_accelerator.v:2705" *) _T_4125;
  assign _T_4173 = _T_4155 & (* src = "crypto_accelerator.v:2706" *) _T_4137;
  assign _T_4177 = _T_4135 & (* src = "crypto_accelerator.v:2708" *) matrix_3_3[0];
  assign _T_4181 = _T_4129 & (* src = "crypto_accelerator.v:2710" *) _T_4157;
  assign _T_4183 = _T_4133 & (* src = "crypto_accelerator.v:2711" *) _T_4123;
  assign _T_4187 = _T_4159 & (* src = "crypto_accelerator.v:2713" *) _T_4149;
  assign _T_4191 = _T_4119 & (* src = "crypto_accelerator.v:2715" *) _T_4131;
  assign _T_4193 = _T_4165 & (* src = "crypto_accelerator.v:2716" *) _T_4161;
  assign _T_4197 = _T_4147 & (* src = "crypto_accelerator.v:2718" *) _T_4143;
  assign _T_4219 = _T_4213 & (* src = "crypto_accelerator.v:2729" *) _T_4209;
  assign _T_4227 = _T_4225 & (* src = "crypto_accelerator.v:2733" *) _T_4223;
  assign _T_4229 = _T_4221 & (* src = "crypto_accelerator.v:2734" *) _T_4217;
  assign _T_4231 = _T_4209 & (* src = "crypto_accelerator.v:2735" *) _T_4215;
  assign _T_4233 = _T_4223 & (* src = "crypto_accelerator.v:2736" *) _T_4231;
  assign _T_4237 = _T_4211 & (* src = "crypto_accelerator.v:2738" *) _T_4213;
  assign _T_4239 = _T_4217 & (* src = "crypto_accelerator.v:2739" *) _T_4237;
  assign _T_4261 = _T_4257 & (* src = "crypto_accelerator.v:2750" *) _T_4125;
  assign _T_4263 = _T_4249 & (* src = "crypto_accelerator.v:2751" *) _T_4137;
  assign _T_4265 = _T_4247 & (* src = "crypto_accelerator.v:2752" *) matrix_3_3[0];
  assign _T_4267 = _T_4255 & (* src = "crypto_accelerator.v:2753" *) _T_4157;
  assign _T_4269 = _T_4245 & (* src = "crypto_accelerator.v:2754" *) _T_4123;
  assign _T_4271 = _T_4243 & (* src = "crypto_accelerator.v:2755" *) _T_4149;
  assign _T_4273 = _T_4253 & (* src = "crypto_accelerator.v:2756" *) _T_4131;
  assign _T_4275 = _T_4259 & (* src = "crypto_accelerator.v:2757" *) _T_4161;
  assign _T_4277 = _T_4251 & (* src = "crypto_accelerator.v:2758" *) _T_4143;
  assign _T_4279 = _T_4257 & (* src = "crypto_accelerator.v:2759" *) _T_4153;
  assign _T_4281 = _T_4249 & (* src = "crypto_accelerator.v:2760" *) _T_4155;
  assign _T_4283 = _T_4247 & (* src = "crypto_accelerator.v:2761" *) _T_4135;
  assign _T_4285 = _T_4255 & (* src = "crypto_accelerator.v:2762" *) _T_4129;
  assign _T_4287 = _T_4245 & (* src = "crypto_accelerator.v:2763" *) _T_4133;
  assign _T_4289 = _T_4243 & (* src = "crypto_accelerator.v:2764" *) _T_4159;
  assign _T_4291 = _T_4253 & (* src = "crypto_accelerator.v:2765" *) _T_4119;
  assign _T_4293 = _T_4259 & (* src = "crypto_accelerator.v:2766" *) _T_4165;
  assign _T_4295 = _T_4251 & (* src = "crypto_accelerator.v:2767" *) _T_4147;
  assign _T_4415 = io_ready & (* src = "crypto_accelerator.v:2840" *) io_dataValid;
  assign _T_133 = _T_115 & (* src = "crypto_accelerator.v:755" *) _T_87;
  assign _T_135 = _T_117 & (* src = "crypto_accelerator.v:756" *) _T_99;
  assign _T_139 = _T_97 & (* src = "crypto_accelerator.v:758" *) matrix_0_0[0];
  assign _T_143 = _T_91 & (* src = "crypto_accelerator.v:760" *) _T_119;
  assign _T_145 = _T_95 & (* src = "crypto_accelerator.v:761" *) _T_85;
  assign _T_149 = _T_121 & (* src = "crypto_accelerator.v:763" *) _T_111;
  assign _T_153 = _T_81 & (* src = "crypto_accelerator.v:765" *) _T_93;
  assign _T_155 = _T_127 & (* src = "crypto_accelerator.v:766" *) _T_123;
  assign _T_159 = _T_109 & (* src = "crypto_accelerator.v:768" *) _T_105;
  assign _T_181 = _T_175 & (* src = "crypto_accelerator.v:779" *) _T_171;
  assign _T_189 = _T_187 & (* src = "crypto_accelerator.v:783" *) _T_185;
  assign _T_191 = _T_183 & (* src = "crypto_accelerator.v:784" *) _T_179;
  assign _T_193 = _T_171 & (* src = "crypto_accelerator.v:785" *) _T_177;
  assign _T_195 = _T_185 & (* src = "crypto_accelerator.v:786" *) _T_193;
  assign _T_199 = _T_173 & (* src = "crypto_accelerator.v:788" *) _T_175;
  assign _T_201 = _T_179 & (* src = "crypto_accelerator.v:789" *) _T_199;
  assign _T_223 = _T_219 & (* src = "crypto_accelerator.v:800" *) _T_87;
  assign _T_225 = _T_211 & (* src = "crypto_accelerator.v:801" *) _T_99;
  assign _T_227 = _T_209 & (* src = "crypto_accelerator.v:802" *) matrix_0_0[0];
  assign _T_229 = _T_217 & (* src = "crypto_accelerator.v:803" *) _T_119;
  assign _T_231 = _T_207 & (* src = "crypto_accelerator.v:804" *) _T_85;
  assign _T_233 = _T_205 & (* src = "crypto_accelerator.v:805" *) _T_111;
  assign _T_235 = _T_215 & (* src = "crypto_accelerator.v:806" *) _T_93;
  assign _T_237 = _T_221 & (* src = "crypto_accelerator.v:807" *) _T_123;
  assign _T_239 = _T_213 & (* src = "crypto_accelerator.v:808" *) _T_105;
  assign _T_241 = _T_219 & (* src = "crypto_accelerator.v:809" *) _T_115;
  assign _T_243 = _T_211 & (* src = "crypto_accelerator.v:810" *) _T_117;
  assign _T_245 = _T_209 & (* src = "crypto_accelerator.v:811" *) _T_97;
  assign _T_247 = _T_217 & (* src = "crypto_accelerator.v:812" *) _T_91;
  assign _T_249 = _T_207 & (* src = "crypto_accelerator.v:813" *) _T_95;
  assign _T_251 = _T_205 & (* src = "crypto_accelerator.v:814" *) _T_121;
  assign _T_253 = _T_215 & (* src = "crypto_accelerator.v:815" *) _T_81;
  assign _T_255 = _T_221 & (* src = "crypto_accelerator.v:816" *) _T_127;
  assign _T_257 = _T_213 & (* src = "crypto_accelerator.v:817" *) _T_109;
  assign _T_402 = _T_384 & (* src = "crypto_accelerator.v:885" *) _T_356;
  assign _T_404 = _T_386 & (* src = "crypto_accelerator.v:886" *) _T_368;
  assign _T_408 = _T_366 & (* src = "crypto_accelerator.v:888" *) matrix_0_1[0];
  assign _T_412 = _T_360 & (* src = "crypto_accelerator.v:890" *) _T_388;
  assign _T_414 = _T_364 & (* src = "crypto_accelerator.v:891" *) _T_354;
  assign _T_418 = _T_390 & (* src = "crypto_accelerator.v:893" *) _T_380;
  assign _T_422 = _T_350 & (* src = "crypto_accelerator.v:895" *) _T_362;
  assign _T_424 = _T_396 & (* src = "crypto_accelerator.v:896" *) _T_392;
  assign _T_428 = _T_378 & (* src = "crypto_accelerator.v:898" *) _T_374;
  assign _T_450 = _T_444 & (* src = "crypto_accelerator.v:909" *) _T_440;
  assign _T_458 = _T_456 & (* src = "crypto_accelerator.v:913" *) _T_454;
  assign _T_460 = _T_452 & (* src = "crypto_accelerator.v:914" *) _T_448;
  assign _T_462 = _T_440 & (* src = "crypto_accelerator.v:915" *) _T_446;
  assign _T_464 = _T_454 & (* src = "crypto_accelerator.v:916" *) _T_462;
  assign _T_468 = _T_442 & (* src = "crypto_accelerator.v:918" *) _T_444;
  assign _T_470 = _T_448 & (* src = "crypto_accelerator.v:919" *) _T_468;
  assign _T_492 = _T_488 & (* src = "crypto_accelerator.v:930" *) _T_356;
  assign _T_494 = _T_480 & (* src = "crypto_accelerator.v:931" *) _T_368;
  assign _T_496 = _T_478 & (* src = "crypto_accelerator.v:932" *) matrix_0_1[0];
  assign _T_498 = _T_486 & (* src = "crypto_accelerator.v:933" *) _T_388;
  assign _T_500 = _T_476 & (* src = "crypto_accelerator.v:934" *) _T_354;
  assign _T_502 = _T_474 & (* src = "crypto_accelerator.v:935" *) _T_380;
  assign _T_504 = _T_484 & (* src = "crypto_accelerator.v:936" *) _T_362;
  assign _T_506 = _T_490 & (* src = "crypto_accelerator.v:937" *) _T_392;
  assign _T_508 = _T_482 & (* src = "crypto_accelerator.v:938" *) _T_374;
  assign _T_510 = _T_488 & (* src = "crypto_accelerator.v:939" *) _T_384;
  assign _T_512 = _T_480 & (* src = "crypto_accelerator.v:940" *) _T_386;
  assign _T_514 = _T_478 & (* src = "crypto_accelerator.v:941" *) _T_366;
  assign _T_516 = _T_486 & (* src = "crypto_accelerator.v:942" *) _T_360;
  assign _T_518 = _T_476 & (* src = "crypto_accelerator.v:943" *) _T_364;
  assign _T_520 = _T_474 & (* src = "crypto_accelerator.v:944" *) _T_390;
  assign _T_522 = _T_484 & (* src = "crypto_accelerator.v:945" *) _T_350;
  assign _T_524 = _T_490 & (* src = "crypto_accelerator.v:946" *) _T_396;
  assign _T_526 = _T_482 & (* src = "crypto_accelerator.v:947" *) _T_378;
  assign _T_4420 = state == (* src = "crypto_accelerator.v:2841" *) 5'b11101;
  assign _T_4421 = state == (* src = "crypto_accelerator.v:2842" *) 5'b10101;
  assign io_outputValid = state == (* src = "crypto_accelerator.v:2886" *) 5'b11110;
  assign _T = ! (* src = "crypto_accelerator.v:685" *) state;
  assign _T_1 = state == (* src = "crypto_accelerator.v:686" *) 1'b1;
  assign _T_836 = ~ (* src = "crypto_accelerator.v:1099" *) _T_835;
  assign _T_846 = ~ (* src = "crypto_accelerator.v:1106" *) _T_845;
  assign _T_854 = ~ (* src = "crypto_accelerator.v:1111" *) _T_853;
  assign _T_861 = ~ (* src = "crypto_accelerator.v:1116" *) _T_860;
  assign _T_1105 = ~ (* src = "crypto_accelerator.v:1229" *) _T_1104;
  assign _T_1115 = ~ (* src = "crypto_accelerator.v:1236" *) _T_1114;
  assign _T_1123 = ~ (* src = "crypto_accelerator.v:1241" *) _T_1122;
  assign _T_1130 = ~ (* src = "crypto_accelerator.v:1246" *) _T_1129;
  assign _T_1375 = ~ (* src = "crypto_accelerator.v:1359" *) _T_1374;
  assign _T_1385 = ~ (* src = "crypto_accelerator.v:1366" *) _T_1384;
  assign _T_1393 = ~ (* src = "crypto_accelerator.v:1371" *) _T_1392;
  assign _T_1400 = ~ (* src = "crypto_accelerator.v:1376" *) _T_1399;
  assign _T_1644 = ~ (* src = "crypto_accelerator.v:1489" *) _T_1643;
  assign _T_1654 = ~ (* src = "crypto_accelerator.v:1496" *) _T_1653;
  assign _T_1662 = ~ (* src = "crypto_accelerator.v:1501" *) _T_1661;
  assign _T_1669 = ~ (* src = "crypto_accelerator.v:1506" *) _T_1668;
  assign _T_1913 = ~ (* src = "crypto_accelerator.v:1619" *) _T_1912;
  assign _T_1923 = ~ (* src = "crypto_accelerator.v:1626" *) _T_1922;
  assign _T_1931 = ~ (* src = "crypto_accelerator.v:1631" *) _T_1930;
  assign _T_1938 = ~ (* src = "crypto_accelerator.v:1636" *) _T_1937;
  assign _T_2182 = ~ (* src = "crypto_accelerator.v:1749" *) _T_2181;
  assign _T_2192 = ~ (* src = "crypto_accelerator.v:1756" *) _T_2191;
  assign _T_2200 = ~ (* src = "crypto_accelerator.v:1761" *) _T_2199;
  assign _T_2207 = ~ (* src = "crypto_accelerator.v:1766" *) _T_2206;
  assign _T_2452 = ~ (* src = "crypto_accelerator.v:1879" *) _T_2451;
  assign _T_2462 = ~ (* src = "crypto_accelerator.v:1886" *) _T_2461;
  assign _T_2470 = ~ (* src = "crypto_accelerator.v:1891" *) _T_2469;
  assign _T_2477 = ~ (* src = "crypto_accelerator.v:1896" *) _T_2476;
  assign _T_2721 = ~ (* src = "crypto_accelerator.v:2009" *) _T_2720;
  assign _T_2731 = ~ (* src = "crypto_accelerator.v:2016" *) _T_2730;
  assign _T_2739 = ~ (* src = "crypto_accelerator.v:2021" *) _T_2738;
  assign _T_2746 = ~ (* src = "crypto_accelerator.v:2026" *) _T_2745;
  assign _T_2990 = ~ (* src = "crypto_accelerator.v:2139" *) _T_2989;
  assign _T_3000 = ~ (* src = "crypto_accelerator.v:2146" *) _T_2999;
  assign _T_3008 = ~ (* src = "crypto_accelerator.v:2151" *) _T_3007;
  assign _T_3015 = ~ (* src = "crypto_accelerator.v:2156" *) _T_3014;
  assign _T_3259 = ~ (* src = "crypto_accelerator.v:2269" *) _T_3258;
  assign _T_3269 = ~ (* src = "crypto_accelerator.v:2276" *) _T_3268;
  assign _T_3277 = ~ (* src = "crypto_accelerator.v:2281" *) _T_3276;
  assign _T_3284 = ~ (* src = "crypto_accelerator.v:2286" *) _T_3283;
  assign _T_3529 = ~ (* src = "crypto_accelerator.v:2399" *) _T_3528;
  assign _T_3539 = ~ (* src = "crypto_accelerator.v:2406" *) _T_3538;
  assign _T_3547 = ~ (* src = "crypto_accelerator.v:2411" *) _T_3546;
  assign _T_3554 = ~ (* src = "crypto_accelerator.v:2416" *) _T_3553;
  assign _T_3798 = ~ (* src = "crypto_accelerator.v:2529" *) _T_3797;
  assign _T_3808 = ~ (* src = "crypto_accelerator.v:2536" *) _T_3807;
  assign _T_3816 = ~ (* src = "crypto_accelerator.v:2541" *) _T_3815;
  assign _T_3823 = ~ (* src = "crypto_accelerator.v:2546" *) _T_3822;
  assign _T_4067 = ~ (* src = "crypto_accelerator.v:2659" *) _T_4066;
  assign _T_4077 = ~ (* src = "crypto_accelerator.v:2666" *) _T_4076;
  assign _T_4085 = ~ (* src = "crypto_accelerator.v:2671" *) _T_4084;
  assign _T_4092 = ~ (* src = "crypto_accelerator.v:2676" *) _T_4091;
  assign _T_4336 = ~ (* src = "crypto_accelerator.v:2789" *) _T_4335;
  assign _T_4346 = ~ (* src = "crypto_accelerator.v:2796" *) _T_4345;
  assign _T_4354 = ~ (* src = "crypto_accelerator.v:2801" *) _T_4353;
  assign _T_4361 = ~ (* src = "crypto_accelerator.v:2806" *) _T_4360;
  assign _T_6 = ~ (* src = "crypto_accelerator.v:689" *) io_ready;
  assign _T_298 = ~ (* src = "crypto_accelerator.v:839" *) _T_297;
  assign _T_308 = ~ (* src = "crypto_accelerator.v:846" *) _T_307;
  assign _T_316 = ~ (* src = "crypto_accelerator.v:851" *) _T_315;
  assign _T_323 = ~ (* src = "crypto_accelerator.v:856" *) _T_322;
  assign _T_567 = ~ (* src = "crypto_accelerator.v:969" *) _T_566;
  assign _T_577 = ~ (* src = "crypto_accelerator.v:976" *) _T_576;
  assign _T_585 = ~ (* src = "crypto_accelerator.v:981" *) _T_584;
  assign _T_592 = ~ (* src = "crypto_accelerator.v:986" *) _T_591;
  assign io_shiftCyc = _T_6 | (* src = "crypto_accelerator.v:2881" *) io_dataValid;
  assign io_ready = _T_2 | (* src = "crypto_accelerator.v:2883" *) io_outputValid;
  assign _T_2 = _T | (* src = "crypto_accelerator.v:687" *) _T_1;
  always @(posedge clock)
      state <= _0016_;
  always @(posedge clock)
      matrix_0_0 <= _0000_;
  always @(posedge clock)
      matrix_0_1 <= _0001_;
  always @(posedge clock)
      matrix_0_2 <= _0002_;
  always @(posedge clock)
      matrix_0_3 <= _0003_;
  always @(posedge clock)
      matrix_1_0 <= _0004_;
  always @(posedge clock)
      matrix_1_1 <= _0005_;
  always @(posedge clock)
      matrix_1_2 <= _0006_;
  always @(posedge clock)
      matrix_1_3 <= _0007_;
  always @(posedge clock)
      matrix_2_0 <= _0008_;
  always @(posedge clock)
      matrix_2_1 <= _0009_;
  always @(posedge clock)
      matrix_2_2 <= _0010_;
  always @(posedge clock)
      matrix_2_3 <= _0011_;
  always @(posedge clock)
      matrix_3_0 <= _0012_;
  always @(posedge clock)
      matrix_3_1 <= _0013_;
  always @(posedge clock)
      matrix_3_2 <= _0014_;
  always @(posedge clock)
      matrix_3_3 <= _0015_;
  assign _0017_ = _T_4415 ? (* src = "crypto_accelerator.v:3164" *) _T_41[7:0] : matrix_3_3;
  assign _0018_ = _T_4422 ? (* src = "crypto_accelerator.v:3159" *) roundPart2_last_3_3 : roundPart2_3_3;
  assign _0019_ = state[0] ? (* src = "crypto_accelerator.v:3157" *) _0018_ : { _T_3257, _T_3284, _T_3259, _T_3262, _T_3263, _T_3280, _T_3277, _T_3269 };
  assign _0015_ = io_ready ? (* src = "crypto_accelerator.v:3156" *) _0017_ : _0019_;
  assign _0020_ = _T_4415 ? (* src = "crypto_accelerator.v:3153" *) _T_41[15:8] : matrix_3_2;
  assign _0021_ = _T_4422 ? (* src = "crypto_accelerator.v:3148" *) roundPart2_last_3_2 : roundPart2_3_2;
  assign _0022_ = state[0] ? (* src = "crypto_accelerator.v:3146" *) _0021_ : { _T_1911, _T_1938, _T_1913, _T_1916, _T_1917, _T_1934, _T_1931, _T_1923 };
  assign _0014_ = io_ready ? (* src = "crypto_accelerator.v:3145" *) _0020_ : _0022_;
  assign _0023_ = _T_4415 ? (* src = "crypto_accelerator.v:3142" *) _T_41[23:16] : matrix_3_1;
  assign _0024_ = _T_4422 ? (* src = "crypto_accelerator.v:3137" *) roundPart2_last_3_1 : roundPart2_3_1;
  assign _0025_ = state[0] ? (* src = "crypto_accelerator.v:3135" *) _0024_ : { _T_565, _T_592, _T_567, _T_570, _T_571, _T_588, _T_585, _T_577 };
  assign _0013_ = io_ready ? (* src = "crypto_accelerator.v:3134" *) _0023_ : _0025_;
  assign _0026_ = _T_4415 ? (* src = "crypto_accelerator.v:3131" *) _T_41[31:24] : matrix_3_0;
  assign _0027_ = _T_4422 ? (* src = "crypto_accelerator.v:3126" *) roundPart2_last_3_0 : roundPart2_3_0;
  assign _0028_ = state[0] ? (* src = "crypto_accelerator.v:3124" *) _0027_ : { _T_3527, _T_3554, _T_3529, _T_3532, _T_3533, _T_3550, _T_3547, _T_3539 };
  assign _0012_ = io_ready ? (* src = "crypto_accelerator.v:3123" *) _0026_ : _0028_;
  assign _0029_ = _T_4415 ? (* src = "crypto_accelerator.v:3120" *) _T_41[39:32] : matrix_2_3;
  assign _0030_ = _T_4422 ? (* src = "crypto_accelerator.v:3115" *) roundPart2_last_2_3 : roundPart2_2_3;
  assign _0031_ = state[0] ? (* src = "crypto_accelerator.v:3113" *) _0030_ : { _T_2180, _T_2207, _T_2182, _T_2185, _T_2186, _T_2203, _T_2200, _T_2192 };
  assign _0011_ = io_ready ? (* src = "crypto_accelerator.v:3112" *) _0029_ : _0031_;
  assign _0032_ = _T_4415 ? (* src = "crypto_accelerator.v:3109" *) _T_41[47:40] : matrix_2_2;
  assign _0033_ = _T_4422 ? (* src = "crypto_accelerator.v:3104" *) roundPart2_last_2_2 : roundPart2_2_2;
  assign _0034_ = state[0] ? (* src = "crypto_accelerator.v:3102" *) _0033_ : { _T_834, _T_861, _T_836, _T_839, _T_840, _T_857, _T_854, _T_846 };
  assign _0010_ = io_ready ? (* src = "crypto_accelerator.v:3101" *) _0032_ : _0034_;
  assign _0035_ = _T_4415 ? (* src = "crypto_accelerator.v:3098" *) _T_41[55:48] : matrix_2_1;
  assign _0036_ = _T_4422 ? (* src = "crypto_accelerator.v:3093" *) roundPart2_last_2_1 : roundPart2_2_1;
  assign _0037_ = state[0] ? (* src = "crypto_accelerator.v:3091" *) _0036_ : { _T_3796, _T_3823, _T_3798, _T_3801, _T_3802, _T_3819, _T_3816, _T_3808 };
  assign _0009_ = io_ready ? (* src = "crypto_accelerator.v:3090" *) _0035_ : _0037_;
  assign _0038_ = _T_4415 ? (* src = "crypto_accelerator.v:3087" *) _T_41[63:56] : matrix_2_0;
  assign _0039_ = _T_4422 ? (* src = "crypto_accelerator.v:3082" *) roundPart2_last_2_0 : roundPart2_2_0;
  assign _0040_ = state[0] ? (* src = "crypto_accelerator.v:3080" *) _0039_ : { _T_2450, _T_2477, _T_2452, _T_2455, _T_2456, _T_2473, _T_2470, _T_2462 };
  assign _0008_ = io_ready ? (* src = "crypto_accelerator.v:3079" *) _0038_ : _0040_;
  assign _0041_ = _T_4415 ? (* src = "crypto_accelerator.v:3076" *) _T_41[71:64] : matrix_1_3;
  assign _0042_ = _T_4422 ? (* src = "crypto_accelerator.v:3071" *) roundPart2_last_1_3 : roundPart2_1_3;
  assign _0043_ = state[0] ? (* src = "crypto_accelerator.v:3069" *) _0042_ : { _T_1103, _T_1130, _T_1105, _T_1108, _T_1109, _T_1126, _T_1123, _T_1115 };
  assign _0007_ = io_ready ? (* src = "crypto_accelerator.v:3068" *) _0041_ : _0043_;
  assign _0044_ = _T_4415 ? (* src = "crypto_accelerator.v:3065" *) _T_41[79:72] : matrix_1_2;
  assign _0045_ = _T_4422 ? (* src = "crypto_accelerator.v:3060" *) roundPart2_last_1_2 : roundPart2_1_2;
  assign _0046_ = state[0] ? (* src = "crypto_accelerator.v:3058" *) _0045_ : { _T_4065, _T_4092, _T_4067, _T_4070, _T_4071, _T_4088, _T_4085, _T_4077 };
  assign _0006_ = io_ready ? (* src = "crypto_accelerator.v:3057" *) _0044_ : _0046_;
  assign _0047_ = _T_4415 ? (* src = "crypto_accelerator.v:3054" *) _T_41[87:80] : matrix_1_1;
  assign _0048_ = _T_4422 ? (* src = "crypto_accelerator.v:3049" *) roundPart2_last_1_1 : roundPart2_1_1;
  assign _0049_ = state[0] ? (* src = "crypto_accelerator.v:3047" *) _0048_ : { _T_2719, _T_2746, _T_2721, _T_2724, _T_2725, _T_2742, _T_2739, _T_2731 };
  assign _0005_ = io_ready ? (* src = "crypto_accelerator.v:3046" *) _0047_ : _0049_;
  assign _0050_ = _T_4415 ? (* src = "crypto_accelerator.v:3043" *) _T_41[95:88] : matrix_1_0;
  assign _0051_ = _T_4422 ? (* src = "crypto_accelerator.v:3038" *) roundPart2_last_1_0 : roundPart2_1_0;
  assign _0052_ = state[0] ? (* src = "crypto_accelerator.v:3036" *) _0051_ : { _T_1373, _T_1400, _T_1375, _T_1378, _T_1379, _T_1396, _T_1393, _T_1385 };
  assign _0004_ = io_ready ? (* src = "crypto_accelerator.v:3035" *) _0050_ : _0052_;
  assign _0053_ = _T_4415 ? (* src = "crypto_accelerator.v:3032" *) _T_41[103:96] : matrix_0_3;
  assign _0054_ = _T_4422 ? (* src = "crypto_accelerator.v:3027" *) roundPart2_last_0_3 : roundPart2_0_3;
  assign _0055_ = state[0] ? (* src = "crypto_accelerator.v:3025" *) _0054_ : { _T_4334, _T_4361, _T_4336, _T_4339, _T_4340, _T_4357, _T_4354, _T_4346 };
  assign _0003_ = io_ready ? (* src = "crypto_accelerator.v:3024" *) _0053_ : _0055_;
  assign _0056_ = _T_4415 ? (* src = "crypto_accelerator.v:3021" *) _T_41[111:104] : matrix_0_2;
  assign _0057_ = _T_4422 ? (* src = "crypto_accelerator.v:3016" *) roundPart2_last_0_2 : roundPart2_0_2;
  assign _0058_ = state[0] ? (* src = "crypto_accelerator.v:3014" *) _0057_ : { _T_2988, _T_3015, _T_2990, _T_2993, _T_2994, _T_3011, _T_3008, _T_3000 };
  assign _0002_ = io_ready ? (* src = "crypto_accelerator.v:3013" *) _0056_ : _0058_;
  assign _0059_ = _T_4415 ? (* src = "crypto_accelerator.v:3010" *) _T_41[119:112] : matrix_0_1;
  assign _0060_ = _T_4422 ? (* src = "crypto_accelerator.v:3005" *) roundPart2_last_0_1 : roundPart2_0_1;
  assign _0061_ = state[0] ? (* src = "crypto_accelerator.v:3003" *) _0060_ : { _T_1642, _T_1669, _T_1644, _T_1647, _T_1648, _T_1665, _T_1662, _T_1654 };
  assign _0001_ = io_ready ? (* src = "crypto_accelerator.v:3002" *) _0059_ : _0061_;
  assign _0062_ = _T_4415 ? (* src = "crypto_accelerator.v:2999" *) _T_41[127:120] : matrix_0_0;
  assign _0063_ = _T_4422 ? (* src = "crypto_accelerator.v:2994" *) roundPart2_last_0_0 : roundPart2_0_0;
  assign _0064_ = state[0] ? (* src = "crypto_accelerator.v:2992" *) _0063_ : { _T_296, _T_323, _T_298, _T_301, _T_302, _T_319, _T_316, _T_308 };
  assign _0000_ = io_ready ? (* src = "crypto_accelerator.v:2991" *) _0062_ : _0064_;
  assign _0065_ = _T_4415 ? (* src = "crypto_accelerator.v:2988" *) 6'b000010 : state;
  assign _0066_ = _T_4422 ? (* src = "crypto_accelerator.v:2983" *) 6'b011110 : _T_4427;
  assign _0067_ = io_ready ? (* src = "crypto_accelerator.v:2982" *) _0065_ : _0066_;
  assign _0016_ = reset ? (* src = "crypto_accelerator.v:2980" *) 6'b000001 : _0067_;
  assign _T_4422 = io_aes256 ? (* src = "crypto_accelerator.v:2843" *) _T_4420 : _T_4421;
  assign _GEN_34 = state[0] ? (* src = "crypto_accelerator.v:2845" *) 1'b1 : _T_4415;
  assign io_shift = io_ready ? (* src = "crypto_accelerator.v:2882" *) _T_4415 : _GEN_34;
  assign _T_641 = matrix_0_2[5] ^ (* src = "crypto_accelerator.v:1000" *) matrix_0_2[2];
  assign _T_643 = _T_621 ^ (* src = "crypto_accelerator.v:1001" *) _T_625;
  assign _T_645 = matrix_0_2[2] ^ (* src = "crypto_accelerator.v:1002" *) _T_629;
  assign _T_647 = matrix_0_2[7] ^ (* src = "crypto_accelerator.v:1003" *) matrix_0_2[2];
  assign _T_649 = matrix_0_2[0] ^ (* src = "crypto_accelerator.v:1004" *) _T_631;
  assign _T_651 = matrix_0_2[1] ^ (* src = "crypto_accelerator.v:1005" *) matrix_0_2[2];
  assign _T_653 = _T_619 ^ (* src = "crypto_accelerator.v:1006" *) _T_651;
  assign _T_655 = _T_623 ^ (* src = "crypto_accelerator.v:1007" *) _T_645;
  assign _T_657 = _T_617 ^ (* src = "crypto_accelerator.v:1008" *) _T_641;
  assign _T_659 = matrix_0_2[7] ^ (* src = "crypto_accelerator.v:1009" *) _T_623;
  assign _T_661 = _T_657 ^ (* src = "crypto_accelerator.v:1010" *) _T_625;
  assign _T_663 = _T_657 ^ (* src = "crypto_accelerator.v:1011" *) _T_629;
  assign _T_665 = _T_629 ^ (* src = "crypto_accelerator.v:1012" *) _T_653;
  assign _T_667 = _T_647 ^ (* src = "crypto_accelerator.v:1013" *) _T_643;
  assign _T_669 = _T_659 ^ (* src = "crypto_accelerator.v:1014" *) _T_649;
  assign _T_675 = _T_639 ^ (* src = "crypto_accelerator.v:1017" *) _T_671;
  assign _T_679 = _T_677 ^ (* src = "crypto_accelerator.v:1019" *) _T_671;
  assign _T_685 = _T_663 ^ (* src = "crypto_accelerator.v:1022" *) _T_681;
  assign _T_689 = _T_687 ^ (* src = "crypto_accelerator.v:1024" *) _T_681;
  assign _T_695 = _T_693 ^ (* src = "crypto_accelerator.v:1027" *) _T_691;
  assign _T_699 = _T_697 ^ (* src = "crypto_accelerator.v:1029" *) _T_691;
  assign _T_701 = _T_675 ^ (* src = "crypto_accelerator.v:1030" *) _T_673;
  assign _T_703 = _T_679 ^ (* src = "crypto_accelerator.v:1031" *) _T_667;
  assign _T_705 = _T_685 ^ (* src = "crypto_accelerator.v:1032" *) _T_683;
  assign _T_707 = _T_689 ^ (* src = "crypto_accelerator.v:1033" *) _T_699;
  assign _T_709 = _T_701 ^ (* src = "crypto_accelerator.v:1034" *) _T_695;
  assign _T_711 = _T_703 ^ (* src = "crypto_accelerator.v:1035" *) _T_699;
  assign _T_713 = _T_705 ^ (* src = "crypto_accelerator.v:1036" *) _T_695;
  assign _T_715 = _T_707 ^ (* src = "crypto_accelerator.v:1037" *) _T_669;
  assign _T_717 = _T_713 ^ (* src = "crypto_accelerator.v:1038" *) _T_715;
  assign _T_721 = _T_711 ^ (* src = "crypto_accelerator.v:1040" *) _T_719;
  assign _T_723 = _T_709 ^ (* src = "crypto_accelerator.v:1041" *) _T_711;
  assign _T_725 = _T_715 ^ (* src = "crypto_accelerator.v:1042" *) _T_719;
  assign _T_735 = _T_723 ^ (* src = "crypto_accelerator.v:1047" *) _T_719;
  assign _T_741 = _T_717 ^ (* src = "crypto_accelerator.v:1050" *) _T_719;
  assign _T_743 = _T_711 ^ (* src = "crypto_accelerator.v:1051" *) _T_727;
  assign _T_745 = _T_733 ^ (* src = "crypto_accelerator.v:1052" *) _T_735;
  assign _T_747 = _T_715 ^ (* src = "crypto_accelerator.v:1053" *) _T_729;
  assign _T_749 = _T_739 ^ (* src = "crypto_accelerator.v:1054" *) _T_741;
  assign _T_751 = _T_745 ^ (* src = "crypto_accelerator.v:1055" *) _T_749;
  assign _T_753 = _T_743 ^ (* src = "crypto_accelerator.v:1056" *) _T_747;
  assign _T_755 = _T_743 ^ (* src = "crypto_accelerator.v:1057" *) _T_745;
  assign _T_757 = _T_747 ^ (* src = "crypto_accelerator.v:1058" *) _T_749;
  assign _T_759 = _T_753 ^ (* src = "crypto_accelerator.v:1059" *) _T_751;
  assign _T_797 = _T_791 ^ (* src = "crypto_accelerator.v:1078" *) _T_793;
  assign _T_799 = _T_769 ^ (* src = "crypto_accelerator.v:1079" *) _T_781;
  assign _T_801 = _T_775 ^ (* src = "crypto_accelerator.v:1080" *) _T_797;
  assign _T_803 = _T_779 ^ (* src = "crypto_accelerator.v:1081" *) _T_799;
  assign _T_805 = _T_765 ^ (* src = "crypto_accelerator.v:1082" *) _T_785;
  assign _T_807 = _T_761 ^ (* src = "crypto_accelerator.v:1083" *) _T_767;
  assign _T_809 = _T_797 ^ (* src = "crypto_accelerator.v:1084" *) _T_807;
  assign _T_811 = _T_763 ^ (* src = "crypto_accelerator.v:1085" *) _T_803;
  assign _T_813 = _T_761 ^ (* src = "crypto_accelerator.v:1086" *) _T_773;
  assign _T_815 = _T_771 ^ (* src = "crypto_accelerator.v:1087" *) _T_787;
  assign _T_817 = _T_777 ^ (* src = "crypto_accelerator.v:1088" *) _T_789;
  assign _T_819 = _T_765 ^ (* src = "crypto_accelerator.v:1089" *) _T_811;
  assign _T_821 = _T_805 ^ (* src = "crypto_accelerator.v:1090" *) _T_817;
  assign _T_823 = _T_783 ^ (* src = "crypto_accelerator.v:1091" *) _T_799;
  assign _T_825 = _T_767 ^ (* src = "crypto_accelerator.v:1092" *) _T_773;
  assign _T_827 = _T_803 ^ (* src = "crypto_accelerator.v:1093" *) _T_825;
  assign _T_829 = _T_795 ^ (* src = "crypto_accelerator.v:1094" *) _T_821;
  assign _T_831 = _T_791 ^ (* src = "crypto_accelerator.v:1095" *) _T_813;
  assign _T_833 = _T_805 ^ (* src = "crypto_accelerator.v:1096" *) _T_815;
  assign _T_834 = _T_801 ^ (* src = "crypto_accelerator.v:1097" *) _T_827;
  assign _T_835 = _T_829 ^ (* src = "crypto_accelerator.v:1098" *) _T_831;
  assign _T_838 = _T_771 ^ (* src = "crypto_accelerator.v:1100" *) _T_797;
  assign _T_839 = _T_809 ^ (* src = "crypto_accelerator.v:1101" *) _T_811;
  assign _T_840 = _T_819 ^ (* src = "crypto_accelerator.v:1102" *) _T_838;
  assign _T_842 = _T_769 ^ (* src = "crypto_accelerator.v:1103" *) _T_785;
  assign _T_844 = _T_807 ^ (* src = "crypto_accelerator.v:1104" *) _T_823;
  assign _T_845 = _T_809 ^ (* src = "crypto_accelerator.v:1105" *) _T_833;
  assign _T_848 = _T_777 ^ (* src = "crypto_accelerator.v:1107" *) _T_815;
  assign _T_850 = _T_842 ^ (* src = "crypto_accelerator.v:1108" *) _T_848;
  assign _T_852 = _T_769 ^ (* src = "crypto_accelerator.v:1109" *) _T_813;
  assign _T_853 = _T_801 ^ (* src = "crypto_accelerator.v:1110" *) _T_850;
  assign _T_856 = _T_821 ^ (* src = "crypto_accelerator.v:1112" *) _T_844;
  assign _T_857 = _T_801 ^ (* src = "crypto_accelerator.v:1113" *) _T_856;
  assign _T_859 = _T_811 ^ (* src = "crypto_accelerator.v:1114" *) _T_852;
  assign _T_860 = _T_801 ^ (* src = "crypto_accelerator.v:1115" *) _T_859;
  assign _T_886 = matrix_0_3[1] ^ (* src = "crypto_accelerator.v:1118" *) matrix_0_3[3];
  assign _T_888 = matrix_0_3[4] ^ (* src = "crypto_accelerator.v:1119" *) matrix_0_3[7];
  assign _T_890 = matrix_0_3[6] ^ (* src = "crypto_accelerator.v:1120" *) matrix_0_3[5];
  assign _T_892 = matrix_0_3[0] ^ (* src = "crypto_accelerator.v:1121" *) _T_890;
  assign _T_894 = _T_886 ^ (* src = "crypto_accelerator.v:1122" *) _T_888;
  assign _T_896 = matrix_0_3[6] ^ (* src = "crypto_accelerator.v:1123" *) matrix_0_3[2];
  assign _T_898 = matrix_0_3[7] ^ (* src = "crypto_accelerator.v:1124" *) matrix_0_3[1];
  assign _T_900 = _T_886 ^ (* src = "crypto_accelerator.v:1125" *) _T_896;
  assign _T_902 = matrix_0_3[1] ^ (* src = "crypto_accelerator.v:1126" *) _T_892;
  assign _T_904 = matrix_0_3[4] ^ (* src = "crypto_accelerator.v:1127" *) _T_892;
  assign _T_906 = matrix_0_3[0] ^ (* src = "crypto_accelerator.v:1128" *) _T_894;
  assign _T_908 = _T_894 ^ (* src = "crypto_accelerator.v:1129" *) _T_896;
  assign _T_910 = matrix_0_3[5] ^ (* src = "crypto_accelerator.v:1130" *) matrix_0_3[2];
  assign _T_912 = _T_890 ^ (* src = "crypto_accelerator.v:1131" *) _T_894;
  assign _T_914 = matrix_0_3[2] ^ (* src = "crypto_accelerator.v:1132" *) _T_898;
  assign _T_916 = matrix_0_3[7] ^ (* src = "crypto_accelerator.v:1133" *) matrix_0_3[2];
  assign _T_918 = matrix_0_3[0] ^ (* src = "crypto_accelerator.v:1134" *) _T_900;
  assign _T_920 = matrix_0_3[1] ^ (* src = "crypto_accelerator.v:1135" *) matrix_0_3[2];
  assign _T_922 = _T_888 ^ (* src = "crypto_accelerator.v:1136" *) _T_920;
  assign _T_924 = _T_892 ^ (* src = "crypto_accelerator.v:1137" *) _T_914;
  assign _T_926 = _T_886 ^ (* src = "crypto_accelerator.v:1138" *) _T_910;
  assign _T_928 = matrix_0_3[7] ^ (* src = "crypto_accelerator.v:1139" *) _T_892;
  assign _T_930 = _T_926 ^ (* src = "crypto_accelerator.v:1140" *) _T_894;
  assign _T_932 = _T_926 ^ (* src = "crypto_accelerator.v:1141" *) _T_898;
  assign _T_934 = _T_898 ^ (* src = "crypto_accelerator.v:1142" *) _T_922;
  assign _T_936 = _T_916 ^ (* src = "crypto_accelerator.v:1143" *) _T_912;
  assign _T_938 = _T_928 ^ (* src = "crypto_accelerator.v:1144" *) _T_918;
  assign _T_944 = _T_908 ^ (* src = "crypto_accelerator.v:1147" *) _T_940;
  assign _T_948 = _T_946 ^ (* src = "crypto_accelerator.v:1149" *) _T_940;
  assign _T_954 = _T_932 ^ (* src = "crypto_accelerator.v:1152" *) _T_950;
  assign _T_958 = _T_956 ^ (* src = "crypto_accelerator.v:1154" *) _T_950;
  assign _T_964 = _T_962 ^ (* src = "crypto_accelerator.v:1157" *) _T_960;
  assign _T_968 = _T_966 ^ (* src = "crypto_accelerator.v:1159" *) _T_960;
  assign _T_970 = _T_944 ^ (* src = "crypto_accelerator.v:1160" *) _T_942;
  assign _T_972 = _T_948 ^ (* src = "crypto_accelerator.v:1161" *) _T_936;
  assign _T_974 = _T_954 ^ (* src = "crypto_accelerator.v:1162" *) _T_952;
  assign _T_976 = _T_958 ^ (* src = "crypto_accelerator.v:1163" *) _T_968;
  assign _T_978 = _T_970 ^ (* src = "crypto_accelerator.v:1164" *) _T_964;
  assign _T_980 = _T_972 ^ (* src = "crypto_accelerator.v:1165" *) _T_968;
  assign _T_982 = _T_974 ^ (* src = "crypto_accelerator.v:1166" *) _T_964;
  assign _T_984 = _T_976 ^ (* src = "crypto_accelerator.v:1167" *) _T_938;
  assign _T_986 = _T_982 ^ (* src = "crypto_accelerator.v:1168" *) _T_984;
  assign _T_990 = _T_980 ^ (* src = "crypto_accelerator.v:1170" *) _T_988;
  assign _T_992 = _T_978 ^ (* src = "crypto_accelerator.v:1171" *) _T_980;
  assign _T_994 = _T_984 ^ (* src = "crypto_accelerator.v:1172" *) _T_988;
  assign _T_1004 = _T_992 ^ (* src = "crypto_accelerator.v:1177" *) _T_988;
  assign _T_1010 = _T_986 ^ (* src = "crypto_accelerator.v:1180" *) _T_988;
  assign _T_1012 = _T_980 ^ (* src = "crypto_accelerator.v:1181" *) _T_996;
  assign _T_1014 = _T_1002 ^ (* src = "crypto_accelerator.v:1182" *) _T_1004;
  assign _T_1016 = _T_984 ^ (* src = "crypto_accelerator.v:1183" *) _T_998;
  assign _T_1018 = _T_1008 ^ (* src = "crypto_accelerator.v:1184" *) _T_1010;
  assign _T_1020 = _T_1014 ^ (* src = "crypto_accelerator.v:1185" *) _T_1018;
  assign _T_1022 = _T_1012 ^ (* src = "crypto_accelerator.v:1186" *) _T_1016;
  assign _T_1024 = _T_1012 ^ (* src = "crypto_accelerator.v:1187" *) _T_1014;
  assign _T_1026 = _T_1016 ^ (* src = "crypto_accelerator.v:1188" *) _T_1018;
  assign _T_1028 = _T_1022 ^ (* src = "crypto_accelerator.v:1189" *) _T_1020;
  assign _T_1066 = _T_1060 ^ (* src = "crypto_accelerator.v:1208" *) _T_1062;
  assign _T_1068 = _T_1038 ^ (* src = "crypto_accelerator.v:1209" *) _T_1050;
  assign _T_1070 = _T_1044 ^ (* src = "crypto_accelerator.v:1210" *) _T_1066;
  assign _T_1072 = _T_1048 ^ (* src = "crypto_accelerator.v:1211" *) _T_1068;
  assign _T_1074 = _T_1034 ^ (* src = "crypto_accelerator.v:1212" *) _T_1054;
  assign _T_1076 = _T_1030 ^ (* src = "crypto_accelerator.v:1213" *) _T_1036;
  assign _T_1078 = _T_1066 ^ (* src = "crypto_accelerator.v:1214" *) _T_1076;
  assign _T_1080 = _T_1032 ^ (* src = "crypto_accelerator.v:1215" *) _T_1072;
  assign _T_1082 = _T_1030 ^ (* src = "crypto_accelerator.v:1216" *) _T_1042;
  assign _T_1084 = _T_1040 ^ (* src = "crypto_accelerator.v:1217" *) _T_1056;
  assign _T_1086 = _T_1046 ^ (* src = "crypto_accelerator.v:1218" *) _T_1058;
  assign _T_1088 = _T_1034 ^ (* src = "crypto_accelerator.v:1219" *) _T_1080;
  assign _T_1090 = _T_1074 ^ (* src = "crypto_accelerator.v:1220" *) _T_1086;
  assign _T_1092 = _T_1052 ^ (* src = "crypto_accelerator.v:1221" *) _T_1068;
  assign _T_1094 = _T_1036 ^ (* src = "crypto_accelerator.v:1222" *) _T_1042;
  assign _T_1096 = _T_1072 ^ (* src = "crypto_accelerator.v:1223" *) _T_1094;
  assign _T_1098 = _T_1064 ^ (* src = "crypto_accelerator.v:1224" *) _T_1090;
  assign _T_1100 = _T_1060 ^ (* src = "crypto_accelerator.v:1225" *) _T_1082;
  assign _T_1102 = _T_1074 ^ (* src = "crypto_accelerator.v:1226" *) _T_1084;
  assign _T_1103 = _T_1070 ^ (* src = "crypto_accelerator.v:1227" *) _T_1096;
  assign _T_1104 = _T_1098 ^ (* src = "crypto_accelerator.v:1228" *) _T_1100;
  assign _T_1107 = _T_1040 ^ (* src = "crypto_accelerator.v:1230" *) _T_1066;
  assign _T_1108 = _T_1078 ^ (* src = "crypto_accelerator.v:1231" *) _T_1080;
  assign _T_1109 = _T_1088 ^ (* src = "crypto_accelerator.v:1232" *) _T_1107;
  assign _T_1111 = _T_1038 ^ (* src = "crypto_accelerator.v:1233" *) _T_1054;
  assign _T_1113 = _T_1076 ^ (* src = "crypto_accelerator.v:1234" *) _T_1092;
  assign _T_1114 = _T_1078 ^ (* src = "crypto_accelerator.v:1235" *) _T_1102;
  assign _T_1117 = _T_1046 ^ (* src = "crypto_accelerator.v:1237" *) _T_1084;
  assign _T_1119 = _T_1111 ^ (* src = "crypto_accelerator.v:1238" *) _T_1117;
  assign _T_1121 = _T_1038 ^ (* src = "crypto_accelerator.v:1239" *) _T_1082;
  assign _T_1122 = _T_1070 ^ (* src = "crypto_accelerator.v:1240" *) _T_1119;
  assign _T_1125 = _T_1090 ^ (* src = "crypto_accelerator.v:1242" *) _T_1113;
  assign _T_1126 = _T_1070 ^ (* src = "crypto_accelerator.v:1243" *) _T_1125;
  assign _T_1128 = _T_1080 ^ (* src = "crypto_accelerator.v:1244" *) _T_1121;
  assign _T_1129 = _T_1070 ^ (* src = "crypto_accelerator.v:1245" *) _T_1128;
  assign _T_1156 = matrix_1_0[1] ^ (* src = "crypto_accelerator.v:1248" *) matrix_1_0[3];
  assign _T_1158 = matrix_1_0[4] ^ (* src = "crypto_accelerator.v:1249" *) matrix_1_0[7];
  assign _T_1160 = matrix_1_0[6] ^ (* src = "crypto_accelerator.v:1250" *) matrix_1_0[5];
  assign _T_1162 = matrix_1_0[0] ^ (* src = "crypto_accelerator.v:1251" *) _T_1160;
  assign _T_1164 = _T_1156 ^ (* src = "crypto_accelerator.v:1252" *) _T_1158;
  assign _T_1166 = matrix_1_0[6] ^ (* src = "crypto_accelerator.v:1253" *) matrix_1_0[2];
  assign _T_1168 = matrix_1_0[7] ^ (* src = "crypto_accelerator.v:1254" *) matrix_1_0[1];
  assign _T_1170 = _T_1156 ^ (* src = "crypto_accelerator.v:1255" *) _T_1166;
  assign _T_1172 = matrix_1_0[1] ^ (* src = "crypto_accelerator.v:1256" *) _T_1162;
  assign _T_1174 = matrix_1_0[4] ^ (* src = "crypto_accelerator.v:1257" *) _T_1162;
  assign _T_1176 = matrix_1_0[0] ^ (* src = "crypto_accelerator.v:1258" *) _T_1164;
  assign _T_1178 = _T_1164 ^ (* src = "crypto_accelerator.v:1259" *) _T_1166;
  assign _T_1180 = matrix_1_0[5] ^ (* src = "crypto_accelerator.v:1260" *) matrix_1_0[2];
  assign _T_1182 = _T_1160 ^ (* src = "crypto_accelerator.v:1261" *) _T_1164;
  assign _T_1184 = matrix_1_0[2] ^ (* src = "crypto_accelerator.v:1262" *) _T_1168;
  assign _T_1186 = matrix_1_0[7] ^ (* src = "crypto_accelerator.v:1263" *) matrix_1_0[2];
  assign _T_1188 = matrix_1_0[0] ^ (* src = "crypto_accelerator.v:1264" *) _T_1170;
  assign _T_1190 = matrix_1_0[1] ^ (* src = "crypto_accelerator.v:1265" *) matrix_1_0[2];
  assign _T_1192 = _T_1158 ^ (* src = "crypto_accelerator.v:1266" *) _T_1190;
  assign _T_1194 = _T_1162 ^ (* src = "crypto_accelerator.v:1267" *) _T_1184;
  assign _T_1196 = _T_1156 ^ (* src = "crypto_accelerator.v:1268" *) _T_1180;
  assign _T_1198 = matrix_1_0[7] ^ (* src = "crypto_accelerator.v:1269" *) _T_1162;
  assign _T_1200 = _T_1196 ^ (* src = "crypto_accelerator.v:1270" *) _T_1164;
  assign _T_1202 = _T_1196 ^ (* src = "crypto_accelerator.v:1271" *) _T_1168;
  assign _T_1204 = _T_1168 ^ (* src = "crypto_accelerator.v:1272" *) _T_1192;
  assign _T_1206 = _T_1186 ^ (* src = "crypto_accelerator.v:1273" *) _T_1182;
  assign _T_1208 = _T_1198 ^ (* src = "crypto_accelerator.v:1274" *) _T_1188;
  assign _T_1214 = _T_1178 ^ (* src = "crypto_accelerator.v:1277" *) _T_1210;
  assign _T_1218 = _T_1216 ^ (* src = "crypto_accelerator.v:1279" *) _T_1210;
  assign _T_1224 = _T_1202 ^ (* src = "crypto_accelerator.v:1282" *) _T_1220;
  assign _T_1228 = _T_1226 ^ (* src = "crypto_accelerator.v:1284" *) _T_1220;
  assign _T_1234 = _T_1232 ^ (* src = "crypto_accelerator.v:1287" *) _T_1230;
  assign _T_1238 = _T_1236 ^ (* src = "crypto_accelerator.v:1289" *) _T_1230;
  assign _T_1240 = _T_1214 ^ (* src = "crypto_accelerator.v:1290" *) _T_1212;
  assign _T_1242 = _T_1218 ^ (* src = "crypto_accelerator.v:1291" *) _T_1206;
  assign _T_1244 = _T_1224 ^ (* src = "crypto_accelerator.v:1292" *) _T_1222;
  assign _T_1246 = _T_1228 ^ (* src = "crypto_accelerator.v:1293" *) _T_1238;
  assign _T_1248 = _T_1240 ^ (* src = "crypto_accelerator.v:1294" *) _T_1234;
  assign _T_1250 = _T_1242 ^ (* src = "crypto_accelerator.v:1295" *) _T_1238;
  assign _T_1252 = _T_1244 ^ (* src = "crypto_accelerator.v:1296" *) _T_1234;
  assign _T_1254 = _T_1246 ^ (* src = "crypto_accelerator.v:1297" *) _T_1208;
  assign _T_1256 = _T_1252 ^ (* src = "crypto_accelerator.v:1298" *) _T_1254;
  assign _T_1260 = _T_1250 ^ (* src = "crypto_accelerator.v:1300" *) _T_1258;
  assign _T_1262 = _T_1248 ^ (* src = "crypto_accelerator.v:1301" *) _T_1250;
  assign _T_1264 = _T_1254 ^ (* src = "crypto_accelerator.v:1302" *) _T_1258;
  assign _T_1274 = _T_1262 ^ (* src = "crypto_accelerator.v:1307" *) _T_1258;
  assign _T_1280 = _T_1256 ^ (* src = "crypto_accelerator.v:1310" *) _T_1258;
  assign _T_1282 = _T_1250 ^ (* src = "crypto_accelerator.v:1311" *) _T_1266;
  assign _T_1284 = _T_1272 ^ (* src = "crypto_accelerator.v:1312" *) _T_1274;
  assign _T_1286 = _T_1254 ^ (* src = "crypto_accelerator.v:1313" *) _T_1268;
  assign _T_1288 = _T_1278 ^ (* src = "crypto_accelerator.v:1314" *) _T_1280;
  assign _T_1290 = _T_1284 ^ (* src = "crypto_accelerator.v:1315" *) _T_1288;
  assign _T_1292 = _T_1282 ^ (* src = "crypto_accelerator.v:1316" *) _T_1286;
  assign _T_1294 = _T_1282 ^ (* src = "crypto_accelerator.v:1317" *) _T_1284;
  assign _T_1296 = _T_1286 ^ (* src = "crypto_accelerator.v:1318" *) _T_1288;
  assign _T_1298 = _T_1292 ^ (* src = "crypto_accelerator.v:1319" *) _T_1290;
  assign _T_1336 = _T_1330 ^ (* src = "crypto_accelerator.v:1338" *) _T_1332;
  assign _T_1338 = _T_1308 ^ (* src = "crypto_accelerator.v:1339" *) _T_1320;
  assign _T_1340 = _T_1314 ^ (* src = "crypto_accelerator.v:1340" *) _T_1336;
  assign _T_1342 = _T_1318 ^ (* src = "crypto_accelerator.v:1341" *) _T_1338;
  assign _T_1344 = _T_1304 ^ (* src = "crypto_accelerator.v:1342" *) _T_1324;
  assign _T_1346 = _T_1300 ^ (* src = "crypto_accelerator.v:1343" *) _T_1306;
  assign _T_1348 = _T_1336 ^ (* src = "crypto_accelerator.v:1344" *) _T_1346;
  assign _T_1350 = _T_1302 ^ (* src = "crypto_accelerator.v:1345" *) _T_1342;
  assign _T_1352 = _T_1300 ^ (* src = "crypto_accelerator.v:1346" *) _T_1312;
  assign _T_1354 = _T_1310 ^ (* src = "crypto_accelerator.v:1347" *) _T_1326;
  assign _T_1356 = _T_1316 ^ (* src = "crypto_accelerator.v:1348" *) _T_1328;
  assign _T_1358 = _T_1304 ^ (* src = "crypto_accelerator.v:1349" *) _T_1350;
  assign _T_1360 = _T_1344 ^ (* src = "crypto_accelerator.v:1350" *) _T_1356;
  assign _T_1362 = _T_1322 ^ (* src = "crypto_accelerator.v:1351" *) _T_1338;
  assign _T_1364 = _T_1306 ^ (* src = "crypto_accelerator.v:1352" *) _T_1312;
  assign _T_1366 = _T_1342 ^ (* src = "crypto_accelerator.v:1353" *) _T_1364;
  assign _T_1368 = _T_1334 ^ (* src = "crypto_accelerator.v:1354" *) _T_1360;
  assign _T_1370 = _T_1330 ^ (* src = "crypto_accelerator.v:1355" *) _T_1352;
  assign _T_1372 = _T_1344 ^ (* src = "crypto_accelerator.v:1356" *) _T_1354;
  assign _T_1373 = _T_1340 ^ (* src = "crypto_accelerator.v:1357" *) _T_1366;
  assign _T_1374 = _T_1368 ^ (* src = "crypto_accelerator.v:1358" *) _T_1370;
  assign _T_1377 = _T_1310 ^ (* src = "crypto_accelerator.v:1360" *) _T_1336;
  assign _T_1378 = _T_1348 ^ (* src = "crypto_accelerator.v:1361" *) _T_1350;
  assign _T_1379 = _T_1358 ^ (* src = "crypto_accelerator.v:1362" *) _T_1377;
  assign _T_1381 = _T_1308 ^ (* src = "crypto_accelerator.v:1363" *) _T_1324;
  assign _T_1383 = _T_1346 ^ (* src = "crypto_accelerator.v:1364" *) _T_1362;
  assign _T_1384 = _T_1348 ^ (* src = "crypto_accelerator.v:1365" *) _T_1372;
  assign _T_1387 = _T_1316 ^ (* src = "crypto_accelerator.v:1367" *) _T_1354;
  assign _T_1389 = _T_1381 ^ (* src = "crypto_accelerator.v:1368" *) _T_1387;
  assign _T_1391 = _T_1308 ^ (* src = "crypto_accelerator.v:1369" *) _T_1352;
  assign _T_1392 = _T_1340 ^ (* src = "crypto_accelerator.v:1370" *) _T_1389;
  assign _T_1395 = _T_1360 ^ (* src = "crypto_accelerator.v:1372" *) _T_1383;
  assign _T_1396 = _T_1340 ^ (* src = "crypto_accelerator.v:1373" *) _T_1395;
  assign _T_1398 = _T_1350 ^ (* src = "crypto_accelerator.v:1374" *) _T_1391;
  assign _T_1399 = _T_1340 ^ (* src = "crypto_accelerator.v:1375" *) _T_1398;
  assign _T_1425 = matrix_1_1[1] ^ (* src = "crypto_accelerator.v:1378" *) matrix_1_1[3];
  assign _T_1427 = matrix_1_1[4] ^ (* src = "crypto_accelerator.v:1379" *) matrix_1_1[7];
  assign _T_1429 = matrix_1_1[6] ^ (* src = "crypto_accelerator.v:1380" *) matrix_1_1[5];
  assign _T_1431 = matrix_1_1[0] ^ (* src = "crypto_accelerator.v:1381" *) _T_1429;
  assign _T_1433 = _T_1425 ^ (* src = "crypto_accelerator.v:1382" *) _T_1427;
  assign _T_1435 = matrix_1_1[6] ^ (* src = "crypto_accelerator.v:1383" *) matrix_1_1[2];
  assign _T_1437 = matrix_1_1[7] ^ (* src = "crypto_accelerator.v:1384" *) matrix_1_1[1];
  assign _T_1439 = _T_1425 ^ (* src = "crypto_accelerator.v:1385" *) _T_1435;
  assign _T_1441 = matrix_1_1[1] ^ (* src = "crypto_accelerator.v:1386" *) _T_1431;
  assign _T_1443 = matrix_1_1[4] ^ (* src = "crypto_accelerator.v:1387" *) _T_1431;
  assign _T_1445 = matrix_1_1[0] ^ (* src = "crypto_accelerator.v:1388" *) _T_1433;
  assign _T_1447 = _T_1433 ^ (* src = "crypto_accelerator.v:1389" *) _T_1435;
  assign _T_1449 = matrix_1_1[5] ^ (* src = "crypto_accelerator.v:1390" *) matrix_1_1[2];
  assign _T_1451 = _T_1429 ^ (* src = "crypto_accelerator.v:1391" *) _T_1433;
  assign _T_1453 = matrix_1_1[2] ^ (* src = "crypto_accelerator.v:1392" *) _T_1437;
  assign _T_1455 = matrix_1_1[7] ^ (* src = "crypto_accelerator.v:1393" *) matrix_1_1[2];
  assign _T_1457 = matrix_1_1[0] ^ (* src = "crypto_accelerator.v:1394" *) _T_1439;
  assign _T_1459 = matrix_1_1[1] ^ (* src = "crypto_accelerator.v:1395" *) matrix_1_1[2];
  assign _T_1461 = _T_1427 ^ (* src = "crypto_accelerator.v:1396" *) _T_1459;
  assign _T_1463 = _T_1431 ^ (* src = "crypto_accelerator.v:1397" *) _T_1453;
  assign _T_1465 = _T_1425 ^ (* src = "crypto_accelerator.v:1398" *) _T_1449;
  assign _T_1467 = matrix_1_1[7] ^ (* src = "crypto_accelerator.v:1399" *) _T_1431;
  assign _T_1469 = _T_1465 ^ (* src = "crypto_accelerator.v:1400" *) _T_1433;
  assign _T_1471 = _T_1465 ^ (* src = "crypto_accelerator.v:1401" *) _T_1437;
  assign _T_1473 = _T_1437 ^ (* src = "crypto_accelerator.v:1402" *) _T_1461;
  assign _T_1475 = _T_1455 ^ (* src = "crypto_accelerator.v:1403" *) _T_1451;
  assign _T_1477 = _T_1467 ^ (* src = "crypto_accelerator.v:1404" *) _T_1457;
  assign _T_1483 = _T_1447 ^ (* src = "crypto_accelerator.v:1407" *) _T_1479;
  assign _T_1487 = _T_1485 ^ (* src = "crypto_accelerator.v:1409" *) _T_1479;
  assign _T_1493 = _T_1471 ^ (* src = "crypto_accelerator.v:1412" *) _T_1489;
  assign _T_1497 = _T_1495 ^ (* src = "crypto_accelerator.v:1414" *) _T_1489;
  assign _T_1503 = _T_1501 ^ (* src = "crypto_accelerator.v:1417" *) _T_1499;
  assign _T_1507 = _T_1505 ^ (* src = "crypto_accelerator.v:1419" *) _T_1499;
  assign _T_1509 = _T_1483 ^ (* src = "crypto_accelerator.v:1420" *) _T_1481;
  assign _T_1511 = _T_1487 ^ (* src = "crypto_accelerator.v:1421" *) _T_1475;
  assign _T_1513 = _T_1493 ^ (* src = "crypto_accelerator.v:1422" *) _T_1491;
  assign _T_1515 = _T_1497 ^ (* src = "crypto_accelerator.v:1423" *) _T_1507;
  assign _T_1517 = _T_1509 ^ (* src = "crypto_accelerator.v:1424" *) _T_1503;
  assign _T_1519 = _T_1511 ^ (* src = "crypto_accelerator.v:1425" *) _T_1507;
  assign _T_1521 = _T_1513 ^ (* src = "crypto_accelerator.v:1426" *) _T_1503;
  assign _T_1523 = _T_1515 ^ (* src = "crypto_accelerator.v:1427" *) _T_1477;
  assign _T_1525 = _T_1521 ^ (* src = "crypto_accelerator.v:1428" *) _T_1523;
  assign _T_1529 = _T_1519 ^ (* src = "crypto_accelerator.v:1430" *) _T_1527;
  assign _T_1531 = _T_1517 ^ (* src = "crypto_accelerator.v:1431" *) _T_1519;
  assign _T_1533 = _T_1523 ^ (* src = "crypto_accelerator.v:1432" *) _T_1527;
  assign _T_1543 = _T_1531 ^ (* src = "crypto_accelerator.v:1437" *) _T_1527;
  assign _T_1549 = _T_1525 ^ (* src = "crypto_accelerator.v:1440" *) _T_1527;
  assign _T_1551 = _T_1519 ^ (* src = "crypto_accelerator.v:1441" *) _T_1535;
  assign _T_1553 = _T_1541 ^ (* src = "crypto_accelerator.v:1442" *) _T_1543;
  assign _T_1555 = _T_1523 ^ (* src = "crypto_accelerator.v:1443" *) _T_1537;
  assign _T_1557 = _T_1547 ^ (* src = "crypto_accelerator.v:1444" *) _T_1549;
  assign _T_1559 = _T_1553 ^ (* src = "crypto_accelerator.v:1445" *) _T_1557;
  assign _T_1561 = _T_1551 ^ (* src = "crypto_accelerator.v:1446" *) _T_1555;
  assign _T_1563 = _T_1551 ^ (* src = "crypto_accelerator.v:1447" *) _T_1553;
  assign _T_1565 = _T_1555 ^ (* src = "crypto_accelerator.v:1448" *) _T_1557;
  assign _T_1567 = _T_1561 ^ (* src = "crypto_accelerator.v:1449" *) _T_1559;
  assign _T_1605 = _T_1599 ^ (* src = "crypto_accelerator.v:1468" *) _T_1601;
  assign _T_1607 = _T_1577 ^ (* src = "crypto_accelerator.v:1469" *) _T_1589;
  assign _T_1609 = _T_1583 ^ (* src = "crypto_accelerator.v:1470" *) _T_1605;
  assign _T_1611 = _T_1587 ^ (* src = "crypto_accelerator.v:1471" *) _T_1607;
  assign _T_1613 = _T_1573 ^ (* src = "crypto_accelerator.v:1472" *) _T_1593;
  assign _T_1615 = _T_1569 ^ (* src = "crypto_accelerator.v:1473" *) _T_1575;
  assign _T_1617 = _T_1605 ^ (* src = "crypto_accelerator.v:1474" *) _T_1615;
  assign _T_1619 = _T_1571 ^ (* src = "crypto_accelerator.v:1475" *) _T_1611;
  assign _T_1621 = _T_1569 ^ (* src = "crypto_accelerator.v:1476" *) _T_1581;
  assign _T_1623 = _T_1579 ^ (* src = "crypto_accelerator.v:1477" *) _T_1595;
  assign _T_1625 = _T_1585 ^ (* src = "crypto_accelerator.v:1478" *) _T_1597;
  assign _T_1627 = _T_1573 ^ (* src = "crypto_accelerator.v:1479" *) _T_1619;
  assign _T_1629 = _T_1613 ^ (* src = "crypto_accelerator.v:1480" *) _T_1625;
  assign _T_1631 = _T_1591 ^ (* src = "crypto_accelerator.v:1481" *) _T_1607;
  assign _T_1633 = _T_1575 ^ (* src = "crypto_accelerator.v:1482" *) _T_1581;
  assign _T_1635 = _T_1611 ^ (* src = "crypto_accelerator.v:1483" *) _T_1633;
  assign _T_1637 = _T_1603 ^ (* src = "crypto_accelerator.v:1484" *) _T_1629;
  assign _T_1639 = _T_1599 ^ (* src = "crypto_accelerator.v:1485" *) _T_1621;
  assign _T_1641 = _T_1613 ^ (* src = "crypto_accelerator.v:1486" *) _T_1623;
  assign _T_1642 = _T_1609 ^ (* src = "crypto_accelerator.v:1487" *) _T_1635;
  assign _T_1643 = _T_1637 ^ (* src = "crypto_accelerator.v:1488" *) _T_1639;
  assign _T_1646 = _T_1579 ^ (* src = "crypto_accelerator.v:1490" *) _T_1605;
  assign _T_1647 = _T_1617 ^ (* src = "crypto_accelerator.v:1491" *) _T_1619;
  assign _T_1648 = _T_1627 ^ (* src = "crypto_accelerator.v:1492" *) _T_1646;
  assign _T_1650 = _T_1577 ^ (* src = "crypto_accelerator.v:1493" *) _T_1593;
  assign _T_1652 = _T_1615 ^ (* src = "crypto_accelerator.v:1494" *) _T_1631;
  assign _T_1653 = _T_1617 ^ (* src = "crypto_accelerator.v:1495" *) _T_1641;
  assign _T_1656 = _T_1585 ^ (* src = "crypto_accelerator.v:1497" *) _T_1623;
  assign _T_1658 = _T_1650 ^ (* src = "crypto_accelerator.v:1498" *) _T_1656;
  assign _T_1660 = _T_1577 ^ (* src = "crypto_accelerator.v:1499" *) _T_1621;
  assign _T_1661 = _T_1609 ^ (* src = "crypto_accelerator.v:1500" *) _T_1658;
  assign _T_1664 = _T_1629 ^ (* src = "crypto_accelerator.v:1502" *) _T_1652;
  assign _T_1665 = _T_1609 ^ (* src = "crypto_accelerator.v:1503" *) _T_1664;
  assign _T_1667 = _T_1619 ^ (* src = "crypto_accelerator.v:1504" *) _T_1660;
  assign _T_1668 = _T_1609 ^ (* src = "crypto_accelerator.v:1505" *) _T_1667;
  assign _T_1694 = matrix_1_2[1] ^ (* src = "crypto_accelerator.v:1508" *) matrix_1_2[3];
  assign _T_1696 = matrix_1_2[4] ^ (* src = "crypto_accelerator.v:1509" *) matrix_1_2[7];
  assign _T_1698 = matrix_1_2[6] ^ (* src = "crypto_accelerator.v:1510" *) matrix_1_2[5];
  assign _T_1700 = matrix_1_2[0] ^ (* src = "crypto_accelerator.v:1511" *) _T_1698;
  assign _T_1702 = _T_1694 ^ (* src = "crypto_accelerator.v:1512" *) _T_1696;
  assign _T_1704 = matrix_1_2[6] ^ (* src = "crypto_accelerator.v:1513" *) matrix_1_2[2];
  assign _T_1706 = matrix_1_2[7] ^ (* src = "crypto_accelerator.v:1514" *) matrix_1_2[1];
  assign _T_1708 = _T_1694 ^ (* src = "crypto_accelerator.v:1515" *) _T_1704;
  assign _T_1710 = matrix_1_2[1] ^ (* src = "crypto_accelerator.v:1516" *) _T_1700;
  assign _T_1712 = matrix_1_2[4] ^ (* src = "crypto_accelerator.v:1517" *) _T_1700;
  assign _T_1714 = matrix_1_2[0] ^ (* src = "crypto_accelerator.v:1518" *) _T_1702;
  assign _T_1716 = _T_1702 ^ (* src = "crypto_accelerator.v:1519" *) _T_1704;
  assign _T_1718 = matrix_1_2[5] ^ (* src = "crypto_accelerator.v:1520" *) matrix_1_2[2];
  assign _T_1720 = _T_1698 ^ (* src = "crypto_accelerator.v:1521" *) _T_1702;
  assign _T_1722 = matrix_1_2[2] ^ (* src = "crypto_accelerator.v:1522" *) _T_1706;
  assign _T_1724 = matrix_1_2[7] ^ (* src = "crypto_accelerator.v:1523" *) matrix_1_2[2];
  assign _T_1726 = matrix_1_2[0] ^ (* src = "crypto_accelerator.v:1524" *) _T_1708;
  assign _T_1728 = matrix_1_2[1] ^ (* src = "crypto_accelerator.v:1525" *) matrix_1_2[2];
  assign _T_1730 = _T_1696 ^ (* src = "crypto_accelerator.v:1526" *) _T_1728;
  assign _T_1732 = _T_1700 ^ (* src = "crypto_accelerator.v:1527" *) _T_1722;
  assign _T_1734 = _T_1694 ^ (* src = "crypto_accelerator.v:1528" *) _T_1718;
  assign _T_1736 = matrix_1_2[7] ^ (* src = "crypto_accelerator.v:1529" *) _T_1700;
  assign _T_1738 = _T_1734 ^ (* src = "crypto_accelerator.v:1530" *) _T_1702;
  assign _T_1740 = _T_1734 ^ (* src = "crypto_accelerator.v:1531" *) _T_1706;
  assign _T_1742 = _T_1706 ^ (* src = "crypto_accelerator.v:1532" *) _T_1730;
  assign _T_1744 = _T_1724 ^ (* src = "crypto_accelerator.v:1533" *) _T_1720;
  assign _T_1746 = _T_1736 ^ (* src = "crypto_accelerator.v:1534" *) _T_1726;
  assign _T_1752 = _T_1716 ^ (* src = "crypto_accelerator.v:1537" *) _T_1748;
  assign _T_1756 = _T_1754 ^ (* src = "crypto_accelerator.v:1539" *) _T_1748;
  assign _T_1762 = _T_1740 ^ (* src = "crypto_accelerator.v:1542" *) _T_1758;
  assign _T_1766 = _T_1764 ^ (* src = "crypto_accelerator.v:1544" *) _T_1758;
  assign _T_1772 = _T_1770 ^ (* src = "crypto_accelerator.v:1547" *) _T_1768;
  assign _T_1776 = _T_1774 ^ (* src = "crypto_accelerator.v:1549" *) _T_1768;
  assign _T_1778 = _T_1752 ^ (* src = "crypto_accelerator.v:1550" *) _T_1750;
  assign _T_1780 = _T_1756 ^ (* src = "crypto_accelerator.v:1551" *) _T_1744;
  assign _T_1782 = _T_1762 ^ (* src = "crypto_accelerator.v:1552" *) _T_1760;
  assign _T_1784 = _T_1766 ^ (* src = "crypto_accelerator.v:1553" *) _T_1776;
  assign _T_1786 = _T_1778 ^ (* src = "crypto_accelerator.v:1554" *) _T_1772;
  assign _T_1788 = _T_1780 ^ (* src = "crypto_accelerator.v:1555" *) _T_1776;
  assign _T_1790 = _T_1782 ^ (* src = "crypto_accelerator.v:1556" *) _T_1772;
  assign _T_1792 = _T_1784 ^ (* src = "crypto_accelerator.v:1557" *) _T_1746;
  assign _T_1794 = _T_1790 ^ (* src = "crypto_accelerator.v:1558" *) _T_1792;
  assign _T_1798 = _T_1788 ^ (* src = "crypto_accelerator.v:1560" *) _T_1796;
  assign _T_1800 = _T_1786 ^ (* src = "crypto_accelerator.v:1561" *) _T_1788;
  assign _T_1802 = _T_1792 ^ (* src = "crypto_accelerator.v:1562" *) _T_1796;
  assign _T_1812 = _T_1800 ^ (* src = "crypto_accelerator.v:1567" *) _T_1796;
  assign _T_1818 = _T_1794 ^ (* src = "crypto_accelerator.v:1570" *) _T_1796;
  assign _T_1820 = _T_1788 ^ (* src = "crypto_accelerator.v:1571" *) _T_1804;
  assign _T_1822 = _T_1810 ^ (* src = "crypto_accelerator.v:1572" *) _T_1812;
  assign _T_1824 = _T_1792 ^ (* src = "crypto_accelerator.v:1573" *) _T_1806;
  assign _T_1826 = _T_1816 ^ (* src = "crypto_accelerator.v:1574" *) _T_1818;
  assign _T_1828 = _T_1822 ^ (* src = "crypto_accelerator.v:1575" *) _T_1826;
  assign _T_1830 = _T_1820 ^ (* src = "crypto_accelerator.v:1576" *) _T_1824;
  assign _T_1832 = _T_1820 ^ (* src = "crypto_accelerator.v:1577" *) _T_1822;
  assign _T_1834 = _T_1824 ^ (* src = "crypto_accelerator.v:1578" *) _T_1826;
  assign _T_1836 = _T_1830 ^ (* src = "crypto_accelerator.v:1579" *) _T_1828;
  assign _T_1874 = _T_1868 ^ (* src = "crypto_accelerator.v:1598" *) _T_1870;
  assign _T_1876 = _T_1846 ^ (* src = "crypto_accelerator.v:1599" *) _T_1858;
  assign _T_1878 = _T_1852 ^ (* src = "crypto_accelerator.v:1600" *) _T_1874;
  assign _T_1880 = _T_1856 ^ (* src = "crypto_accelerator.v:1601" *) _T_1876;
  assign _T_1882 = _T_1842 ^ (* src = "crypto_accelerator.v:1602" *) _T_1862;
  assign _T_1884 = _T_1838 ^ (* src = "crypto_accelerator.v:1603" *) _T_1844;
  assign _T_1886 = _T_1874 ^ (* src = "crypto_accelerator.v:1604" *) _T_1884;
  assign _T_1888 = _T_1840 ^ (* src = "crypto_accelerator.v:1605" *) _T_1880;
  assign _T_1890 = _T_1838 ^ (* src = "crypto_accelerator.v:1606" *) _T_1850;
  assign _T_1892 = _T_1848 ^ (* src = "crypto_accelerator.v:1607" *) _T_1864;
  assign _T_1894 = _T_1854 ^ (* src = "crypto_accelerator.v:1608" *) _T_1866;
  assign _T_1896 = _T_1842 ^ (* src = "crypto_accelerator.v:1609" *) _T_1888;
  assign _T_1898 = _T_1882 ^ (* src = "crypto_accelerator.v:1610" *) _T_1894;
  assign _T_1900 = _T_1860 ^ (* src = "crypto_accelerator.v:1611" *) _T_1876;
  assign _T_1902 = _T_1844 ^ (* src = "crypto_accelerator.v:1612" *) _T_1850;
  assign _T_1904 = _T_1880 ^ (* src = "crypto_accelerator.v:1613" *) _T_1902;
  assign _T_1906 = _T_1872 ^ (* src = "crypto_accelerator.v:1614" *) _T_1898;
  assign _T_1908 = _T_1868 ^ (* src = "crypto_accelerator.v:1615" *) _T_1890;
  assign _T_1910 = _T_1882 ^ (* src = "crypto_accelerator.v:1616" *) _T_1892;
  assign _T_1911 = _T_1878 ^ (* src = "crypto_accelerator.v:1617" *) _T_1904;
  assign _T_1912 = _T_1906 ^ (* src = "crypto_accelerator.v:1618" *) _T_1908;
  assign _T_1915 = _T_1848 ^ (* src = "crypto_accelerator.v:1620" *) _T_1874;
  assign _T_1916 = _T_1886 ^ (* src = "crypto_accelerator.v:1621" *) _T_1888;
  assign _T_1917 = _T_1896 ^ (* src = "crypto_accelerator.v:1622" *) _T_1915;
  assign _T_1919 = _T_1846 ^ (* src = "crypto_accelerator.v:1623" *) _T_1862;
  assign _T_1921 = _T_1884 ^ (* src = "crypto_accelerator.v:1624" *) _T_1900;
  assign _T_1922 = _T_1886 ^ (* src = "crypto_accelerator.v:1625" *) _T_1910;
  assign _T_1925 = _T_1854 ^ (* src = "crypto_accelerator.v:1627" *) _T_1892;
  assign _T_1927 = _T_1919 ^ (* src = "crypto_accelerator.v:1628" *) _T_1925;
  assign _T_1929 = _T_1846 ^ (* src = "crypto_accelerator.v:1629" *) _T_1890;
  assign _T_1930 = _T_1878 ^ (* src = "crypto_accelerator.v:1630" *) _T_1927;
  assign _T_1933 = _T_1898 ^ (* src = "crypto_accelerator.v:1632" *) _T_1921;
  assign _T_1934 = _T_1878 ^ (* src = "crypto_accelerator.v:1633" *) _T_1933;
  assign _T_1936 = _T_1888 ^ (* src = "crypto_accelerator.v:1634" *) _T_1929;
  assign _T_1937 = _T_1878 ^ (* src = "crypto_accelerator.v:1635" *) _T_1936;
  assign _T_1963 = matrix_1_3[1] ^ (* src = "crypto_accelerator.v:1638" *) matrix_1_3[3];
  assign _T_1965 = matrix_1_3[4] ^ (* src = "crypto_accelerator.v:1639" *) matrix_1_3[7];
  assign _T_1967 = matrix_1_3[6] ^ (* src = "crypto_accelerator.v:1640" *) matrix_1_3[5];
  assign _T_1969 = matrix_1_3[0] ^ (* src = "crypto_accelerator.v:1641" *) _T_1967;
  assign _T_1971 = _T_1963 ^ (* src = "crypto_accelerator.v:1642" *) _T_1965;
  assign _T_1973 = matrix_1_3[6] ^ (* src = "crypto_accelerator.v:1643" *) matrix_1_3[2];
  assign _T_1975 = matrix_1_3[7] ^ (* src = "crypto_accelerator.v:1644" *) matrix_1_3[1];
  assign _T_1977 = _T_1963 ^ (* src = "crypto_accelerator.v:1645" *) _T_1973;
  assign _T_1979 = matrix_1_3[1] ^ (* src = "crypto_accelerator.v:1646" *) _T_1969;
  assign _T_1981 = matrix_1_3[4] ^ (* src = "crypto_accelerator.v:1647" *) _T_1969;
  assign _T_1983 = matrix_1_3[0] ^ (* src = "crypto_accelerator.v:1648" *) _T_1971;
  assign _T_1985 = _T_1971 ^ (* src = "crypto_accelerator.v:1649" *) _T_1973;
  assign _T_1987 = matrix_1_3[5] ^ (* src = "crypto_accelerator.v:1650" *) matrix_1_3[2];
  assign _T_1989 = _T_1967 ^ (* src = "crypto_accelerator.v:1651" *) _T_1971;
  assign _T_1991 = matrix_1_3[2] ^ (* src = "crypto_accelerator.v:1652" *) _T_1975;
  assign _T_1993 = matrix_1_3[7] ^ (* src = "crypto_accelerator.v:1653" *) matrix_1_3[2];
  assign _T_1995 = matrix_1_3[0] ^ (* src = "crypto_accelerator.v:1654" *) _T_1977;
  assign _T_1997 = matrix_1_3[1] ^ (* src = "crypto_accelerator.v:1655" *) matrix_1_3[2];
  assign _T_1999 = _T_1965 ^ (* src = "crypto_accelerator.v:1656" *) _T_1997;
  assign _T_2001 = _T_1969 ^ (* src = "crypto_accelerator.v:1657" *) _T_1991;
  assign _T_2003 = _T_1963 ^ (* src = "crypto_accelerator.v:1658" *) _T_1987;
  assign _T_2005 = matrix_1_3[7] ^ (* src = "crypto_accelerator.v:1659" *) _T_1969;
  assign _T_2007 = _T_2003 ^ (* src = "crypto_accelerator.v:1660" *) _T_1971;
  assign _T_2009 = _T_2003 ^ (* src = "crypto_accelerator.v:1661" *) _T_1975;
  assign _T_2011 = _T_1975 ^ (* src = "crypto_accelerator.v:1662" *) _T_1999;
  assign _T_2013 = _T_1993 ^ (* src = "crypto_accelerator.v:1663" *) _T_1989;
  assign _T_2015 = _T_2005 ^ (* src = "crypto_accelerator.v:1664" *) _T_1995;
  assign _T_2021 = _T_1985 ^ (* src = "crypto_accelerator.v:1667" *) _T_2017;
  assign _T_2025 = _T_2023 ^ (* src = "crypto_accelerator.v:1669" *) _T_2017;
  assign _T_2031 = _T_2009 ^ (* src = "crypto_accelerator.v:1672" *) _T_2027;
  assign _T_2035 = _T_2033 ^ (* src = "crypto_accelerator.v:1674" *) _T_2027;
  assign _T_2041 = _T_2039 ^ (* src = "crypto_accelerator.v:1677" *) _T_2037;
  assign _T_2045 = _T_2043 ^ (* src = "crypto_accelerator.v:1679" *) _T_2037;
  assign _T_2047 = _T_2021 ^ (* src = "crypto_accelerator.v:1680" *) _T_2019;
  assign _T_2049 = _T_2025 ^ (* src = "crypto_accelerator.v:1681" *) _T_2013;
  assign _T_2051 = _T_2031 ^ (* src = "crypto_accelerator.v:1682" *) _T_2029;
  assign _T_2053 = _T_2035 ^ (* src = "crypto_accelerator.v:1683" *) _T_2045;
  assign _T_2055 = _T_2047 ^ (* src = "crypto_accelerator.v:1684" *) _T_2041;
  assign _T_2057 = _T_2049 ^ (* src = "crypto_accelerator.v:1685" *) _T_2045;
  assign _T_2059 = _T_2051 ^ (* src = "crypto_accelerator.v:1686" *) _T_2041;
  assign _T_2061 = _T_2053 ^ (* src = "crypto_accelerator.v:1687" *) _T_2015;
  assign _T_2063 = _T_2059 ^ (* src = "crypto_accelerator.v:1688" *) _T_2061;
  assign _T_2067 = _T_2057 ^ (* src = "crypto_accelerator.v:1690" *) _T_2065;
  assign _T_2069 = _T_2055 ^ (* src = "crypto_accelerator.v:1691" *) _T_2057;
  assign _T_2071 = _T_2061 ^ (* src = "crypto_accelerator.v:1692" *) _T_2065;
  assign _T_2081 = _T_2069 ^ (* src = "crypto_accelerator.v:1697" *) _T_2065;
  assign _T_2087 = _T_2063 ^ (* src = "crypto_accelerator.v:1700" *) _T_2065;
  assign _T_2089 = _T_2057 ^ (* src = "crypto_accelerator.v:1701" *) _T_2073;
  assign _T_2091 = _T_2079 ^ (* src = "crypto_accelerator.v:1702" *) _T_2081;
  assign _T_2093 = _T_2061 ^ (* src = "crypto_accelerator.v:1703" *) _T_2075;
  assign _T_2095 = _T_2085 ^ (* src = "crypto_accelerator.v:1704" *) _T_2087;
  assign _T_2097 = _T_2091 ^ (* src = "crypto_accelerator.v:1705" *) _T_2095;
  assign _T_2099 = _T_2089 ^ (* src = "crypto_accelerator.v:1706" *) _T_2093;
  assign _T_2101 = _T_2089 ^ (* src = "crypto_accelerator.v:1707" *) _T_2091;
  assign _T_2103 = _T_2093 ^ (* src = "crypto_accelerator.v:1708" *) _T_2095;
  assign _T_2105 = _T_2099 ^ (* src = "crypto_accelerator.v:1709" *) _T_2097;
  assign _T_2143 = _T_2137 ^ (* src = "crypto_accelerator.v:1728" *) _T_2139;
  assign _T_2145 = _T_2115 ^ (* src = "crypto_accelerator.v:1729" *) _T_2127;
  assign _T_2147 = _T_2121 ^ (* src = "crypto_accelerator.v:1730" *) _T_2143;
  assign _T_2149 = _T_2125 ^ (* src = "crypto_accelerator.v:1731" *) _T_2145;
  assign _T_2151 = _T_2111 ^ (* src = "crypto_accelerator.v:1732" *) _T_2131;
  assign _T_2153 = _T_2107 ^ (* src = "crypto_accelerator.v:1733" *) _T_2113;
  assign _T_2155 = _T_2143 ^ (* src = "crypto_accelerator.v:1734" *) _T_2153;
  assign _T_2157 = _T_2109 ^ (* src = "crypto_accelerator.v:1735" *) _T_2149;
  assign _T_2159 = _T_2107 ^ (* src = "crypto_accelerator.v:1736" *) _T_2119;
  assign _T_2161 = _T_2117 ^ (* src = "crypto_accelerator.v:1737" *) _T_2133;
  assign _T_2163 = _T_2123 ^ (* src = "crypto_accelerator.v:1738" *) _T_2135;
  assign _T_2165 = _T_2111 ^ (* src = "crypto_accelerator.v:1739" *) _T_2157;
  assign _T_2167 = _T_2151 ^ (* src = "crypto_accelerator.v:1740" *) _T_2163;
  assign _T_2169 = _T_2129 ^ (* src = "crypto_accelerator.v:1741" *) _T_2145;
  assign _T_2171 = _T_2113 ^ (* src = "crypto_accelerator.v:1742" *) _T_2119;
  assign _T_2173 = _T_2149 ^ (* src = "crypto_accelerator.v:1743" *) _T_2171;
  assign _T_2175 = _T_2141 ^ (* src = "crypto_accelerator.v:1744" *) _T_2167;
  assign _T_2177 = _T_2137 ^ (* src = "crypto_accelerator.v:1745" *) _T_2159;
  assign _T_2179 = _T_2151 ^ (* src = "crypto_accelerator.v:1746" *) _T_2161;
  assign _T_2180 = _T_2147 ^ (* src = "crypto_accelerator.v:1747" *) _T_2173;
  assign _T_2181 = _T_2175 ^ (* src = "crypto_accelerator.v:1748" *) _T_2177;
  assign _T_2184 = _T_2117 ^ (* src = "crypto_accelerator.v:1750" *) _T_2143;
  assign _T_2185 = _T_2155 ^ (* src = "crypto_accelerator.v:1751" *) _T_2157;
  assign _T_2186 = _T_2165 ^ (* src = "crypto_accelerator.v:1752" *) _T_2184;
  assign _T_2188 = _T_2115 ^ (* src = "crypto_accelerator.v:1753" *) _T_2131;
  assign _T_2190 = _T_2153 ^ (* src = "crypto_accelerator.v:1754" *) _T_2169;
  assign _T_2191 = _T_2155 ^ (* src = "crypto_accelerator.v:1755" *) _T_2179;
  assign _T_2194 = _T_2123 ^ (* src = "crypto_accelerator.v:1757" *) _T_2161;
  assign _T_2196 = _T_2188 ^ (* src = "crypto_accelerator.v:1758" *) _T_2194;
  assign _T_2198 = _T_2115 ^ (* src = "crypto_accelerator.v:1759" *) _T_2159;
  assign _T_2199 = _T_2147 ^ (* src = "crypto_accelerator.v:1760" *) _T_2196;
  assign _T_2202 = _T_2167 ^ (* src = "crypto_accelerator.v:1762" *) _T_2190;
  assign _T_2203 = _T_2147 ^ (* src = "crypto_accelerator.v:1763" *) _T_2202;
  assign _T_2205 = _T_2157 ^ (* src = "crypto_accelerator.v:1764" *) _T_2198;
  assign _T_2206 = _T_2147 ^ (* src = "crypto_accelerator.v:1765" *) _T_2205;
  assign _T_2233 = matrix_2_0[1] ^ (* src = "crypto_accelerator.v:1768" *) matrix_2_0[3];
  assign _T_2235 = matrix_2_0[4] ^ (* src = "crypto_accelerator.v:1769" *) matrix_2_0[7];
  assign _T_2237 = matrix_2_0[6] ^ (* src = "crypto_accelerator.v:1770" *) matrix_2_0[5];
  assign _T_2239 = matrix_2_0[0] ^ (* src = "crypto_accelerator.v:1771" *) _T_2237;
  assign _T_2241 = _T_2233 ^ (* src = "crypto_accelerator.v:1772" *) _T_2235;
  assign _T_2243 = matrix_2_0[6] ^ (* src = "crypto_accelerator.v:1773" *) matrix_2_0[2];
  assign _T_2245 = matrix_2_0[7] ^ (* src = "crypto_accelerator.v:1774" *) matrix_2_0[1];
  assign _T_2247 = _T_2233 ^ (* src = "crypto_accelerator.v:1775" *) _T_2243;
  assign _T_2249 = matrix_2_0[1] ^ (* src = "crypto_accelerator.v:1776" *) _T_2239;
  assign _T_2251 = matrix_2_0[4] ^ (* src = "crypto_accelerator.v:1777" *) _T_2239;
  assign _T_2253 = matrix_2_0[0] ^ (* src = "crypto_accelerator.v:1778" *) _T_2241;
  assign _T_2255 = _T_2241 ^ (* src = "crypto_accelerator.v:1779" *) _T_2243;
  assign _T_2257 = matrix_2_0[5] ^ (* src = "crypto_accelerator.v:1780" *) matrix_2_0[2];
  assign _T_2259 = _T_2237 ^ (* src = "crypto_accelerator.v:1781" *) _T_2241;
  assign _T_2261 = matrix_2_0[2] ^ (* src = "crypto_accelerator.v:1782" *) _T_2245;
  assign _T_2263 = matrix_2_0[7] ^ (* src = "crypto_accelerator.v:1783" *) matrix_2_0[2];
  assign _T_2265 = matrix_2_0[0] ^ (* src = "crypto_accelerator.v:1784" *) _T_2247;
  assign _T_2267 = matrix_2_0[1] ^ (* src = "crypto_accelerator.v:1785" *) matrix_2_0[2];
  assign _T_2269 = _T_2235 ^ (* src = "crypto_accelerator.v:1786" *) _T_2267;
  assign _T_2271 = _T_2239 ^ (* src = "crypto_accelerator.v:1787" *) _T_2261;
  assign _T_2273 = _T_2233 ^ (* src = "crypto_accelerator.v:1788" *) _T_2257;
  assign _T_2275 = matrix_2_0[7] ^ (* src = "crypto_accelerator.v:1789" *) _T_2239;
  assign _T_2277 = _T_2273 ^ (* src = "crypto_accelerator.v:1790" *) _T_2241;
  assign _T_2279 = _T_2273 ^ (* src = "crypto_accelerator.v:1791" *) _T_2245;
  assign _T_2281 = _T_2245 ^ (* src = "crypto_accelerator.v:1792" *) _T_2269;
  assign _T_2283 = _T_2263 ^ (* src = "crypto_accelerator.v:1793" *) _T_2259;
  assign _T_2285 = _T_2275 ^ (* src = "crypto_accelerator.v:1794" *) _T_2265;
  assign _T_2291 = _T_2255 ^ (* src = "crypto_accelerator.v:1797" *) _T_2287;
  assign _T_2295 = _T_2293 ^ (* src = "crypto_accelerator.v:1799" *) _T_2287;
  assign _T_2301 = _T_2279 ^ (* src = "crypto_accelerator.v:1802" *) _T_2297;
  assign _T_2305 = _T_2303 ^ (* src = "crypto_accelerator.v:1804" *) _T_2297;
  assign _T_2311 = _T_2309 ^ (* src = "crypto_accelerator.v:1807" *) _T_2307;
  assign _T_2315 = _T_2313 ^ (* src = "crypto_accelerator.v:1809" *) _T_2307;
  assign _T_2317 = _T_2291 ^ (* src = "crypto_accelerator.v:1810" *) _T_2289;
  assign _T_2319 = _T_2295 ^ (* src = "crypto_accelerator.v:1811" *) _T_2283;
  assign _T_2321 = _T_2301 ^ (* src = "crypto_accelerator.v:1812" *) _T_2299;
  assign _T_2323 = _T_2305 ^ (* src = "crypto_accelerator.v:1813" *) _T_2315;
  assign _T_2325 = _T_2317 ^ (* src = "crypto_accelerator.v:1814" *) _T_2311;
  assign _T_2327 = _T_2319 ^ (* src = "crypto_accelerator.v:1815" *) _T_2315;
  assign _T_2329 = _T_2321 ^ (* src = "crypto_accelerator.v:1816" *) _T_2311;
  assign _T_2331 = _T_2323 ^ (* src = "crypto_accelerator.v:1817" *) _T_2285;
  assign _T_2333 = _T_2329 ^ (* src = "crypto_accelerator.v:1818" *) _T_2331;
  assign _T_2337 = _T_2327 ^ (* src = "crypto_accelerator.v:1820" *) _T_2335;
  assign _T_2339 = _T_2325 ^ (* src = "crypto_accelerator.v:1821" *) _T_2327;
  assign _T_2341 = _T_2331 ^ (* src = "crypto_accelerator.v:1822" *) _T_2335;
  assign _T_2351 = _T_2339 ^ (* src = "crypto_accelerator.v:1827" *) _T_2335;
  assign _T_2357 = _T_2333 ^ (* src = "crypto_accelerator.v:1830" *) _T_2335;
  assign _T_2359 = _T_2327 ^ (* src = "crypto_accelerator.v:1831" *) _T_2343;
  assign _T_2361 = _T_2349 ^ (* src = "crypto_accelerator.v:1832" *) _T_2351;
  assign _T_2363 = _T_2331 ^ (* src = "crypto_accelerator.v:1833" *) _T_2345;
  assign _T_2365 = _T_2355 ^ (* src = "crypto_accelerator.v:1834" *) _T_2357;
  assign _T_2367 = _T_2361 ^ (* src = "crypto_accelerator.v:1835" *) _T_2365;
  assign _T_2369 = _T_2359 ^ (* src = "crypto_accelerator.v:1836" *) _T_2363;
  assign _T_2371 = _T_2359 ^ (* src = "crypto_accelerator.v:1837" *) _T_2361;
  assign _T_2373 = _T_2363 ^ (* src = "crypto_accelerator.v:1838" *) _T_2365;
  assign _T_2375 = _T_2369 ^ (* src = "crypto_accelerator.v:1839" *) _T_2367;
  assign _T_2413 = _T_2407 ^ (* src = "crypto_accelerator.v:1858" *) _T_2409;
  assign _T_2415 = _T_2385 ^ (* src = "crypto_accelerator.v:1859" *) _T_2397;
  assign _T_2417 = _T_2391 ^ (* src = "crypto_accelerator.v:1860" *) _T_2413;
  assign _T_2419 = _T_2395 ^ (* src = "crypto_accelerator.v:1861" *) _T_2415;
  assign _T_2421 = _T_2381 ^ (* src = "crypto_accelerator.v:1862" *) _T_2401;
  assign _T_2423 = _T_2377 ^ (* src = "crypto_accelerator.v:1863" *) _T_2383;
  assign _T_2425 = _T_2413 ^ (* src = "crypto_accelerator.v:1864" *) _T_2423;
  assign _T_2427 = _T_2379 ^ (* src = "crypto_accelerator.v:1865" *) _T_2419;
  assign _T_2429 = _T_2377 ^ (* src = "crypto_accelerator.v:1866" *) _T_2389;
  assign _T_2431 = _T_2387 ^ (* src = "crypto_accelerator.v:1867" *) _T_2403;
  assign _T_2433 = _T_2393 ^ (* src = "crypto_accelerator.v:1868" *) _T_2405;
  assign _T_2435 = _T_2381 ^ (* src = "crypto_accelerator.v:1869" *) _T_2427;
  assign _T_2437 = _T_2421 ^ (* src = "crypto_accelerator.v:1870" *) _T_2433;
  assign _T_2439 = _T_2399 ^ (* src = "crypto_accelerator.v:1871" *) _T_2415;
  assign _T_2441 = _T_2383 ^ (* src = "crypto_accelerator.v:1872" *) _T_2389;
  assign _T_2443 = _T_2419 ^ (* src = "crypto_accelerator.v:1873" *) _T_2441;
  assign _T_2445 = _T_2411 ^ (* src = "crypto_accelerator.v:1874" *) _T_2437;
  assign _T_2447 = _T_2407 ^ (* src = "crypto_accelerator.v:1875" *) _T_2429;
  assign _T_2449 = _T_2421 ^ (* src = "crypto_accelerator.v:1876" *) _T_2431;
  assign _T_2450 = _T_2417 ^ (* src = "crypto_accelerator.v:1877" *) _T_2443;
  assign _T_2451 = _T_2445 ^ (* src = "crypto_accelerator.v:1878" *) _T_2447;
  assign _T_2454 = _T_2387 ^ (* src = "crypto_accelerator.v:1880" *) _T_2413;
  assign _T_2455 = _T_2425 ^ (* src = "crypto_accelerator.v:1881" *) _T_2427;
  assign _T_2456 = _T_2435 ^ (* src = "crypto_accelerator.v:1882" *) _T_2454;
  assign _T_2458 = _T_2385 ^ (* src = "crypto_accelerator.v:1883" *) _T_2401;
  assign _T_2460 = _T_2423 ^ (* src = "crypto_accelerator.v:1884" *) _T_2439;
  assign _T_2461 = _T_2425 ^ (* src = "crypto_accelerator.v:1885" *) _T_2449;
  assign _T_2464 = _T_2393 ^ (* src = "crypto_accelerator.v:1887" *) _T_2431;
  assign _T_2466 = _T_2458 ^ (* src = "crypto_accelerator.v:1888" *) _T_2464;
  assign _T_2468 = _T_2385 ^ (* src = "crypto_accelerator.v:1889" *) _T_2429;
  assign _T_2469 = _T_2417 ^ (* src = "crypto_accelerator.v:1890" *) _T_2466;
  assign _T_2472 = _T_2437 ^ (* src = "crypto_accelerator.v:1892" *) _T_2460;
  assign _T_2473 = _T_2417 ^ (* src = "crypto_accelerator.v:1893" *) _T_2472;
  assign _T_2475 = _T_2427 ^ (* src = "crypto_accelerator.v:1894" *) _T_2468;
  assign _T_2476 = _T_2417 ^ (* src = "crypto_accelerator.v:1895" *) _T_2475;
  assign _T_2502 = matrix_2_1[1] ^ (* src = "crypto_accelerator.v:1898" *) matrix_2_1[3];
  assign _T_2504 = matrix_2_1[4] ^ (* src = "crypto_accelerator.v:1899" *) matrix_2_1[7];
  assign _T_2506 = matrix_2_1[6] ^ (* src = "crypto_accelerator.v:1900" *) matrix_2_1[5];
  assign _T_2508 = matrix_2_1[0] ^ (* src = "crypto_accelerator.v:1901" *) _T_2506;
  assign _T_2510 = _T_2502 ^ (* src = "crypto_accelerator.v:1902" *) _T_2504;
  assign _T_2512 = matrix_2_1[6] ^ (* src = "crypto_accelerator.v:1903" *) matrix_2_1[2];
  assign _T_2514 = matrix_2_1[7] ^ (* src = "crypto_accelerator.v:1904" *) matrix_2_1[1];
  assign _T_2516 = _T_2502 ^ (* src = "crypto_accelerator.v:1905" *) _T_2512;
  assign _T_2518 = matrix_2_1[1] ^ (* src = "crypto_accelerator.v:1906" *) _T_2508;
  assign _T_2520 = matrix_2_1[4] ^ (* src = "crypto_accelerator.v:1907" *) _T_2508;
  assign _T_2522 = matrix_2_1[0] ^ (* src = "crypto_accelerator.v:1908" *) _T_2510;
  assign _T_2524 = _T_2510 ^ (* src = "crypto_accelerator.v:1909" *) _T_2512;
  assign _T_2526 = matrix_2_1[5] ^ (* src = "crypto_accelerator.v:1910" *) matrix_2_1[2];
  assign _T_2528 = _T_2506 ^ (* src = "crypto_accelerator.v:1911" *) _T_2510;
  assign _T_2530 = matrix_2_1[2] ^ (* src = "crypto_accelerator.v:1912" *) _T_2514;
  assign _T_2532 = matrix_2_1[7] ^ (* src = "crypto_accelerator.v:1913" *) matrix_2_1[2];
  assign _T_2534 = matrix_2_1[0] ^ (* src = "crypto_accelerator.v:1914" *) _T_2516;
  assign _T_2536 = matrix_2_1[1] ^ (* src = "crypto_accelerator.v:1915" *) matrix_2_1[2];
  assign _T_2538 = _T_2504 ^ (* src = "crypto_accelerator.v:1916" *) _T_2536;
  assign _T_2540 = _T_2508 ^ (* src = "crypto_accelerator.v:1917" *) _T_2530;
  assign _T_2542 = _T_2502 ^ (* src = "crypto_accelerator.v:1918" *) _T_2526;
  assign _T_2544 = matrix_2_1[7] ^ (* src = "crypto_accelerator.v:1919" *) _T_2508;
  assign _T_2546 = _T_2542 ^ (* src = "crypto_accelerator.v:1920" *) _T_2510;
  assign _T_2548 = _T_2542 ^ (* src = "crypto_accelerator.v:1921" *) _T_2514;
  assign _T_2550 = _T_2514 ^ (* src = "crypto_accelerator.v:1922" *) _T_2538;
  assign _T_2552 = _T_2532 ^ (* src = "crypto_accelerator.v:1923" *) _T_2528;
  assign _T_2554 = _T_2544 ^ (* src = "crypto_accelerator.v:1924" *) _T_2534;
  assign _T_2560 = _T_2524 ^ (* src = "crypto_accelerator.v:1927" *) _T_2556;
  assign _T_2564 = _T_2562 ^ (* src = "crypto_accelerator.v:1929" *) _T_2556;
  assign _T_2570 = _T_2548 ^ (* src = "crypto_accelerator.v:1932" *) _T_2566;
  assign _T_2574 = _T_2572 ^ (* src = "crypto_accelerator.v:1934" *) _T_2566;
  assign _T_2580 = _T_2578 ^ (* src = "crypto_accelerator.v:1937" *) _T_2576;
  assign _T_2584 = _T_2582 ^ (* src = "crypto_accelerator.v:1939" *) _T_2576;
  assign _T_2586 = _T_2560 ^ (* src = "crypto_accelerator.v:1940" *) _T_2558;
  assign _T_2588 = _T_2564 ^ (* src = "crypto_accelerator.v:1941" *) _T_2552;
  assign _T_2590 = _T_2570 ^ (* src = "crypto_accelerator.v:1942" *) _T_2568;
  assign _T_2592 = _T_2574 ^ (* src = "crypto_accelerator.v:1943" *) _T_2584;
  assign _T_2594 = _T_2586 ^ (* src = "crypto_accelerator.v:1944" *) _T_2580;
  assign _T_2596 = _T_2588 ^ (* src = "crypto_accelerator.v:1945" *) _T_2584;
  assign _T_2598 = _T_2590 ^ (* src = "crypto_accelerator.v:1946" *) _T_2580;
  assign _T_2600 = _T_2592 ^ (* src = "crypto_accelerator.v:1947" *) _T_2554;
  assign _T_2602 = _T_2598 ^ (* src = "crypto_accelerator.v:1948" *) _T_2600;
  assign _T_2606 = _T_2596 ^ (* src = "crypto_accelerator.v:1950" *) _T_2604;
  assign _T_2608 = _T_2594 ^ (* src = "crypto_accelerator.v:1951" *) _T_2596;
  assign _T_2610 = _T_2600 ^ (* src = "crypto_accelerator.v:1952" *) _T_2604;
  assign _T_2620 = _T_2608 ^ (* src = "crypto_accelerator.v:1957" *) _T_2604;
  assign _T_2626 = _T_2602 ^ (* src = "crypto_accelerator.v:1960" *) _T_2604;
  assign _T_2628 = _T_2596 ^ (* src = "crypto_accelerator.v:1961" *) _T_2612;
  assign _T_2630 = _T_2618 ^ (* src = "crypto_accelerator.v:1962" *) _T_2620;
  assign _T_2632 = _T_2600 ^ (* src = "crypto_accelerator.v:1963" *) _T_2614;
  assign _T_2634 = _T_2624 ^ (* src = "crypto_accelerator.v:1964" *) _T_2626;
  assign _T_2636 = _T_2630 ^ (* src = "crypto_accelerator.v:1965" *) _T_2634;
  assign _T_2638 = _T_2628 ^ (* src = "crypto_accelerator.v:1966" *) _T_2632;
  assign _T_2640 = _T_2628 ^ (* src = "crypto_accelerator.v:1967" *) _T_2630;
  assign _T_2642 = _T_2632 ^ (* src = "crypto_accelerator.v:1968" *) _T_2634;
  assign _T_2644 = _T_2638 ^ (* src = "crypto_accelerator.v:1969" *) _T_2636;
  assign _T_2682 = _T_2676 ^ (* src = "crypto_accelerator.v:1988" *) _T_2678;
  assign _T_2684 = _T_2654 ^ (* src = "crypto_accelerator.v:1989" *) _T_2666;
  assign _T_2686 = _T_2660 ^ (* src = "crypto_accelerator.v:1990" *) _T_2682;
  assign _T_2688 = _T_2664 ^ (* src = "crypto_accelerator.v:1991" *) _T_2684;
  assign _T_2690 = _T_2650 ^ (* src = "crypto_accelerator.v:1992" *) _T_2670;
  assign _T_2692 = _T_2646 ^ (* src = "crypto_accelerator.v:1993" *) _T_2652;
  assign _T_2694 = _T_2682 ^ (* src = "crypto_accelerator.v:1994" *) _T_2692;
  assign _T_2696 = _T_2648 ^ (* src = "crypto_accelerator.v:1995" *) _T_2688;
  assign _T_2698 = _T_2646 ^ (* src = "crypto_accelerator.v:1996" *) _T_2658;
  assign _T_2700 = _T_2656 ^ (* src = "crypto_accelerator.v:1997" *) _T_2672;
  assign _T_2702 = _T_2662 ^ (* src = "crypto_accelerator.v:1998" *) _T_2674;
  assign _T_2704 = _T_2650 ^ (* src = "crypto_accelerator.v:1999" *) _T_2696;
  assign _T_2706 = _T_2690 ^ (* src = "crypto_accelerator.v:2000" *) _T_2702;
  assign _T_2708 = _T_2668 ^ (* src = "crypto_accelerator.v:2001" *) _T_2684;
  assign _T_2710 = _T_2652 ^ (* src = "crypto_accelerator.v:2002" *) _T_2658;
  assign _T_2712 = _T_2688 ^ (* src = "crypto_accelerator.v:2003" *) _T_2710;
  assign _T_2714 = _T_2680 ^ (* src = "crypto_accelerator.v:2004" *) _T_2706;
  assign _T_2716 = _T_2676 ^ (* src = "crypto_accelerator.v:2005" *) _T_2698;
  assign _T_2718 = _T_2690 ^ (* src = "crypto_accelerator.v:2006" *) _T_2700;
  assign _T_2719 = _T_2686 ^ (* src = "crypto_accelerator.v:2007" *) _T_2712;
  assign _T_2720 = _T_2714 ^ (* src = "crypto_accelerator.v:2008" *) _T_2716;
  assign _T_2723 = _T_2656 ^ (* src = "crypto_accelerator.v:2010" *) _T_2682;
  assign _T_2724 = _T_2694 ^ (* src = "crypto_accelerator.v:2011" *) _T_2696;
  assign _T_2725 = _T_2704 ^ (* src = "crypto_accelerator.v:2012" *) _T_2723;
  assign _T_2727 = _T_2654 ^ (* src = "crypto_accelerator.v:2013" *) _T_2670;
  assign _T_2729 = _T_2692 ^ (* src = "crypto_accelerator.v:2014" *) _T_2708;
  assign _T_2730 = _T_2694 ^ (* src = "crypto_accelerator.v:2015" *) _T_2718;
  assign _T_2733 = _T_2662 ^ (* src = "crypto_accelerator.v:2017" *) _T_2700;
  assign _T_2735 = _T_2727 ^ (* src = "crypto_accelerator.v:2018" *) _T_2733;
  assign _T_2737 = _T_2654 ^ (* src = "crypto_accelerator.v:2019" *) _T_2698;
  assign _T_2738 = _T_2686 ^ (* src = "crypto_accelerator.v:2020" *) _T_2735;
  assign _T_2741 = _T_2706 ^ (* src = "crypto_accelerator.v:2022" *) _T_2729;
  assign _T_2742 = _T_2686 ^ (* src = "crypto_accelerator.v:2023" *) _T_2741;
  assign _T_2744 = _T_2696 ^ (* src = "crypto_accelerator.v:2024" *) _T_2737;
  assign _T_2745 = _T_2686 ^ (* src = "crypto_accelerator.v:2025" *) _T_2744;
  assign _T_2771 = matrix_2_2[1] ^ (* src = "crypto_accelerator.v:2028" *) matrix_2_2[3];
  assign _T_2773 = matrix_2_2[4] ^ (* src = "crypto_accelerator.v:2029" *) matrix_2_2[7];
  assign _T_2775 = matrix_2_2[6] ^ (* src = "crypto_accelerator.v:2030" *) matrix_2_2[5];
  assign _T_2777 = matrix_2_2[0] ^ (* src = "crypto_accelerator.v:2031" *) _T_2775;
  assign _T_2779 = _T_2771 ^ (* src = "crypto_accelerator.v:2032" *) _T_2773;
  assign _T_2781 = matrix_2_2[6] ^ (* src = "crypto_accelerator.v:2033" *) matrix_2_2[2];
  assign _T_2783 = matrix_2_2[7] ^ (* src = "crypto_accelerator.v:2034" *) matrix_2_2[1];
  assign _T_2785 = _T_2771 ^ (* src = "crypto_accelerator.v:2035" *) _T_2781;
  assign _T_2787 = matrix_2_2[1] ^ (* src = "crypto_accelerator.v:2036" *) _T_2777;
  assign _T_2789 = matrix_2_2[4] ^ (* src = "crypto_accelerator.v:2037" *) _T_2777;
  assign _T_2791 = matrix_2_2[0] ^ (* src = "crypto_accelerator.v:2038" *) _T_2779;
  assign _T_2793 = _T_2779 ^ (* src = "crypto_accelerator.v:2039" *) _T_2781;
  assign _T_2795 = matrix_2_2[5] ^ (* src = "crypto_accelerator.v:2040" *) matrix_2_2[2];
  assign _T_2797 = _T_2775 ^ (* src = "crypto_accelerator.v:2041" *) _T_2779;
  assign _T_2799 = matrix_2_2[2] ^ (* src = "crypto_accelerator.v:2042" *) _T_2783;
  assign _T_2801 = matrix_2_2[7] ^ (* src = "crypto_accelerator.v:2043" *) matrix_2_2[2];
  assign _T_2803 = matrix_2_2[0] ^ (* src = "crypto_accelerator.v:2044" *) _T_2785;
  assign _T_2805 = matrix_2_2[1] ^ (* src = "crypto_accelerator.v:2045" *) matrix_2_2[2];
  assign _T_2807 = _T_2773 ^ (* src = "crypto_accelerator.v:2046" *) _T_2805;
  assign _T_2809 = _T_2777 ^ (* src = "crypto_accelerator.v:2047" *) _T_2799;
  assign _T_2811 = _T_2771 ^ (* src = "crypto_accelerator.v:2048" *) _T_2795;
  assign _T_2813 = matrix_2_2[7] ^ (* src = "crypto_accelerator.v:2049" *) _T_2777;
  assign _T_2815 = _T_2811 ^ (* src = "crypto_accelerator.v:2050" *) _T_2779;
  assign _T_2817 = _T_2811 ^ (* src = "crypto_accelerator.v:2051" *) _T_2783;
  assign _T_2819 = _T_2783 ^ (* src = "crypto_accelerator.v:2052" *) _T_2807;
  assign _T_2821 = _T_2801 ^ (* src = "crypto_accelerator.v:2053" *) _T_2797;
  assign _T_2823 = _T_2813 ^ (* src = "crypto_accelerator.v:2054" *) _T_2803;
  assign _T_2829 = _T_2793 ^ (* src = "crypto_accelerator.v:2057" *) _T_2825;
  assign _T_2833 = _T_2831 ^ (* src = "crypto_accelerator.v:2059" *) _T_2825;
  assign _T_2839 = _T_2817 ^ (* src = "crypto_accelerator.v:2062" *) _T_2835;
  assign _T_2843 = _T_2841 ^ (* src = "crypto_accelerator.v:2064" *) _T_2835;
  assign _T_2849 = _T_2847 ^ (* src = "crypto_accelerator.v:2067" *) _T_2845;
  assign _T_2853 = _T_2851 ^ (* src = "crypto_accelerator.v:2069" *) _T_2845;
  assign _T_2855 = _T_2829 ^ (* src = "crypto_accelerator.v:2070" *) _T_2827;
  assign _T_2857 = _T_2833 ^ (* src = "crypto_accelerator.v:2071" *) _T_2821;
  assign _T_2859 = _T_2839 ^ (* src = "crypto_accelerator.v:2072" *) _T_2837;
  assign _T_2861 = _T_2843 ^ (* src = "crypto_accelerator.v:2073" *) _T_2853;
  assign _T_2863 = _T_2855 ^ (* src = "crypto_accelerator.v:2074" *) _T_2849;
  assign _T_2865 = _T_2857 ^ (* src = "crypto_accelerator.v:2075" *) _T_2853;
  assign _T_2867 = _T_2859 ^ (* src = "crypto_accelerator.v:2076" *) _T_2849;
  assign _T_2869 = _T_2861 ^ (* src = "crypto_accelerator.v:2077" *) _T_2823;
  assign _T_2871 = _T_2867 ^ (* src = "crypto_accelerator.v:2078" *) _T_2869;
  assign _T_2875 = _T_2865 ^ (* src = "crypto_accelerator.v:2080" *) _T_2873;
  assign _T_2877 = _T_2863 ^ (* src = "crypto_accelerator.v:2081" *) _T_2865;
  assign _T_2879 = _T_2869 ^ (* src = "crypto_accelerator.v:2082" *) _T_2873;
  assign _T_2889 = _T_2877 ^ (* src = "crypto_accelerator.v:2087" *) _T_2873;
  assign _T_2895 = _T_2871 ^ (* src = "crypto_accelerator.v:2090" *) _T_2873;
  assign _T_2897 = _T_2865 ^ (* src = "crypto_accelerator.v:2091" *) _T_2881;
  assign _T_2899 = _T_2887 ^ (* src = "crypto_accelerator.v:2092" *) _T_2889;
  assign _T_2901 = _T_2869 ^ (* src = "crypto_accelerator.v:2093" *) _T_2883;
  assign _T_2903 = _T_2893 ^ (* src = "crypto_accelerator.v:2094" *) _T_2895;
  assign _T_2905 = _T_2899 ^ (* src = "crypto_accelerator.v:2095" *) _T_2903;
  assign _T_2907 = _T_2897 ^ (* src = "crypto_accelerator.v:2096" *) _T_2901;
  assign _T_2909 = _T_2897 ^ (* src = "crypto_accelerator.v:2097" *) _T_2899;
  assign _T_2911 = _T_2901 ^ (* src = "crypto_accelerator.v:2098" *) _T_2903;
  assign _T_2913 = _T_2907 ^ (* src = "crypto_accelerator.v:2099" *) _T_2905;
  assign _T_2951 = _T_2945 ^ (* src = "crypto_accelerator.v:2118" *) _T_2947;
  assign _T_2953 = _T_2923 ^ (* src = "crypto_accelerator.v:2119" *) _T_2935;
  assign _T_2955 = _T_2929 ^ (* src = "crypto_accelerator.v:2120" *) _T_2951;
  assign _T_2957 = _T_2933 ^ (* src = "crypto_accelerator.v:2121" *) _T_2953;
  assign _T_2959 = _T_2919 ^ (* src = "crypto_accelerator.v:2122" *) _T_2939;
  assign _T_2961 = _T_2915 ^ (* src = "crypto_accelerator.v:2123" *) _T_2921;
  assign _T_2963 = _T_2951 ^ (* src = "crypto_accelerator.v:2124" *) _T_2961;
  assign _T_2965 = _T_2917 ^ (* src = "crypto_accelerator.v:2125" *) _T_2957;
  assign _T_2967 = _T_2915 ^ (* src = "crypto_accelerator.v:2126" *) _T_2927;
  assign _T_2969 = _T_2925 ^ (* src = "crypto_accelerator.v:2127" *) _T_2941;
  assign _T_2971 = _T_2931 ^ (* src = "crypto_accelerator.v:2128" *) _T_2943;
  assign _T_2973 = _T_2919 ^ (* src = "crypto_accelerator.v:2129" *) _T_2965;
  assign _T_2975 = _T_2959 ^ (* src = "crypto_accelerator.v:2130" *) _T_2971;
  assign _T_2977 = _T_2937 ^ (* src = "crypto_accelerator.v:2131" *) _T_2953;
  assign _T_2979 = _T_2921 ^ (* src = "crypto_accelerator.v:2132" *) _T_2927;
  assign _T_2981 = _T_2957 ^ (* src = "crypto_accelerator.v:2133" *) _T_2979;
  assign _T_2983 = _T_2949 ^ (* src = "crypto_accelerator.v:2134" *) _T_2975;
  assign _T_2985 = _T_2945 ^ (* src = "crypto_accelerator.v:2135" *) _T_2967;
  assign _T_2987 = _T_2959 ^ (* src = "crypto_accelerator.v:2136" *) _T_2969;
  assign _T_2988 = _T_2955 ^ (* src = "crypto_accelerator.v:2137" *) _T_2981;
  assign _T_2989 = _T_2983 ^ (* src = "crypto_accelerator.v:2138" *) _T_2985;
  assign _T_2992 = _T_2925 ^ (* src = "crypto_accelerator.v:2140" *) _T_2951;
  assign _T_2993 = _T_2963 ^ (* src = "crypto_accelerator.v:2141" *) _T_2965;
  assign _T_2994 = _T_2973 ^ (* src = "crypto_accelerator.v:2142" *) _T_2992;
  assign _T_2996 = _T_2923 ^ (* src = "crypto_accelerator.v:2143" *) _T_2939;
  assign _T_2998 = _T_2961 ^ (* src = "crypto_accelerator.v:2144" *) _T_2977;
  assign _T_2999 = _T_2963 ^ (* src = "crypto_accelerator.v:2145" *) _T_2987;
  assign _T_3002 = _T_2931 ^ (* src = "crypto_accelerator.v:2147" *) _T_2969;
  assign _T_3004 = _T_2996 ^ (* src = "crypto_accelerator.v:2148" *) _T_3002;
  assign _T_3006 = _T_2923 ^ (* src = "crypto_accelerator.v:2149" *) _T_2967;
  assign _T_3007 = _T_2955 ^ (* src = "crypto_accelerator.v:2150" *) _T_3004;
  assign _T_3010 = _T_2975 ^ (* src = "crypto_accelerator.v:2152" *) _T_2998;
  assign _T_3011 = _T_2955 ^ (* src = "crypto_accelerator.v:2153" *) _T_3010;
  assign _T_3013 = _T_2965 ^ (* src = "crypto_accelerator.v:2154" *) _T_3006;
  assign _T_3014 = _T_2955 ^ (* src = "crypto_accelerator.v:2155" *) _T_3013;
  assign _T_3040 = matrix_2_3[1] ^ (* src = "crypto_accelerator.v:2158" *) matrix_2_3[3];
  assign _T_3042 = matrix_2_3[4] ^ (* src = "crypto_accelerator.v:2159" *) matrix_2_3[7];
  assign _T_3044 = matrix_2_3[6] ^ (* src = "crypto_accelerator.v:2160" *) matrix_2_3[5];
  assign _T_3046 = matrix_2_3[0] ^ (* src = "crypto_accelerator.v:2161" *) _T_3044;
  assign _T_3048 = _T_3040 ^ (* src = "crypto_accelerator.v:2162" *) _T_3042;
  assign _T_3050 = matrix_2_3[6] ^ (* src = "crypto_accelerator.v:2163" *) matrix_2_3[2];
  assign _T_3052 = matrix_2_3[7] ^ (* src = "crypto_accelerator.v:2164" *) matrix_2_3[1];
  assign _T_3054 = _T_3040 ^ (* src = "crypto_accelerator.v:2165" *) _T_3050;
  assign _T_3056 = matrix_2_3[1] ^ (* src = "crypto_accelerator.v:2166" *) _T_3046;
  assign _T_3058 = matrix_2_3[4] ^ (* src = "crypto_accelerator.v:2167" *) _T_3046;
  assign _T_3060 = matrix_2_3[0] ^ (* src = "crypto_accelerator.v:2168" *) _T_3048;
  assign _T_3062 = _T_3048 ^ (* src = "crypto_accelerator.v:2169" *) _T_3050;
  assign _T_3064 = matrix_2_3[5] ^ (* src = "crypto_accelerator.v:2170" *) matrix_2_3[2];
  assign _T_3066 = _T_3044 ^ (* src = "crypto_accelerator.v:2171" *) _T_3048;
  assign _T_3068 = matrix_2_3[2] ^ (* src = "crypto_accelerator.v:2172" *) _T_3052;
  assign _T_3070 = matrix_2_3[7] ^ (* src = "crypto_accelerator.v:2173" *) matrix_2_3[2];
  assign _T_3072 = matrix_2_3[0] ^ (* src = "crypto_accelerator.v:2174" *) _T_3054;
  assign _T_3074 = matrix_2_3[1] ^ (* src = "crypto_accelerator.v:2175" *) matrix_2_3[2];
  assign _T_3076 = _T_3042 ^ (* src = "crypto_accelerator.v:2176" *) _T_3074;
  assign _T_3078 = _T_3046 ^ (* src = "crypto_accelerator.v:2177" *) _T_3068;
  assign _T_3080 = _T_3040 ^ (* src = "crypto_accelerator.v:2178" *) _T_3064;
  assign _T_3082 = matrix_2_3[7] ^ (* src = "crypto_accelerator.v:2179" *) _T_3046;
  assign _T_3084 = _T_3080 ^ (* src = "crypto_accelerator.v:2180" *) _T_3048;
  assign _T_3086 = _T_3080 ^ (* src = "crypto_accelerator.v:2181" *) _T_3052;
  assign _T_3088 = _T_3052 ^ (* src = "crypto_accelerator.v:2182" *) _T_3076;
  assign _T_3090 = _T_3070 ^ (* src = "crypto_accelerator.v:2183" *) _T_3066;
  assign _T_3092 = _T_3082 ^ (* src = "crypto_accelerator.v:2184" *) _T_3072;
  assign _T_3098 = _T_3062 ^ (* src = "crypto_accelerator.v:2187" *) _T_3094;
  assign _T_3102 = _T_3100 ^ (* src = "crypto_accelerator.v:2189" *) _T_3094;
  assign _T_3108 = _T_3086 ^ (* src = "crypto_accelerator.v:2192" *) _T_3104;
  assign _T_3112 = _T_3110 ^ (* src = "crypto_accelerator.v:2194" *) _T_3104;
  assign _T_3118 = _T_3116 ^ (* src = "crypto_accelerator.v:2197" *) _T_3114;
  assign _T_3122 = _T_3120 ^ (* src = "crypto_accelerator.v:2199" *) _T_3114;
  assign _T_3124 = _T_3098 ^ (* src = "crypto_accelerator.v:2200" *) _T_3096;
  assign _T_3126 = _T_3102 ^ (* src = "crypto_accelerator.v:2201" *) _T_3090;
  assign _T_3128 = _T_3108 ^ (* src = "crypto_accelerator.v:2202" *) _T_3106;
  assign _T_3130 = _T_3112 ^ (* src = "crypto_accelerator.v:2203" *) _T_3122;
  assign _T_3132 = _T_3124 ^ (* src = "crypto_accelerator.v:2204" *) _T_3118;
  assign _T_3134 = _T_3126 ^ (* src = "crypto_accelerator.v:2205" *) _T_3122;
  assign _T_3136 = _T_3128 ^ (* src = "crypto_accelerator.v:2206" *) _T_3118;
  assign _T_3138 = _T_3130 ^ (* src = "crypto_accelerator.v:2207" *) _T_3092;
  assign _T_3140 = _T_3136 ^ (* src = "crypto_accelerator.v:2208" *) _T_3138;
  assign _T_3144 = _T_3134 ^ (* src = "crypto_accelerator.v:2210" *) _T_3142;
  assign _T_3146 = _T_3132 ^ (* src = "crypto_accelerator.v:2211" *) _T_3134;
  assign _T_3148 = _T_3138 ^ (* src = "crypto_accelerator.v:2212" *) _T_3142;
  assign _T_3158 = _T_3146 ^ (* src = "crypto_accelerator.v:2217" *) _T_3142;
  assign _T_3164 = _T_3140 ^ (* src = "crypto_accelerator.v:2220" *) _T_3142;
  assign _T_3166 = _T_3134 ^ (* src = "crypto_accelerator.v:2221" *) _T_3150;
  assign _T_3168 = _T_3156 ^ (* src = "crypto_accelerator.v:2222" *) _T_3158;
  assign _T_3170 = _T_3138 ^ (* src = "crypto_accelerator.v:2223" *) _T_3152;
  assign _T_3172 = _T_3162 ^ (* src = "crypto_accelerator.v:2224" *) _T_3164;
  assign _T_3174 = _T_3168 ^ (* src = "crypto_accelerator.v:2225" *) _T_3172;
  assign _T_3176 = _T_3166 ^ (* src = "crypto_accelerator.v:2226" *) _T_3170;
  assign _T_3178 = _T_3166 ^ (* src = "crypto_accelerator.v:2227" *) _T_3168;
  assign _T_3180 = _T_3170 ^ (* src = "crypto_accelerator.v:2228" *) _T_3172;
  assign _T_3182 = _T_3176 ^ (* src = "crypto_accelerator.v:2229" *) _T_3174;
  assign _T_3220 = _T_3214 ^ (* src = "crypto_accelerator.v:2248" *) _T_3216;
  assign _T_3222 = _T_3192 ^ (* src = "crypto_accelerator.v:2249" *) _T_3204;
  assign _T_3224 = _T_3198 ^ (* src = "crypto_accelerator.v:2250" *) _T_3220;
  assign _T_3226 = _T_3202 ^ (* src = "crypto_accelerator.v:2251" *) _T_3222;
  assign _T_3228 = _T_3188 ^ (* src = "crypto_accelerator.v:2252" *) _T_3208;
  assign _T_3230 = _T_3184 ^ (* src = "crypto_accelerator.v:2253" *) _T_3190;
  assign _T_3232 = _T_3220 ^ (* src = "crypto_accelerator.v:2254" *) _T_3230;
  assign _T_3234 = _T_3186 ^ (* src = "crypto_accelerator.v:2255" *) _T_3226;
  assign _T_3236 = _T_3184 ^ (* src = "crypto_accelerator.v:2256" *) _T_3196;
  assign _T_3238 = _T_3194 ^ (* src = "crypto_accelerator.v:2257" *) _T_3210;
  assign _T_3240 = _T_3200 ^ (* src = "crypto_accelerator.v:2258" *) _T_3212;
  assign _T_3242 = _T_3188 ^ (* src = "crypto_accelerator.v:2259" *) _T_3234;
  assign _T_3244 = _T_3228 ^ (* src = "crypto_accelerator.v:2260" *) _T_3240;
  assign _T_3246 = _T_3206 ^ (* src = "crypto_accelerator.v:2261" *) _T_3222;
  assign _T_3248 = _T_3190 ^ (* src = "crypto_accelerator.v:2262" *) _T_3196;
  assign _T_3250 = _T_3226 ^ (* src = "crypto_accelerator.v:2263" *) _T_3248;
  assign _T_3252 = _T_3218 ^ (* src = "crypto_accelerator.v:2264" *) _T_3244;
  assign _T_3254 = _T_3214 ^ (* src = "crypto_accelerator.v:2265" *) _T_3236;
  assign _T_3256 = _T_3228 ^ (* src = "crypto_accelerator.v:2266" *) _T_3238;
  assign _T_3257 = _T_3224 ^ (* src = "crypto_accelerator.v:2267" *) _T_3250;
  assign _T_3258 = _T_3252 ^ (* src = "crypto_accelerator.v:2268" *) _T_3254;
  assign _T_3261 = _T_3194 ^ (* src = "crypto_accelerator.v:2270" *) _T_3220;
  assign _T_3262 = _T_3232 ^ (* src = "crypto_accelerator.v:2271" *) _T_3234;
  assign _T_3263 = _T_3242 ^ (* src = "crypto_accelerator.v:2272" *) _T_3261;
  assign _T_3265 = _T_3192 ^ (* src = "crypto_accelerator.v:2273" *) _T_3208;
  assign _T_3267 = _T_3230 ^ (* src = "crypto_accelerator.v:2274" *) _T_3246;
  assign _T_3268 = _T_3232 ^ (* src = "crypto_accelerator.v:2275" *) _T_3256;
  assign _T_3271 = _T_3200 ^ (* src = "crypto_accelerator.v:2277" *) _T_3238;
  assign _T_3273 = _T_3265 ^ (* src = "crypto_accelerator.v:2278" *) _T_3271;
  assign _T_3275 = _T_3192 ^ (* src = "crypto_accelerator.v:2279" *) _T_3236;
  assign _T_3276 = _T_3224 ^ (* src = "crypto_accelerator.v:2280" *) _T_3273;
  assign _T_3279 = _T_3244 ^ (* src = "crypto_accelerator.v:2282" *) _T_3267;
  assign _T_3280 = _T_3224 ^ (* src = "crypto_accelerator.v:2283" *) _T_3279;
  assign _T_3282 = _T_3234 ^ (* src = "crypto_accelerator.v:2284" *) _T_3275;
  assign _T_3283 = _T_3224 ^ (* src = "crypto_accelerator.v:2285" *) _T_3282;
  assign _T_3310 = matrix_3_0[1] ^ (* src = "crypto_accelerator.v:2288" *) matrix_3_0[3];
  assign _T_3312 = matrix_3_0[4] ^ (* src = "crypto_accelerator.v:2289" *) matrix_3_0[7];
  assign _T_3314 = matrix_3_0[6] ^ (* src = "crypto_accelerator.v:2290" *) matrix_3_0[5];
  assign _T_3316 = matrix_3_0[0] ^ (* src = "crypto_accelerator.v:2291" *) _T_3314;
  assign _T_3318 = _T_3310 ^ (* src = "crypto_accelerator.v:2292" *) _T_3312;
  assign _T_3320 = matrix_3_0[6] ^ (* src = "crypto_accelerator.v:2293" *) matrix_3_0[2];
  assign _T_3322 = matrix_3_0[7] ^ (* src = "crypto_accelerator.v:2294" *) matrix_3_0[1];
  assign _T_3324 = _T_3310 ^ (* src = "crypto_accelerator.v:2295" *) _T_3320;
  assign _T_3326 = matrix_3_0[1] ^ (* src = "crypto_accelerator.v:2296" *) _T_3316;
  assign _T_3328 = matrix_3_0[4] ^ (* src = "crypto_accelerator.v:2297" *) _T_3316;
  assign _T_3330 = matrix_3_0[0] ^ (* src = "crypto_accelerator.v:2298" *) _T_3318;
  assign _T_3332 = _T_3318 ^ (* src = "crypto_accelerator.v:2299" *) _T_3320;
  assign _T_3334 = matrix_3_0[5] ^ (* src = "crypto_accelerator.v:2300" *) matrix_3_0[2];
  assign _T_3336 = _T_3314 ^ (* src = "crypto_accelerator.v:2301" *) _T_3318;
  assign _T_3338 = matrix_3_0[2] ^ (* src = "crypto_accelerator.v:2302" *) _T_3322;
  assign _T_3340 = matrix_3_0[7] ^ (* src = "crypto_accelerator.v:2303" *) matrix_3_0[2];
  assign _T_3342 = matrix_3_0[0] ^ (* src = "crypto_accelerator.v:2304" *) _T_3324;
  assign _T_3344 = matrix_3_0[1] ^ (* src = "crypto_accelerator.v:2305" *) matrix_3_0[2];
  assign _T_3346 = _T_3312 ^ (* src = "crypto_accelerator.v:2306" *) _T_3344;
  assign _T_3348 = _T_3316 ^ (* src = "crypto_accelerator.v:2307" *) _T_3338;
  assign _T_3350 = _T_3310 ^ (* src = "crypto_accelerator.v:2308" *) _T_3334;
  assign _T_3352 = matrix_3_0[7] ^ (* src = "crypto_accelerator.v:2309" *) _T_3316;
  assign _T_3354 = _T_3350 ^ (* src = "crypto_accelerator.v:2310" *) _T_3318;
  assign _T_3356 = _T_3350 ^ (* src = "crypto_accelerator.v:2311" *) _T_3322;
  assign _T_3358 = _T_3322 ^ (* src = "crypto_accelerator.v:2312" *) _T_3346;
  assign _T_3360 = _T_3340 ^ (* src = "crypto_accelerator.v:2313" *) _T_3336;
  assign _T_3362 = _T_3352 ^ (* src = "crypto_accelerator.v:2314" *) _T_3342;
  assign _T_3368 = _T_3332 ^ (* src = "crypto_accelerator.v:2317" *) _T_3364;
  assign _T_3372 = _T_3370 ^ (* src = "crypto_accelerator.v:2319" *) _T_3364;
  assign _T_3378 = _T_3356 ^ (* src = "crypto_accelerator.v:2322" *) _T_3374;
  assign _T_3382 = _T_3380 ^ (* src = "crypto_accelerator.v:2324" *) _T_3374;
  assign _T_3388 = _T_3386 ^ (* src = "crypto_accelerator.v:2327" *) _T_3384;
  assign _T_3392 = _T_3390 ^ (* src = "crypto_accelerator.v:2329" *) _T_3384;
  assign _T_3394 = _T_3368 ^ (* src = "crypto_accelerator.v:2330" *) _T_3366;
  assign _T_3396 = _T_3372 ^ (* src = "crypto_accelerator.v:2331" *) _T_3360;
  assign _T_3398 = _T_3378 ^ (* src = "crypto_accelerator.v:2332" *) _T_3376;
  assign _T_3400 = _T_3382 ^ (* src = "crypto_accelerator.v:2333" *) _T_3392;
  assign _T_3402 = _T_3394 ^ (* src = "crypto_accelerator.v:2334" *) _T_3388;
  assign _T_3404 = _T_3396 ^ (* src = "crypto_accelerator.v:2335" *) _T_3392;
  assign _T_3406 = _T_3398 ^ (* src = "crypto_accelerator.v:2336" *) _T_3388;
  assign _T_3408 = _T_3400 ^ (* src = "crypto_accelerator.v:2337" *) _T_3362;
  assign _T_3410 = _T_3406 ^ (* src = "crypto_accelerator.v:2338" *) _T_3408;
  assign _T_3414 = _T_3404 ^ (* src = "crypto_accelerator.v:2340" *) _T_3412;
  assign _T_3416 = _T_3402 ^ (* src = "crypto_accelerator.v:2341" *) _T_3404;
  assign _T_3418 = _T_3408 ^ (* src = "crypto_accelerator.v:2342" *) _T_3412;
  assign _T_3428 = _T_3416 ^ (* src = "crypto_accelerator.v:2347" *) _T_3412;
  assign _T_3434 = _T_3410 ^ (* src = "crypto_accelerator.v:2350" *) _T_3412;
  assign _T_3436 = _T_3404 ^ (* src = "crypto_accelerator.v:2351" *) _T_3420;
  assign _T_3438 = _T_3426 ^ (* src = "crypto_accelerator.v:2352" *) _T_3428;
  assign _T_3440 = _T_3408 ^ (* src = "crypto_accelerator.v:2353" *) _T_3422;
  assign _T_3442 = _T_3432 ^ (* src = "crypto_accelerator.v:2354" *) _T_3434;
  assign _T_3444 = _T_3438 ^ (* src = "crypto_accelerator.v:2355" *) _T_3442;
  assign _T_3446 = _T_3436 ^ (* src = "crypto_accelerator.v:2356" *) _T_3440;
  assign _T_3448 = _T_3436 ^ (* src = "crypto_accelerator.v:2357" *) _T_3438;
  assign _T_3450 = _T_3440 ^ (* src = "crypto_accelerator.v:2358" *) _T_3442;
  assign _T_3452 = _T_3446 ^ (* src = "crypto_accelerator.v:2359" *) _T_3444;
  assign _T_3490 = _T_3484 ^ (* src = "crypto_accelerator.v:2378" *) _T_3486;
  assign _T_3492 = _T_3462 ^ (* src = "crypto_accelerator.v:2379" *) _T_3474;
  assign _T_3494 = _T_3468 ^ (* src = "crypto_accelerator.v:2380" *) _T_3490;
  assign _T_3496 = _T_3472 ^ (* src = "crypto_accelerator.v:2381" *) _T_3492;
  assign _T_3498 = _T_3458 ^ (* src = "crypto_accelerator.v:2382" *) _T_3478;
  assign _T_3500 = _T_3454 ^ (* src = "crypto_accelerator.v:2383" *) _T_3460;
  assign _T_3502 = _T_3490 ^ (* src = "crypto_accelerator.v:2384" *) _T_3500;
  assign _T_3504 = _T_3456 ^ (* src = "crypto_accelerator.v:2385" *) _T_3496;
  assign _T_3506 = _T_3454 ^ (* src = "crypto_accelerator.v:2386" *) _T_3466;
  assign _T_3508 = _T_3464 ^ (* src = "crypto_accelerator.v:2387" *) _T_3480;
  assign _T_3510 = _T_3470 ^ (* src = "crypto_accelerator.v:2388" *) _T_3482;
  assign _T_3512 = _T_3458 ^ (* src = "crypto_accelerator.v:2389" *) _T_3504;
  assign _T_3514 = _T_3498 ^ (* src = "crypto_accelerator.v:2390" *) _T_3510;
  assign _T_3516 = _T_3476 ^ (* src = "crypto_accelerator.v:2391" *) _T_3492;
  assign _T_3518 = _T_3460 ^ (* src = "crypto_accelerator.v:2392" *) _T_3466;
  assign _T_3520 = _T_3496 ^ (* src = "crypto_accelerator.v:2393" *) _T_3518;
  assign _T_3522 = _T_3488 ^ (* src = "crypto_accelerator.v:2394" *) _T_3514;
  assign _T_3524 = _T_3484 ^ (* src = "crypto_accelerator.v:2395" *) _T_3506;
  assign _T_3526 = _T_3498 ^ (* src = "crypto_accelerator.v:2396" *) _T_3508;
  assign _T_3527 = _T_3494 ^ (* src = "crypto_accelerator.v:2397" *) _T_3520;
  assign _T_3528 = _T_3522 ^ (* src = "crypto_accelerator.v:2398" *) _T_3524;
  assign _T_3531 = _T_3464 ^ (* src = "crypto_accelerator.v:2400" *) _T_3490;
  assign _T_3532 = _T_3502 ^ (* src = "crypto_accelerator.v:2401" *) _T_3504;
  assign _T_3533 = _T_3512 ^ (* src = "crypto_accelerator.v:2402" *) _T_3531;
  assign _T_3535 = _T_3462 ^ (* src = "crypto_accelerator.v:2403" *) _T_3478;
  assign _T_3537 = _T_3500 ^ (* src = "crypto_accelerator.v:2404" *) _T_3516;
  assign _T_3538 = _T_3502 ^ (* src = "crypto_accelerator.v:2405" *) _T_3526;
  assign _T_3541 = _T_3470 ^ (* src = "crypto_accelerator.v:2407" *) _T_3508;
  assign _T_3543 = _T_3535 ^ (* src = "crypto_accelerator.v:2408" *) _T_3541;
  assign _T_3545 = _T_3462 ^ (* src = "crypto_accelerator.v:2409" *) _T_3506;
  assign _T_3546 = _T_3494 ^ (* src = "crypto_accelerator.v:2410" *) _T_3543;
  assign _T_3549 = _T_3514 ^ (* src = "crypto_accelerator.v:2412" *) _T_3537;
  assign _T_3550 = _T_3494 ^ (* src = "crypto_accelerator.v:2413" *) _T_3549;
  assign _T_3552 = _T_3504 ^ (* src = "crypto_accelerator.v:2414" *) _T_3545;
  assign _T_3553 = _T_3494 ^ (* src = "crypto_accelerator.v:2415" *) _T_3552;
  assign _T_3579 = matrix_3_1[1] ^ (* src = "crypto_accelerator.v:2418" *) matrix_3_1[3];
  assign _T_3581 = matrix_3_1[4] ^ (* src = "crypto_accelerator.v:2419" *) matrix_3_1[7];
  assign _T_3583 = matrix_3_1[6] ^ (* src = "crypto_accelerator.v:2420" *) matrix_3_1[5];
  assign _T_3585 = matrix_3_1[0] ^ (* src = "crypto_accelerator.v:2421" *) _T_3583;
  assign _T_3587 = _T_3579 ^ (* src = "crypto_accelerator.v:2422" *) _T_3581;
  assign _T_3589 = matrix_3_1[6] ^ (* src = "crypto_accelerator.v:2423" *) matrix_3_1[2];
  assign _T_3591 = matrix_3_1[7] ^ (* src = "crypto_accelerator.v:2424" *) matrix_3_1[1];
  assign _T_3593 = _T_3579 ^ (* src = "crypto_accelerator.v:2425" *) _T_3589;
  assign _T_3595 = matrix_3_1[1] ^ (* src = "crypto_accelerator.v:2426" *) _T_3585;
  assign _T_3597 = matrix_3_1[4] ^ (* src = "crypto_accelerator.v:2427" *) _T_3585;
  assign _T_3599 = matrix_3_1[0] ^ (* src = "crypto_accelerator.v:2428" *) _T_3587;
  assign _T_3601 = _T_3587 ^ (* src = "crypto_accelerator.v:2429" *) _T_3589;
  assign _T_3603 = matrix_3_1[5] ^ (* src = "crypto_accelerator.v:2430" *) matrix_3_1[2];
  assign _T_3605 = _T_3583 ^ (* src = "crypto_accelerator.v:2431" *) _T_3587;
  assign _T_3607 = matrix_3_1[2] ^ (* src = "crypto_accelerator.v:2432" *) _T_3591;
  assign _T_3609 = matrix_3_1[7] ^ (* src = "crypto_accelerator.v:2433" *) matrix_3_1[2];
  assign _T_3611 = matrix_3_1[0] ^ (* src = "crypto_accelerator.v:2434" *) _T_3593;
  assign _T_3613 = matrix_3_1[1] ^ (* src = "crypto_accelerator.v:2435" *) matrix_3_1[2];
  assign _T_3615 = _T_3581 ^ (* src = "crypto_accelerator.v:2436" *) _T_3613;
  assign _T_3617 = _T_3585 ^ (* src = "crypto_accelerator.v:2437" *) _T_3607;
  assign _T_3619 = _T_3579 ^ (* src = "crypto_accelerator.v:2438" *) _T_3603;
  assign _T_3621 = matrix_3_1[7] ^ (* src = "crypto_accelerator.v:2439" *) _T_3585;
  assign _T_3623 = _T_3619 ^ (* src = "crypto_accelerator.v:2440" *) _T_3587;
  assign _T_3625 = _T_3619 ^ (* src = "crypto_accelerator.v:2441" *) _T_3591;
  assign _T_3627 = _T_3591 ^ (* src = "crypto_accelerator.v:2442" *) _T_3615;
  assign _T_3629 = _T_3609 ^ (* src = "crypto_accelerator.v:2443" *) _T_3605;
  assign _T_3631 = _T_3621 ^ (* src = "crypto_accelerator.v:2444" *) _T_3611;
  assign _T_3637 = _T_3601 ^ (* src = "crypto_accelerator.v:2447" *) _T_3633;
  assign _T_3641 = _T_3639 ^ (* src = "crypto_accelerator.v:2449" *) _T_3633;
  assign _T_3647 = _T_3625 ^ (* src = "crypto_accelerator.v:2452" *) _T_3643;
  assign _T_3651 = _T_3649 ^ (* src = "crypto_accelerator.v:2454" *) _T_3643;
  assign _T_3657 = _T_3655 ^ (* src = "crypto_accelerator.v:2457" *) _T_3653;
  assign _T_3661 = _T_3659 ^ (* src = "crypto_accelerator.v:2459" *) _T_3653;
  assign _T_3663 = _T_3637 ^ (* src = "crypto_accelerator.v:2460" *) _T_3635;
  assign _T_3665 = _T_3641 ^ (* src = "crypto_accelerator.v:2461" *) _T_3629;
  assign _T_3667 = _T_3647 ^ (* src = "crypto_accelerator.v:2462" *) _T_3645;
  assign _T_3669 = _T_3651 ^ (* src = "crypto_accelerator.v:2463" *) _T_3661;
  assign _T_3671 = _T_3663 ^ (* src = "crypto_accelerator.v:2464" *) _T_3657;
  assign _T_3673 = _T_3665 ^ (* src = "crypto_accelerator.v:2465" *) _T_3661;
  assign _T_3675 = _T_3667 ^ (* src = "crypto_accelerator.v:2466" *) _T_3657;
  assign _T_3677 = _T_3669 ^ (* src = "crypto_accelerator.v:2467" *) _T_3631;
  assign _T_3679 = _T_3675 ^ (* src = "crypto_accelerator.v:2468" *) _T_3677;
  assign _T_3683 = _T_3673 ^ (* src = "crypto_accelerator.v:2470" *) _T_3681;
  assign _T_3685 = _T_3671 ^ (* src = "crypto_accelerator.v:2471" *) _T_3673;
  assign _T_3687 = _T_3677 ^ (* src = "crypto_accelerator.v:2472" *) _T_3681;
  assign _T_3697 = _T_3685 ^ (* src = "crypto_accelerator.v:2477" *) _T_3681;
  assign _T_3703 = _T_3679 ^ (* src = "crypto_accelerator.v:2480" *) _T_3681;
  assign _T_3705 = _T_3673 ^ (* src = "crypto_accelerator.v:2481" *) _T_3689;
  assign _T_3707 = _T_3695 ^ (* src = "crypto_accelerator.v:2482" *) _T_3697;
  assign _T_3709 = _T_3677 ^ (* src = "crypto_accelerator.v:2483" *) _T_3691;
  assign _T_3711 = _T_3701 ^ (* src = "crypto_accelerator.v:2484" *) _T_3703;
  assign _T_3713 = _T_3707 ^ (* src = "crypto_accelerator.v:2485" *) _T_3711;
  assign _T_3715 = _T_3705 ^ (* src = "crypto_accelerator.v:2486" *) _T_3709;
  assign _T_3717 = _T_3705 ^ (* src = "crypto_accelerator.v:2487" *) _T_3707;
  assign _T_3719 = _T_3709 ^ (* src = "crypto_accelerator.v:2488" *) _T_3711;
  assign _T_3721 = _T_3715 ^ (* src = "crypto_accelerator.v:2489" *) _T_3713;
  assign _T_3759 = _T_3753 ^ (* src = "crypto_accelerator.v:2508" *) _T_3755;
  assign _T_3761 = _T_3731 ^ (* src = "crypto_accelerator.v:2509" *) _T_3743;
  assign _T_3763 = _T_3737 ^ (* src = "crypto_accelerator.v:2510" *) _T_3759;
  assign _T_3765 = _T_3741 ^ (* src = "crypto_accelerator.v:2511" *) _T_3761;
  assign _T_3767 = _T_3727 ^ (* src = "crypto_accelerator.v:2512" *) _T_3747;
  assign _T_3769 = _T_3723 ^ (* src = "crypto_accelerator.v:2513" *) _T_3729;
  assign _T_3771 = _T_3759 ^ (* src = "crypto_accelerator.v:2514" *) _T_3769;
  assign _T_3773 = _T_3725 ^ (* src = "crypto_accelerator.v:2515" *) _T_3765;
  assign _T_3775 = _T_3723 ^ (* src = "crypto_accelerator.v:2516" *) _T_3735;
  assign _T_3777 = _T_3733 ^ (* src = "crypto_accelerator.v:2517" *) _T_3749;
  assign _T_3779 = _T_3739 ^ (* src = "crypto_accelerator.v:2518" *) _T_3751;
  assign _T_3781 = _T_3727 ^ (* src = "crypto_accelerator.v:2519" *) _T_3773;
  assign _T_3783 = _T_3767 ^ (* src = "crypto_accelerator.v:2520" *) _T_3779;
  assign _T_3785 = _T_3745 ^ (* src = "crypto_accelerator.v:2521" *) _T_3761;
  assign _T_3787 = _T_3729 ^ (* src = "crypto_accelerator.v:2522" *) _T_3735;
  assign _T_3789 = _T_3765 ^ (* src = "crypto_accelerator.v:2523" *) _T_3787;
  assign _T_3791 = _T_3757 ^ (* src = "crypto_accelerator.v:2524" *) _T_3783;
  assign _T_3793 = _T_3753 ^ (* src = "crypto_accelerator.v:2525" *) _T_3775;
  assign _T_3795 = _T_3767 ^ (* src = "crypto_accelerator.v:2526" *) _T_3777;
  assign _T_3796 = _T_3763 ^ (* src = "crypto_accelerator.v:2527" *) _T_3789;
  assign _T_3797 = _T_3791 ^ (* src = "crypto_accelerator.v:2528" *) _T_3793;
  assign _T_3800 = _T_3733 ^ (* src = "crypto_accelerator.v:2530" *) _T_3759;
  assign _T_3801 = _T_3771 ^ (* src = "crypto_accelerator.v:2531" *) _T_3773;
  assign _T_3802 = _T_3781 ^ (* src = "crypto_accelerator.v:2532" *) _T_3800;
  assign _T_3804 = _T_3731 ^ (* src = "crypto_accelerator.v:2533" *) _T_3747;
  assign _T_3806 = _T_3769 ^ (* src = "crypto_accelerator.v:2534" *) _T_3785;
  assign _T_3807 = _T_3771 ^ (* src = "crypto_accelerator.v:2535" *) _T_3795;
  assign _T_3810 = _T_3739 ^ (* src = "crypto_accelerator.v:2537" *) _T_3777;
  assign _T_3812 = _T_3804 ^ (* src = "crypto_accelerator.v:2538" *) _T_3810;
  assign _T_3814 = _T_3731 ^ (* src = "crypto_accelerator.v:2539" *) _T_3775;
  assign _T_3815 = _T_3763 ^ (* src = "crypto_accelerator.v:2540" *) _T_3812;
  assign _T_3818 = _T_3783 ^ (* src = "crypto_accelerator.v:2542" *) _T_3806;
  assign _T_3819 = _T_3763 ^ (* src = "crypto_accelerator.v:2543" *) _T_3818;
  assign _T_3821 = _T_3773 ^ (* src = "crypto_accelerator.v:2544" *) _T_3814;
  assign _T_3822 = _T_3763 ^ (* src = "crypto_accelerator.v:2545" *) _T_3821;
  assign _T_3848 = matrix_3_2[1] ^ (* src = "crypto_accelerator.v:2548" *) matrix_3_2[3];
  assign _T_3850 = matrix_3_2[4] ^ (* src = "crypto_accelerator.v:2549" *) matrix_3_2[7];
  assign _T_3852 = matrix_3_2[6] ^ (* src = "crypto_accelerator.v:2550" *) matrix_3_2[5];
  assign _T_3854 = matrix_3_2[0] ^ (* src = "crypto_accelerator.v:2551" *) _T_3852;
  assign _T_3856 = _T_3848 ^ (* src = "crypto_accelerator.v:2552" *) _T_3850;
  assign _T_3858 = matrix_3_2[6] ^ (* src = "crypto_accelerator.v:2553" *) matrix_3_2[2];
  assign _T_3860 = matrix_3_2[7] ^ (* src = "crypto_accelerator.v:2554" *) matrix_3_2[1];
  assign _T_3862 = _T_3848 ^ (* src = "crypto_accelerator.v:2555" *) _T_3858;
  assign _T_3864 = matrix_3_2[1] ^ (* src = "crypto_accelerator.v:2556" *) _T_3854;
  assign _T_3866 = matrix_3_2[4] ^ (* src = "crypto_accelerator.v:2557" *) _T_3854;
  assign _T_3868 = matrix_3_2[0] ^ (* src = "crypto_accelerator.v:2558" *) _T_3856;
  assign _T_3870 = _T_3856 ^ (* src = "crypto_accelerator.v:2559" *) _T_3858;
  assign _T_3872 = matrix_3_2[5] ^ (* src = "crypto_accelerator.v:2560" *) matrix_3_2[2];
  assign _T_3874 = _T_3852 ^ (* src = "crypto_accelerator.v:2561" *) _T_3856;
  assign _T_3876 = matrix_3_2[2] ^ (* src = "crypto_accelerator.v:2562" *) _T_3860;
  assign _T_3878 = matrix_3_2[7] ^ (* src = "crypto_accelerator.v:2563" *) matrix_3_2[2];
  assign _T_3880 = matrix_3_2[0] ^ (* src = "crypto_accelerator.v:2564" *) _T_3862;
  assign _T_3882 = matrix_3_2[1] ^ (* src = "crypto_accelerator.v:2565" *) matrix_3_2[2];
  assign _T_3884 = _T_3850 ^ (* src = "crypto_accelerator.v:2566" *) _T_3882;
  assign _T_3886 = _T_3854 ^ (* src = "crypto_accelerator.v:2567" *) _T_3876;
  assign _T_3888 = _T_3848 ^ (* src = "crypto_accelerator.v:2568" *) _T_3872;
  assign _T_3890 = matrix_3_2[7] ^ (* src = "crypto_accelerator.v:2569" *) _T_3854;
  assign _T_3892 = _T_3888 ^ (* src = "crypto_accelerator.v:2570" *) _T_3856;
  assign _T_3894 = _T_3888 ^ (* src = "crypto_accelerator.v:2571" *) _T_3860;
  assign _T_3896 = _T_3860 ^ (* src = "crypto_accelerator.v:2572" *) _T_3884;
  assign _T_3898 = _T_3878 ^ (* src = "crypto_accelerator.v:2573" *) _T_3874;
  assign _T_3900 = _T_3890 ^ (* src = "crypto_accelerator.v:2574" *) _T_3880;
  assign _T_3906 = _T_3870 ^ (* src = "crypto_accelerator.v:2577" *) _T_3902;
  assign _T_3910 = _T_3908 ^ (* src = "crypto_accelerator.v:2579" *) _T_3902;
  assign _T_3916 = _T_3894 ^ (* src = "crypto_accelerator.v:2582" *) _T_3912;
  assign _T_3920 = _T_3918 ^ (* src = "crypto_accelerator.v:2584" *) _T_3912;
  assign _T_3926 = _T_3924 ^ (* src = "crypto_accelerator.v:2587" *) _T_3922;
  assign _T_3930 = _T_3928 ^ (* src = "crypto_accelerator.v:2589" *) _T_3922;
  assign _T_3932 = _T_3906 ^ (* src = "crypto_accelerator.v:2590" *) _T_3904;
  assign _T_3934 = _T_3910 ^ (* src = "crypto_accelerator.v:2591" *) _T_3898;
  assign _T_3936 = _T_3916 ^ (* src = "crypto_accelerator.v:2592" *) _T_3914;
  assign _T_3938 = _T_3920 ^ (* src = "crypto_accelerator.v:2593" *) _T_3930;
  assign _T_3940 = _T_3932 ^ (* src = "crypto_accelerator.v:2594" *) _T_3926;
  assign _T_3942 = _T_3934 ^ (* src = "crypto_accelerator.v:2595" *) _T_3930;
  assign _T_3944 = _T_3936 ^ (* src = "crypto_accelerator.v:2596" *) _T_3926;
  assign _T_3946 = _T_3938 ^ (* src = "crypto_accelerator.v:2597" *) _T_3900;
  assign _T_3948 = _T_3944 ^ (* src = "crypto_accelerator.v:2598" *) _T_3946;
  assign _T_3952 = _T_3942 ^ (* src = "crypto_accelerator.v:2600" *) _T_3950;
  assign _T_3954 = _T_3940 ^ (* src = "crypto_accelerator.v:2601" *) _T_3942;
  assign _T_3956 = _T_3946 ^ (* src = "crypto_accelerator.v:2602" *) _T_3950;
  assign _T_3966 = _T_3954 ^ (* src = "crypto_accelerator.v:2607" *) _T_3950;
  assign _T_3972 = _T_3948 ^ (* src = "crypto_accelerator.v:2610" *) _T_3950;
  assign _T_3974 = _T_3942 ^ (* src = "crypto_accelerator.v:2611" *) _T_3958;
  assign _T_3976 = _T_3964 ^ (* src = "crypto_accelerator.v:2612" *) _T_3966;
  assign _T_3978 = _T_3946 ^ (* src = "crypto_accelerator.v:2613" *) _T_3960;
  assign _T_3980 = _T_3970 ^ (* src = "crypto_accelerator.v:2614" *) _T_3972;
  assign _T_3982 = _T_3976 ^ (* src = "crypto_accelerator.v:2615" *) _T_3980;
  assign _T_3984 = _T_3974 ^ (* src = "crypto_accelerator.v:2616" *) _T_3978;
  assign _T_3986 = _T_3974 ^ (* src = "crypto_accelerator.v:2617" *) _T_3976;
  assign _T_3988 = _T_3978 ^ (* src = "crypto_accelerator.v:2618" *) _T_3980;
  assign _T_3990 = _T_3984 ^ (* src = "crypto_accelerator.v:2619" *) _T_3982;
  assign _T_4028 = _T_4022 ^ (* src = "crypto_accelerator.v:2638" *) _T_4024;
  assign _T_4030 = _T_4000 ^ (* src = "crypto_accelerator.v:2639" *) _T_4012;
  assign _T_4032 = _T_4006 ^ (* src = "crypto_accelerator.v:2640" *) _T_4028;
  assign _T_4034 = _T_4010 ^ (* src = "crypto_accelerator.v:2641" *) _T_4030;
  assign _T_4036 = _T_3996 ^ (* src = "crypto_accelerator.v:2642" *) _T_4016;
  assign _T_4038 = _T_3992 ^ (* src = "crypto_accelerator.v:2643" *) _T_3998;
  assign _T_4040 = _T_4028 ^ (* src = "crypto_accelerator.v:2644" *) _T_4038;
  assign _T_4042 = _T_3994 ^ (* src = "crypto_accelerator.v:2645" *) _T_4034;
  assign _T_4044 = _T_3992 ^ (* src = "crypto_accelerator.v:2646" *) _T_4004;
  assign _T_4046 = _T_4002 ^ (* src = "crypto_accelerator.v:2647" *) _T_4018;
  assign _T_4048 = _T_4008 ^ (* src = "crypto_accelerator.v:2648" *) _T_4020;
  assign _T_4050 = _T_3996 ^ (* src = "crypto_accelerator.v:2649" *) _T_4042;
  assign _T_4052 = _T_4036 ^ (* src = "crypto_accelerator.v:2650" *) _T_4048;
  assign _T_4054 = _T_4014 ^ (* src = "crypto_accelerator.v:2651" *) _T_4030;
  assign _T_4056 = _T_3998 ^ (* src = "crypto_accelerator.v:2652" *) _T_4004;
  assign _T_4058 = _T_4034 ^ (* src = "crypto_accelerator.v:2653" *) _T_4056;
  assign _T_4060 = _T_4026 ^ (* src = "crypto_accelerator.v:2654" *) _T_4052;
  assign _T_4062 = _T_4022 ^ (* src = "crypto_accelerator.v:2655" *) _T_4044;
  assign _T_4064 = _T_4036 ^ (* src = "crypto_accelerator.v:2656" *) _T_4046;
  assign _T_4065 = _T_4032 ^ (* src = "crypto_accelerator.v:2657" *) _T_4058;
  assign _T_4066 = _T_4060 ^ (* src = "crypto_accelerator.v:2658" *) _T_4062;
  assign _T_4069 = _T_4002 ^ (* src = "crypto_accelerator.v:2660" *) _T_4028;
  assign _T_4070 = _T_4040 ^ (* src = "crypto_accelerator.v:2661" *) _T_4042;
  assign _T_4071 = _T_4050 ^ (* src = "crypto_accelerator.v:2662" *) _T_4069;
  assign _T_4073 = _T_4000 ^ (* src = "crypto_accelerator.v:2663" *) _T_4016;
  assign _T_4075 = _T_4038 ^ (* src = "crypto_accelerator.v:2664" *) _T_4054;
  assign _T_4076 = _T_4040 ^ (* src = "crypto_accelerator.v:2665" *) _T_4064;
  assign _T_4079 = _T_4008 ^ (* src = "crypto_accelerator.v:2667" *) _T_4046;
  assign _T_4081 = _T_4073 ^ (* src = "crypto_accelerator.v:2668" *) _T_4079;
  assign _T_4083 = _T_4000 ^ (* src = "crypto_accelerator.v:2669" *) _T_4044;
  assign _T_4084 = _T_4032 ^ (* src = "crypto_accelerator.v:2670" *) _T_4081;
  assign _T_4087 = _T_4052 ^ (* src = "crypto_accelerator.v:2672" *) _T_4075;
  assign _T_4088 = _T_4032 ^ (* src = "crypto_accelerator.v:2673" *) _T_4087;
  assign _T_4090 = _T_4042 ^ (* src = "crypto_accelerator.v:2674" *) _T_4083;
  assign _T_4091 = _T_4032 ^ (* src = "crypto_accelerator.v:2675" *) _T_4090;
  assign _T_4117 = matrix_3_3[1] ^ (* src = "crypto_accelerator.v:2678" *) matrix_3_3[3];
  assign _T_4119 = matrix_3_3[4] ^ (* src = "crypto_accelerator.v:2679" *) matrix_3_3[7];
  assign _T_4121 = matrix_3_3[6] ^ (* src = "crypto_accelerator.v:2680" *) matrix_3_3[5];
  assign _T_4123 = matrix_3_3[0] ^ (* src = "crypto_accelerator.v:2681" *) _T_4121;
  assign _T_4125 = _T_4117 ^ (* src = "crypto_accelerator.v:2682" *) _T_4119;
  assign _T_4127 = matrix_3_3[6] ^ (* src = "crypto_accelerator.v:2683" *) matrix_3_3[2];
  assign _T_4129 = matrix_3_3[7] ^ (* src = "crypto_accelerator.v:2684" *) matrix_3_3[1];
  assign _T_4131 = _T_4117 ^ (* src = "crypto_accelerator.v:2685" *) _T_4127;
  assign _T_4133 = matrix_3_3[1] ^ (* src = "crypto_accelerator.v:2686" *) _T_4123;
  assign _T_4135 = matrix_3_3[4] ^ (* src = "crypto_accelerator.v:2687" *) _T_4123;
  assign _T_4137 = matrix_3_3[0] ^ (* src = "crypto_accelerator.v:2688" *) _T_4125;
  assign _T_4139 = _T_4125 ^ (* src = "crypto_accelerator.v:2689" *) _T_4127;
  assign _T_4141 = matrix_3_3[5] ^ (* src = "crypto_accelerator.v:2690" *) matrix_3_3[2];
  assign _T_4143 = _T_4121 ^ (* src = "crypto_accelerator.v:2691" *) _T_4125;
  assign _T_4145 = matrix_3_3[2] ^ (* src = "crypto_accelerator.v:2692" *) _T_4129;
  assign _T_4147 = matrix_3_3[7] ^ (* src = "crypto_accelerator.v:2693" *) matrix_3_3[2];
  assign _T_4149 = matrix_3_3[0] ^ (* src = "crypto_accelerator.v:2694" *) _T_4131;
  assign _T_4151 = matrix_3_3[1] ^ (* src = "crypto_accelerator.v:2695" *) matrix_3_3[2];
  assign _T_4153 = _T_4119 ^ (* src = "crypto_accelerator.v:2696" *) _T_4151;
  assign _T_4155 = _T_4123 ^ (* src = "crypto_accelerator.v:2697" *) _T_4145;
  assign _T_4157 = _T_4117 ^ (* src = "crypto_accelerator.v:2698" *) _T_4141;
  assign _T_4159 = matrix_3_3[7] ^ (* src = "crypto_accelerator.v:2699" *) _T_4123;
  assign _T_4161 = _T_4157 ^ (* src = "crypto_accelerator.v:2700" *) _T_4125;
  assign _T_4163 = _T_4157 ^ (* src = "crypto_accelerator.v:2701" *) _T_4129;
  assign _T_4165 = _T_4129 ^ (* src = "crypto_accelerator.v:2702" *) _T_4153;
  assign _T_4167 = _T_4147 ^ (* src = "crypto_accelerator.v:2703" *) _T_4143;
  assign _T_4169 = _T_4159 ^ (* src = "crypto_accelerator.v:2704" *) _T_4149;
  assign _T_4175 = _T_4139 ^ (* src = "crypto_accelerator.v:2707" *) _T_4171;
  assign _T_4179 = _T_4177 ^ (* src = "crypto_accelerator.v:2709" *) _T_4171;
  assign _T_4185 = _T_4163 ^ (* src = "crypto_accelerator.v:2712" *) _T_4181;
  assign _T_4189 = _T_4187 ^ (* src = "crypto_accelerator.v:2714" *) _T_4181;
  assign _T_4195 = _T_4193 ^ (* src = "crypto_accelerator.v:2717" *) _T_4191;
  assign _T_4199 = _T_4197 ^ (* src = "crypto_accelerator.v:2719" *) _T_4191;
  assign _T_4201 = _T_4175 ^ (* src = "crypto_accelerator.v:2720" *) _T_4173;
  assign _T_4203 = _T_4179 ^ (* src = "crypto_accelerator.v:2721" *) _T_4167;
  assign _T_4205 = _T_4185 ^ (* src = "crypto_accelerator.v:2722" *) _T_4183;
  assign _T_4207 = _T_4189 ^ (* src = "crypto_accelerator.v:2723" *) _T_4199;
  assign _T_4209 = _T_4201 ^ (* src = "crypto_accelerator.v:2724" *) _T_4195;
  assign _T_4211 = _T_4203 ^ (* src = "crypto_accelerator.v:2725" *) _T_4199;
  assign _T_4213 = _T_4205 ^ (* src = "crypto_accelerator.v:2726" *) _T_4195;
  assign _T_4215 = _T_4207 ^ (* src = "crypto_accelerator.v:2727" *) _T_4169;
  assign _T_4217 = _T_4213 ^ (* src = "crypto_accelerator.v:2728" *) _T_4215;
  assign _T_4221 = _T_4211 ^ (* src = "crypto_accelerator.v:2730" *) _T_4219;
  assign _T_4223 = _T_4209 ^ (* src = "crypto_accelerator.v:2731" *) _T_4211;
  assign _T_4225 = _T_4215 ^ (* src = "crypto_accelerator.v:2732" *) _T_4219;
  assign _T_4235 = _T_4223 ^ (* src = "crypto_accelerator.v:2737" *) _T_4219;
  assign _T_4241 = _T_4217 ^ (* src = "crypto_accelerator.v:2740" *) _T_4219;
  assign _T_4243 = _T_4211 ^ (* src = "crypto_accelerator.v:2741" *) _T_4227;
  assign _T_4245 = _T_4233 ^ (* src = "crypto_accelerator.v:2742" *) _T_4235;
  assign _T_4247 = _T_4215 ^ (* src = "crypto_accelerator.v:2743" *) _T_4229;
  assign _T_4249 = _T_4239 ^ (* src = "crypto_accelerator.v:2744" *) _T_4241;
  assign _T_4251 = _T_4245 ^ (* src = "crypto_accelerator.v:2745" *) _T_4249;
  assign _T_4253 = _T_4243 ^ (* src = "crypto_accelerator.v:2746" *) _T_4247;
  assign _T_4255 = _T_4243 ^ (* src = "crypto_accelerator.v:2747" *) _T_4245;
  assign _T_4257 = _T_4247 ^ (* src = "crypto_accelerator.v:2748" *) _T_4249;
  assign _T_4259 = _T_4253 ^ (* src = "crypto_accelerator.v:2749" *) _T_4251;
  assign _T_4297 = _T_4291 ^ (* src = "crypto_accelerator.v:2768" *) _T_4293;
  assign _T_4299 = _T_4269 ^ (* src = "crypto_accelerator.v:2769" *) _T_4281;
  assign _T_4301 = _T_4275 ^ (* src = "crypto_accelerator.v:2770" *) _T_4297;
  assign _T_4303 = _T_4279 ^ (* src = "crypto_accelerator.v:2771" *) _T_4299;
  assign _T_4305 = _T_4265 ^ (* src = "crypto_accelerator.v:2772" *) _T_4285;
  assign _T_4307 = _T_4261 ^ (* src = "crypto_accelerator.v:2773" *) _T_4267;
  assign _T_4309 = _T_4297 ^ (* src = "crypto_accelerator.v:2774" *) _T_4307;
  assign _T_4311 = _T_4263 ^ (* src = "crypto_accelerator.v:2775" *) _T_4303;
  assign _T_4313 = _T_4261 ^ (* src = "crypto_accelerator.v:2776" *) _T_4273;
  assign _T_4315 = _T_4271 ^ (* src = "crypto_accelerator.v:2777" *) _T_4287;
  assign _T_4317 = _T_4277 ^ (* src = "crypto_accelerator.v:2778" *) _T_4289;
  assign _T_4319 = _T_4265 ^ (* src = "crypto_accelerator.v:2779" *) _T_4311;
  assign _T_4321 = _T_4305 ^ (* src = "crypto_accelerator.v:2780" *) _T_4317;
  assign _T_4323 = _T_4283 ^ (* src = "crypto_accelerator.v:2781" *) _T_4299;
  assign _T_4325 = _T_4267 ^ (* src = "crypto_accelerator.v:2782" *) _T_4273;
  assign _T_4327 = _T_4303 ^ (* src = "crypto_accelerator.v:2783" *) _T_4325;
  assign _T_4329 = _T_4295 ^ (* src = "crypto_accelerator.v:2784" *) _T_4321;
  assign _T_4331 = _T_4291 ^ (* src = "crypto_accelerator.v:2785" *) _T_4313;
  assign _T_4333 = _T_4305 ^ (* src = "crypto_accelerator.v:2786" *) _T_4315;
  assign _T_4334 = _T_4301 ^ (* src = "crypto_accelerator.v:2787" *) _T_4327;
  assign _T_4335 = _T_4329 ^ (* src = "crypto_accelerator.v:2788" *) _T_4331;
  assign _T_4338 = _T_4271 ^ (* src = "crypto_accelerator.v:2790" *) _T_4297;
  assign _T_4339 = _T_4309 ^ (* src = "crypto_accelerator.v:2791" *) _T_4311;
  assign _T_4340 = _T_4319 ^ (* src = "crypto_accelerator.v:2792" *) _T_4338;
  assign _T_4342 = _T_4269 ^ (* src = "crypto_accelerator.v:2793" *) _T_4285;
  assign _T_4344 = _T_4307 ^ (* src = "crypto_accelerator.v:2794" *) _T_4323;
  assign _T_4345 = _T_4309 ^ (* src = "crypto_accelerator.v:2795" *) _T_4333;
  assign _T_4348 = _T_4277 ^ (* src = "crypto_accelerator.v:2797" *) _T_4315;
  assign _T_4350 = _T_4342 ^ (* src = "crypto_accelerator.v:2798" *) _T_4348;
  assign _T_4352 = _T_4269 ^ (* src = "crypto_accelerator.v:2799" *) _T_4313;
  assign _T_4353 = _T_4301 ^ (* src = "crypto_accelerator.v:2800" *) _T_4350;
  assign _T_4356 = _T_4321 ^ (* src = "crypto_accelerator.v:2802" *) _T_4344;
  assign _T_4357 = _T_4301 ^ (* src = "crypto_accelerator.v:2803" *) _T_4356;
  assign _T_4359 = _T_4311 ^ (* src = "crypto_accelerator.v:2804" *) _T_4352;
  assign _T_4360 = _T_4301 ^ (* src = "crypto_accelerator.v:2805" *) _T_4359;
  assign roundPart2_0_0 = MixColsModule_io_out_0_0 ^ (* src = "crypto_accelerator.v:2808" *) io_keys_0_0_0;
  assign roundPart2_0_1 = MixColsModule_io_out_0_1 ^ (* src = "crypto_accelerator.v:2809" *) io_keys_0_0_1;
  assign roundPart2_0_2 = MixColsModule_io_out_0_2 ^ (* src = "crypto_accelerator.v:2810" *) io_keys_0_0_2;
  assign roundPart2_0_3 = MixColsModule_io_out_0_3 ^ (* src = "crypto_accelerator.v:2811" *) io_keys_0_0_3;
  assign roundPart2_1_0 = MixColsModule_io_out_1_0 ^ (* src = "crypto_accelerator.v:2812" *) io_keys_0_1_0;
  assign roundPart2_1_1 = MixColsModule_io_out_1_1 ^ (* src = "crypto_accelerator.v:2813" *) io_keys_0_1_1;
  assign roundPart2_1_2 = MixColsModule_io_out_1_2 ^ (* src = "crypto_accelerator.v:2814" *) io_keys_0_1_2;
  assign roundPart2_1_3 = MixColsModule_io_out_1_3 ^ (* src = "crypto_accelerator.v:2815" *) io_keys_0_1_3;
  assign roundPart2_2_0 = MixColsModule_io_out_2_0 ^ (* src = "crypto_accelerator.v:2816" *) io_keys_0_2_0;
  assign roundPart2_2_1 = MixColsModule_io_out_2_1 ^ (* src = "crypto_accelerator.v:2817" *) io_keys_0_2_1;
  assign roundPart2_2_2 = MixColsModule_io_out_2_2 ^ (* src = "crypto_accelerator.v:2818" *) io_keys_0_2_2;
  assign roundPart2_2_3 = MixColsModule_io_out_2_3 ^ (* src = "crypto_accelerator.v:2819" *) io_keys_0_2_3;
  assign roundPart2_3_0 = MixColsModule_io_out_3_0 ^ (* src = "crypto_accelerator.v:2820" *) io_keys_0_3_0;
  assign roundPart2_3_1 = MixColsModule_io_out_3_1 ^ (* src = "crypto_accelerator.v:2821" *) io_keys_0_3_1;
  assign roundPart2_3_2 = MixColsModule_io_out_3_2 ^ (* src = "crypto_accelerator.v:2822" *) io_keys_0_3_2;
  assign roundPart2_3_3 = MixColsModule_io_out_3_3 ^ (* src = "crypto_accelerator.v:2823" *) io_keys_0_3_3;
  assign roundPart2_last_0_0 = matrix_0_0 ^ (* src = "crypto_accelerator.v:2824" *) io_keys_0_0_0;
  assign roundPart2_last_0_1 = matrix_0_1 ^ (* src = "crypto_accelerator.v:2825" *) io_keys_0_0_1;
  assign roundPart2_last_0_2 = matrix_0_2 ^ (* src = "crypto_accelerator.v:2826" *) io_keys_0_0_2;
  assign roundPart2_last_0_3 = matrix_0_3 ^ (* src = "crypto_accelerator.v:2827" *) io_keys_0_0_3;
  assign roundPart2_last_1_0 = matrix_1_0 ^ (* src = "crypto_accelerator.v:2828" *) io_keys_0_1_0;
  assign roundPart2_last_1_1 = matrix_1_1 ^ (* src = "crypto_accelerator.v:2829" *) io_keys_0_1_1;
  assign roundPart2_last_1_2 = matrix_1_2 ^ (* src = "crypto_accelerator.v:2830" *) io_keys_0_1_2;
  assign roundPart2_last_1_3 = matrix_1_3 ^ (* src = "crypto_accelerator.v:2831" *) io_keys_0_1_3;
  assign roundPart2_last_2_0 = matrix_2_0 ^ (* src = "crypto_accelerator.v:2832" *) io_keys_0_2_0;
  assign roundPart2_last_2_1 = matrix_2_1 ^ (* src = "crypto_accelerator.v:2833" *) io_keys_0_2_1;
  assign roundPart2_last_2_2 = matrix_2_2 ^ (* src = "crypto_accelerator.v:2834" *) io_keys_0_2_2;
  assign roundPart2_last_2_3 = matrix_2_3 ^ (* src = "crypto_accelerator.v:2835" *) io_keys_0_2_3;
  assign roundPart2_last_3_0 = matrix_3_0 ^ (* src = "crypto_accelerator.v:2836" *) io_keys_0_3_0;
  assign roundPart2_last_3_1 = matrix_3_1 ^ (* src = "crypto_accelerator.v:2837" *) io_keys_0_3_1;
  assign roundPart2_last_3_2 = matrix_3_2 ^ (* src = "crypto_accelerator.v:2838" *) io_keys_0_3_2;
  assign roundPart2_last_3_3 = matrix_3_3 ^ (* src = "crypto_accelerator.v:2839" *) io_keys_0_3_3;
  assign _T_25 = io_dataIn ^ (* src = "crypto_accelerator.v:708" *) io_ivIn;
  assign _T_41 = _T_25 ^ (* src = "crypto_accelerator.v:711" *) { io_keys_0_0_0, io_keys_0_0_1, io_keys_0_0_2, io_keys_0_0_3, io_keys_0_1_0, io_keys_0_1_1, io_keys_0_1_2, io_keys_0_1_3, io_keys_0_2_0, io_keys_0_2_1, io_keys_0_2_2, io_keys_0_2_3, io_keys_0_3_0, io_keys_0_3_1, io_keys_0_3_2, io_keys_0_3_3 };
  assign _T_79 = matrix_0_0[1] ^ (* src = "crypto_accelerator.v:728" *) matrix_0_0[3];
  assign _T_81 = matrix_0_0[4] ^ (* src = "crypto_accelerator.v:729" *) matrix_0_0[7];
  assign _T_83 = matrix_0_0[6] ^ (* src = "crypto_accelerator.v:730" *) matrix_0_0[5];
  assign _T_85 = matrix_0_0[0] ^ (* src = "crypto_accelerator.v:731" *) _T_83;
  assign _T_87 = _T_79 ^ (* src = "crypto_accelerator.v:732" *) _T_81;
  assign _T_89 = matrix_0_0[6] ^ (* src = "crypto_accelerator.v:733" *) matrix_0_0[2];
  assign _T_91 = matrix_0_0[7] ^ (* src = "crypto_accelerator.v:734" *) matrix_0_0[1];
  assign _T_93 = _T_79 ^ (* src = "crypto_accelerator.v:735" *) _T_89;
  assign _T_95 = matrix_0_0[1] ^ (* src = "crypto_accelerator.v:736" *) _T_85;
  assign _T_97 = matrix_0_0[4] ^ (* src = "crypto_accelerator.v:737" *) _T_85;
  assign _T_99 = matrix_0_0[0] ^ (* src = "crypto_accelerator.v:738" *) _T_87;
  assign _T_101 = _T_87 ^ (* src = "crypto_accelerator.v:739" *) _T_89;
  assign _T_103 = matrix_0_0[5] ^ (* src = "crypto_accelerator.v:740" *) matrix_0_0[2];
  assign _T_105 = _T_83 ^ (* src = "crypto_accelerator.v:741" *) _T_87;
  assign _T_107 = matrix_0_0[2] ^ (* src = "crypto_accelerator.v:742" *) _T_91;
  assign _T_109 = matrix_0_0[7] ^ (* src = "crypto_accelerator.v:743" *) matrix_0_0[2];
  assign _T_111 = matrix_0_0[0] ^ (* src = "crypto_accelerator.v:744" *) _T_93;
  assign _T_113 = matrix_0_0[1] ^ (* src = "crypto_accelerator.v:745" *) matrix_0_0[2];
  assign _T_115 = _T_81 ^ (* src = "crypto_accelerator.v:746" *) _T_113;
  assign _T_117 = _T_85 ^ (* src = "crypto_accelerator.v:747" *) _T_107;
  assign _T_119 = _T_79 ^ (* src = "crypto_accelerator.v:748" *) _T_103;
  assign _T_121 = matrix_0_0[7] ^ (* src = "crypto_accelerator.v:749" *) _T_85;
  assign _T_123 = _T_119 ^ (* src = "crypto_accelerator.v:750" *) _T_87;
  assign _T_125 = _T_119 ^ (* src = "crypto_accelerator.v:751" *) _T_91;
  assign _T_127 = _T_91 ^ (* src = "crypto_accelerator.v:752" *) _T_115;
  assign _T_129 = _T_109 ^ (* src = "crypto_accelerator.v:753" *) _T_105;
  assign _T_131 = _T_121 ^ (* src = "crypto_accelerator.v:754" *) _T_111;
  assign _T_137 = _T_101 ^ (* src = "crypto_accelerator.v:757" *) _T_133;
  assign _T_141 = _T_139 ^ (* src = "crypto_accelerator.v:759" *) _T_133;
  assign _T_147 = _T_125 ^ (* src = "crypto_accelerator.v:762" *) _T_143;
  assign _T_151 = _T_149 ^ (* src = "crypto_accelerator.v:764" *) _T_143;
  assign _T_157 = _T_155 ^ (* src = "crypto_accelerator.v:767" *) _T_153;
  assign _T_161 = _T_159 ^ (* src = "crypto_accelerator.v:769" *) _T_153;
  assign _T_163 = _T_137 ^ (* src = "crypto_accelerator.v:770" *) _T_135;
  assign _T_165 = _T_141 ^ (* src = "crypto_accelerator.v:771" *) _T_129;
  assign _T_167 = _T_147 ^ (* src = "crypto_accelerator.v:772" *) _T_145;
  assign _T_169 = _T_151 ^ (* src = "crypto_accelerator.v:773" *) _T_161;
  assign _T_171 = _T_163 ^ (* src = "crypto_accelerator.v:774" *) _T_157;
  assign _T_173 = _T_165 ^ (* src = "crypto_accelerator.v:775" *) _T_161;
  assign _T_175 = _T_167 ^ (* src = "crypto_accelerator.v:776" *) _T_157;
  assign _T_177 = _T_169 ^ (* src = "crypto_accelerator.v:777" *) _T_131;
  assign _T_179 = _T_175 ^ (* src = "crypto_accelerator.v:778" *) _T_177;
  assign _T_183 = _T_173 ^ (* src = "crypto_accelerator.v:780" *) _T_181;
  assign _T_185 = _T_171 ^ (* src = "crypto_accelerator.v:781" *) _T_173;
  assign _T_187 = _T_177 ^ (* src = "crypto_accelerator.v:782" *) _T_181;
  assign _T_197 = _T_185 ^ (* src = "crypto_accelerator.v:787" *) _T_181;
  assign _T_203 = _T_179 ^ (* src = "crypto_accelerator.v:790" *) _T_181;
  assign _T_205 = _T_173 ^ (* src = "crypto_accelerator.v:791" *) _T_189;
  assign _T_207 = _T_195 ^ (* src = "crypto_accelerator.v:792" *) _T_197;
  assign _T_209 = _T_177 ^ (* src = "crypto_accelerator.v:793" *) _T_191;
  assign _T_211 = _T_201 ^ (* src = "crypto_accelerator.v:794" *) _T_203;
  assign _T_213 = _T_207 ^ (* src = "crypto_accelerator.v:795" *) _T_211;
  assign _T_215 = _T_205 ^ (* src = "crypto_accelerator.v:796" *) _T_209;
  assign _T_217 = _T_205 ^ (* src = "crypto_accelerator.v:797" *) _T_207;
  assign _T_219 = _T_209 ^ (* src = "crypto_accelerator.v:798" *) _T_211;
  assign _T_221 = _T_215 ^ (* src = "crypto_accelerator.v:799" *) _T_213;
  assign _T_259 = _T_253 ^ (* src = "crypto_accelerator.v:818" *) _T_255;
  assign _T_261 = _T_231 ^ (* src = "crypto_accelerator.v:819" *) _T_243;
  assign _T_263 = _T_237 ^ (* src = "crypto_accelerator.v:820" *) _T_259;
  assign _T_265 = _T_241 ^ (* src = "crypto_accelerator.v:821" *) _T_261;
  assign _T_267 = _T_227 ^ (* src = "crypto_accelerator.v:822" *) _T_247;
  assign _T_269 = _T_223 ^ (* src = "crypto_accelerator.v:823" *) _T_229;
  assign _T_271 = _T_259 ^ (* src = "crypto_accelerator.v:824" *) _T_269;
  assign _T_273 = _T_225 ^ (* src = "crypto_accelerator.v:825" *) _T_265;
  assign _T_275 = _T_223 ^ (* src = "crypto_accelerator.v:826" *) _T_235;
  assign _T_277 = _T_233 ^ (* src = "crypto_accelerator.v:827" *) _T_249;
  assign _T_279 = _T_239 ^ (* src = "crypto_accelerator.v:828" *) _T_251;
  assign _T_281 = _T_227 ^ (* src = "crypto_accelerator.v:829" *) _T_273;
  assign _T_283 = _T_267 ^ (* src = "crypto_accelerator.v:830" *) _T_279;
  assign _T_285 = _T_245 ^ (* src = "crypto_accelerator.v:831" *) _T_261;
  assign _T_287 = _T_229 ^ (* src = "crypto_accelerator.v:832" *) _T_235;
  assign _T_289 = _T_265 ^ (* src = "crypto_accelerator.v:833" *) _T_287;
  assign _T_291 = _T_257 ^ (* src = "crypto_accelerator.v:834" *) _T_283;
  assign _T_293 = _T_253 ^ (* src = "crypto_accelerator.v:835" *) _T_275;
  assign _T_295 = _T_267 ^ (* src = "crypto_accelerator.v:836" *) _T_277;
  assign _T_296 = _T_263 ^ (* src = "crypto_accelerator.v:837" *) _T_289;
  assign _T_297 = _T_291 ^ (* src = "crypto_accelerator.v:838" *) _T_293;
  assign _T_300 = _T_233 ^ (* src = "crypto_accelerator.v:840" *) _T_259;
  assign _T_301 = _T_271 ^ (* src = "crypto_accelerator.v:841" *) _T_273;
  assign _T_302 = _T_281 ^ (* src = "crypto_accelerator.v:842" *) _T_300;
  assign _T_304 = _T_231 ^ (* src = "crypto_accelerator.v:843" *) _T_247;
  assign _T_306 = _T_269 ^ (* src = "crypto_accelerator.v:844" *) _T_285;
  assign _T_307 = _T_271 ^ (* src = "crypto_accelerator.v:845" *) _T_295;
  assign _T_310 = _T_239 ^ (* src = "crypto_accelerator.v:847" *) _T_277;
  assign _T_312 = _T_304 ^ (* src = "crypto_accelerator.v:848" *) _T_310;
  assign _T_314 = _T_231 ^ (* src = "crypto_accelerator.v:849" *) _T_275;
  assign _T_315 = _T_263 ^ (* src = "crypto_accelerator.v:850" *) _T_312;
  assign _T_318 = _T_283 ^ (* src = "crypto_accelerator.v:852" *) _T_306;
  assign _T_319 = _T_263 ^ (* src = "crypto_accelerator.v:853" *) _T_318;
  assign _T_321 = _T_273 ^ (* src = "crypto_accelerator.v:854" *) _T_314;
  assign _T_322 = _T_263 ^ (* src = "crypto_accelerator.v:855" *) _T_321;
  assign _T_348 = matrix_0_1[1] ^ (* src = "crypto_accelerator.v:858" *) matrix_0_1[3];
  assign _T_350 = matrix_0_1[4] ^ (* src = "crypto_accelerator.v:859" *) matrix_0_1[7];
  assign _T_352 = matrix_0_1[6] ^ (* src = "crypto_accelerator.v:860" *) matrix_0_1[5];
  assign _T_354 = matrix_0_1[0] ^ (* src = "crypto_accelerator.v:861" *) _T_352;
  assign _T_356 = _T_348 ^ (* src = "crypto_accelerator.v:862" *) _T_350;
  assign _T_358 = matrix_0_1[6] ^ (* src = "crypto_accelerator.v:863" *) matrix_0_1[2];
  assign _T_360 = matrix_0_1[7] ^ (* src = "crypto_accelerator.v:864" *) matrix_0_1[1];
  assign _T_362 = _T_348 ^ (* src = "crypto_accelerator.v:865" *) _T_358;
  assign _T_364 = matrix_0_1[1] ^ (* src = "crypto_accelerator.v:866" *) _T_354;
  assign _T_366 = matrix_0_1[4] ^ (* src = "crypto_accelerator.v:867" *) _T_354;
  assign _T_368 = matrix_0_1[0] ^ (* src = "crypto_accelerator.v:868" *) _T_356;
  assign _T_370 = _T_356 ^ (* src = "crypto_accelerator.v:869" *) _T_358;
  assign _T_372 = matrix_0_1[5] ^ (* src = "crypto_accelerator.v:870" *) matrix_0_1[2];
  assign _T_374 = _T_352 ^ (* src = "crypto_accelerator.v:871" *) _T_356;
  assign _T_376 = matrix_0_1[2] ^ (* src = "crypto_accelerator.v:872" *) _T_360;
  assign _T_378 = matrix_0_1[7] ^ (* src = "crypto_accelerator.v:873" *) matrix_0_1[2];
  assign _T_380 = matrix_0_1[0] ^ (* src = "crypto_accelerator.v:874" *) _T_362;
  assign _T_382 = matrix_0_1[1] ^ (* src = "crypto_accelerator.v:875" *) matrix_0_1[2];
  assign _T_384 = _T_350 ^ (* src = "crypto_accelerator.v:876" *) _T_382;
  assign _T_386 = _T_354 ^ (* src = "crypto_accelerator.v:877" *) _T_376;
  assign _T_388 = _T_348 ^ (* src = "crypto_accelerator.v:878" *) _T_372;
  assign _T_390 = matrix_0_1[7] ^ (* src = "crypto_accelerator.v:879" *) _T_354;
  assign _T_392 = _T_388 ^ (* src = "crypto_accelerator.v:880" *) _T_356;
  assign _T_394 = _T_388 ^ (* src = "crypto_accelerator.v:881" *) _T_360;
  assign _T_396 = _T_360 ^ (* src = "crypto_accelerator.v:882" *) _T_384;
  assign _T_398 = _T_378 ^ (* src = "crypto_accelerator.v:883" *) _T_374;
  assign _T_400 = _T_390 ^ (* src = "crypto_accelerator.v:884" *) _T_380;
  assign _T_406 = _T_370 ^ (* src = "crypto_accelerator.v:887" *) _T_402;
  assign _T_410 = _T_408 ^ (* src = "crypto_accelerator.v:889" *) _T_402;
  assign _T_416 = _T_394 ^ (* src = "crypto_accelerator.v:892" *) _T_412;
  assign _T_420 = _T_418 ^ (* src = "crypto_accelerator.v:894" *) _T_412;
  assign _T_426 = _T_424 ^ (* src = "crypto_accelerator.v:897" *) _T_422;
  assign _T_430 = _T_428 ^ (* src = "crypto_accelerator.v:899" *) _T_422;
  assign _T_432 = _T_406 ^ (* src = "crypto_accelerator.v:900" *) _T_404;
  assign _T_434 = _T_410 ^ (* src = "crypto_accelerator.v:901" *) _T_398;
  assign _T_436 = _T_416 ^ (* src = "crypto_accelerator.v:902" *) _T_414;
  assign _T_438 = _T_420 ^ (* src = "crypto_accelerator.v:903" *) _T_430;
  assign _T_440 = _T_432 ^ (* src = "crypto_accelerator.v:904" *) _T_426;
  assign _T_442 = _T_434 ^ (* src = "crypto_accelerator.v:905" *) _T_430;
  assign _T_444 = _T_436 ^ (* src = "crypto_accelerator.v:906" *) _T_426;
  assign _T_446 = _T_438 ^ (* src = "crypto_accelerator.v:907" *) _T_400;
  assign _T_448 = _T_444 ^ (* src = "crypto_accelerator.v:908" *) _T_446;
  assign _T_452 = _T_442 ^ (* src = "crypto_accelerator.v:910" *) _T_450;
  assign _T_454 = _T_440 ^ (* src = "crypto_accelerator.v:911" *) _T_442;
  assign _T_456 = _T_446 ^ (* src = "crypto_accelerator.v:912" *) _T_450;
  assign _T_466 = _T_454 ^ (* src = "crypto_accelerator.v:917" *) _T_450;
  assign _T_472 = _T_448 ^ (* src = "crypto_accelerator.v:920" *) _T_450;
  assign _T_474 = _T_442 ^ (* src = "crypto_accelerator.v:921" *) _T_458;
  assign _T_476 = _T_464 ^ (* src = "crypto_accelerator.v:922" *) _T_466;
  assign _T_478 = _T_446 ^ (* src = "crypto_accelerator.v:923" *) _T_460;
  assign _T_480 = _T_470 ^ (* src = "crypto_accelerator.v:924" *) _T_472;
  assign _T_482 = _T_476 ^ (* src = "crypto_accelerator.v:925" *) _T_480;
  assign _T_484 = _T_474 ^ (* src = "crypto_accelerator.v:926" *) _T_478;
  assign _T_486 = _T_474 ^ (* src = "crypto_accelerator.v:927" *) _T_476;
  assign _T_488 = _T_478 ^ (* src = "crypto_accelerator.v:928" *) _T_480;
  assign _T_490 = _T_484 ^ (* src = "crypto_accelerator.v:929" *) _T_482;
  assign _T_528 = _T_522 ^ (* src = "crypto_accelerator.v:948" *) _T_524;
  assign _T_530 = _T_500 ^ (* src = "crypto_accelerator.v:949" *) _T_512;
  assign _T_532 = _T_506 ^ (* src = "crypto_accelerator.v:950" *) _T_528;
  assign _T_534 = _T_510 ^ (* src = "crypto_accelerator.v:951" *) _T_530;
  assign _T_536 = _T_496 ^ (* src = "crypto_accelerator.v:952" *) _T_516;
  assign _T_538 = _T_492 ^ (* src = "crypto_accelerator.v:953" *) _T_498;
  assign _T_540 = _T_528 ^ (* src = "crypto_accelerator.v:954" *) _T_538;
  assign _T_542 = _T_494 ^ (* src = "crypto_accelerator.v:955" *) _T_534;
  assign _T_544 = _T_492 ^ (* src = "crypto_accelerator.v:956" *) _T_504;
  assign _T_546 = _T_502 ^ (* src = "crypto_accelerator.v:957" *) _T_518;
  assign _T_548 = _T_508 ^ (* src = "crypto_accelerator.v:958" *) _T_520;
  assign _T_550 = _T_496 ^ (* src = "crypto_accelerator.v:959" *) _T_542;
  assign _T_552 = _T_536 ^ (* src = "crypto_accelerator.v:960" *) _T_548;
  assign _T_554 = _T_514 ^ (* src = "crypto_accelerator.v:961" *) _T_530;
  assign _T_556 = _T_498 ^ (* src = "crypto_accelerator.v:962" *) _T_504;
  assign _T_558 = _T_534 ^ (* src = "crypto_accelerator.v:963" *) _T_556;
  assign _T_560 = _T_526 ^ (* src = "crypto_accelerator.v:964" *) _T_552;
  assign _T_562 = _T_522 ^ (* src = "crypto_accelerator.v:965" *) _T_544;
  assign _T_564 = _T_536 ^ (* src = "crypto_accelerator.v:966" *) _T_546;
  assign _T_565 = _T_532 ^ (* src = "crypto_accelerator.v:967" *) _T_558;
  assign _T_566 = _T_560 ^ (* src = "crypto_accelerator.v:968" *) _T_562;
  assign _T_569 = _T_502 ^ (* src = "crypto_accelerator.v:970" *) _T_528;
  assign _T_570 = _T_540 ^ (* src = "crypto_accelerator.v:971" *) _T_542;
  assign _T_571 = _T_550 ^ (* src = "crypto_accelerator.v:972" *) _T_569;
  assign _T_573 = _T_500 ^ (* src = "crypto_accelerator.v:973" *) _T_516;
  assign _T_575 = _T_538 ^ (* src = "crypto_accelerator.v:974" *) _T_554;
  assign _T_576 = _T_540 ^ (* src = "crypto_accelerator.v:975" *) _T_564;
  assign _T_579 = _T_508 ^ (* src = "crypto_accelerator.v:977" *) _T_546;
  assign _T_581 = _T_573 ^ (* src = "crypto_accelerator.v:978" *) _T_579;
  assign _T_583 = _T_500 ^ (* src = "crypto_accelerator.v:979" *) _T_544;
  assign _T_584 = _T_532 ^ (* src = "crypto_accelerator.v:980" *) _T_581;
  assign _T_587 = _T_552 ^ (* src = "crypto_accelerator.v:982" *) _T_575;
  assign _T_588 = _T_532 ^ (* src = "crypto_accelerator.v:983" *) _T_587;
  assign _T_590 = _T_542 ^ (* src = "crypto_accelerator.v:984" *) _T_583;
  assign _T_591 = _T_532 ^ (* src = "crypto_accelerator.v:985" *) _T_590;
  assign _T_617 = matrix_0_2[1] ^ (* src = "crypto_accelerator.v:988" *) matrix_0_2[3];
  assign _T_619 = matrix_0_2[4] ^ (* src = "crypto_accelerator.v:989" *) matrix_0_2[7];
  assign _T_621 = matrix_0_2[6] ^ (* src = "crypto_accelerator.v:990" *) matrix_0_2[5];
  assign _T_623 = matrix_0_2[0] ^ (* src = "crypto_accelerator.v:991" *) _T_621;
  assign _T_625 = _T_617 ^ (* src = "crypto_accelerator.v:992" *) _T_619;
  assign _T_627 = matrix_0_2[6] ^ (* src = "crypto_accelerator.v:993" *) matrix_0_2[2];
  assign _T_629 = matrix_0_2[7] ^ (* src = "crypto_accelerator.v:994" *) matrix_0_2[1];
  assign _T_631 = _T_617 ^ (* src = "crypto_accelerator.v:995" *) _T_627;
  assign _T_633 = matrix_0_2[1] ^ (* src = "crypto_accelerator.v:996" *) _T_623;
  assign _T_635 = matrix_0_2[4] ^ (* src = "crypto_accelerator.v:997" *) _T_623;
  assign _T_637 = matrix_0_2[0] ^ (* src = "crypto_accelerator.v:998" *) _T_625;
  assign _T_639 = _T_625 ^ (* src = "crypto_accelerator.v:999" *) _T_627;
  (* src = "crypto_accelerator.v:2847" *)
  MixColsModule MixColsModule (
    .io_in_0_0(matrix_0_0),
    .io_in_0_1(matrix_0_1),
    .io_in_0_2(matrix_0_2),
    .io_in_0_3(matrix_0_3),
    .io_in_1_0(matrix_1_0),
    .io_in_1_1(matrix_1_1),
    .io_in_1_2(matrix_1_2),
    .io_in_1_3(matrix_1_3),
    .io_in_2_0(matrix_2_0),
    .io_in_2_1(matrix_2_1),
    .io_in_2_2(matrix_2_2),
    .io_in_2_3(matrix_2_3),
    .io_in_3_0(matrix_3_0),
    .io_in_3_1(matrix_3_1),
    .io_in_3_2(matrix_3_2),
    .io_in_3_3(matrix_3_3),
    .io_out_0_0(MixColsModule_io_out_0_0),
    .io_out_0_1(MixColsModule_io_out_0_1),
    .io_out_0_2(MixColsModule_io_out_0_2),
    .io_out_0_3(MixColsModule_io_out_0_3),
    .io_out_1_0(MixColsModule_io_out_1_0),
    .io_out_1_1(MixColsModule_io_out_1_1),
    .io_out_1_2(MixColsModule_io_out_1_2),
    .io_out_1_3(MixColsModule_io_out_1_3),
    .io_out_2_0(MixColsModule_io_out_2_0),
    .io_out_2_1(MixColsModule_io_out_2_1),
    .io_out_2_2(MixColsModule_io_out_2_2),
    .io_out_2_3(MixColsModule_io_out_2_3),
    .io_out_3_0(MixColsModule_io_out_3_0),
    .io_out_3_1(MixColsModule_io_out_3_1),
    .io_out_3_2(MixColsModule_io_out_3_2),
    .io_out_3_3(MixColsModule_io_out_3_3)
  );
  assign MixColsModule_io_in_0_0 = matrix_0_0;
  assign MixColsModule_io_in_0_1 = matrix_0_1;
  assign MixColsModule_io_in_0_2 = matrix_0_2;
  assign MixColsModule_io_in_0_3 = matrix_0_3;
  assign MixColsModule_io_in_1_0 = matrix_1_0;
  assign MixColsModule_io_in_1_1 = matrix_1_1;
  assign MixColsModule_io_in_1_2 = matrix_1_2;
  assign MixColsModule_io_in_1_3 = matrix_1_3;
  assign MixColsModule_io_in_2_0 = matrix_2_0;
  assign MixColsModule_io_in_2_1 = matrix_2_1;
  assign MixColsModule_io_in_2_2 = matrix_2_2;
  assign MixColsModule_io_in_2_3 = matrix_2_3;
  assign MixColsModule_io_in_3_0 = matrix_3_0;
  assign MixColsModule_io_in_3_1 = matrix_3_1;
  assign MixColsModule_io_in_3_2 = matrix_3_2;
  assign MixColsModule_io_in_3_3 = matrix_3_3;
  assign _T_16 = { matrix_2_0, matrix_2_1, matrix_2_2, matrix_2_3, matrix_3_0, matrix_3_1, matrix_3_2, matrix_3_3 };
  assign _T_23 = { matrix_0_0, matrix_0_1, matrix_0_2, matrix_0_3, matrix_1_0, matrix_1_1, matrix_1_2, matrix_1_3 };
  assign _T_3 = io_outputValid;
  assign _T_32 = { io_keys_0_2_0, io_keys_0_2_1, io_keys_0_2_2, io_keys_0_2_3, io_keys_0_3_0, io_keys_0_3_1, io_keys_0_3_2, io_keys_0_3_3 };
  assign _T_40 = { io_keys_0_0_0, io_keys_0_0_1, io_keys_0_0_2, io_keys_0_0_3, io_keys_0_1_0, io_keys_0_1_1, io_keys_0_1_2, io_keys_0_1_3, io_keys_0_2_0, io_keys_0_2_1, io_keys_0_2_2, io_keys_0_2_3, io_keys_0_3_0, io_keys_0_3_1, io_keys_0_3_2, io_keys_0_3_3 };
  assign initOut_0_0 = _T_41[127:120];
  assign initOut_0_1 = _T_41[119:112];
  assign initOut_0_2 = _T_41[111:104];
  assign initOut_0_3 = _T_41[103:96];
  assign initOut_1_0 = _T_41[95:88];
  assign initOut_1_1 = _T_41[87:80];
  assign initOut_1_2 = _T_41[79:72];
  assign initOut_1_3 = _T_41[71:64];
  assign initOut_2_0 = _T_41[63:56];
  assign initOut_2_1 = _T_41[55:48];
  assign initOut_2_2 = _T_41[47:40];
  assign initOut_2_3 = _T_41[39:32];
  assign initOut_3_0 = _T_41[31:24];
  assign initOut_3_1 = _T_41[23:16];
  assign initOut_3_2 = _T_41[15:8];
  assign initOut_3_3 = _T_41[7:0];
  assign io_dataOut = { matrix_0_0, matrix_0_1, matrix_0_2, matrix_0_3, matrix_1_0, matrix_1_1, matrix_1_2, matrix_1_3, matrix_2_0, matrix_2_1, matrix_2_2, matrix_2_3, matrix_3_0, matrix_3_1, matrix_3_2, matrix_3_3 };
  assign io_ivOut = { matrix_0_0, matrix_0_1, matrix_0_2, matrix_0_3, matrix_1_0, matrix_1_1, matrix_1_2, matrix_1_3, matrix_2_0, matrix_2_1, matrix_2_2, matrix_2_3, matrix_3_0, matrix_3_1, matrix_3_2, matrix_3_3 };
  assign roundPart1_0_0 = { _T_296, _T_323, _T_298, _T_301, _T_302, _T_319, _T_316, _T_308 };
  assign roundPart1_0_1 = { _T_1642, _T_1669, _T_1644, _T_1647, _T_1648, _T_1665, _T_1662, _T_1654 };
  assign roundPart1_0_2 = { _T_2988, _T_3015, _T_2990, _T_2993, _T_2994, _T_3011, _T_3008, _T_3000 };
  assign roundPart1_0_3 = { _T_4334, _T_4361, _T_4336, _T_4339, _T_4340, _T_4357, _T_4354, _T_4346 };
  assign roundPart1_1_0 = { _T_1373, _T_1400, _T_1375, _T_1378, _T_1379, _T_1396, _T_1393, _T_1385 };
  assign roundPart1_1_1 = { _T_2719, _T_2746, _T_2721, _T_2724, _T_2725, _T_2742, _T_2739, _T_2731 };
  assign roundPart1_1_2 = { _T_4065, _T_4092, _T_4067, _T_4070, _T_4071, _T_4088, _T_4085, _T_4077 };
  assign roundPart1_1_3 = { _T_1103, _T_1130, _T_1105, _T_1108, _T_1109, _T_1126, _T_1123, _T_1115 };
  assign roundPart1_2_0 = { _T_2450, _T_2477, _T_2452, _T_2455, _T_2456, _T_2473, _T_2470, _T_2462 };
  assign roundPart1_2_1 = { _T_3796, _T_3823, _T_3798, _T_3801, _T_3802, _T_3819, _T_3816, _T_3808 };
  assign roundPart1_2_2 = { _T_834, _T_861, _T_836, _T_839, _T_840, _T_857, _T_854, _T_846 };
  assign roundPart1_2_3 = { _T_2180, _T_2207, _T_2182, _T_2185, _T_2186, _T_2203, _T_2200, _T_2192 };
  assign roundPart1_3_0 = { _T_3527, _T_3554, _T_3529, _T_3532, _T_3533, _T_3550, _T_3547, _T_3539 };
  assign roundPart1_3_1 = { _T_565, _T_592, _T_567, _T_570, _T_571, _T_588, _T_585, _T_577 };
  assign roundPart1_3_2 = { _T_1911, _T_1938, _T_1913, _T_1916, _T_1917, _T_1934, _T_1931, _T_1923 };
  assign roundPart1_3_3 = { _T_3257, _T_3284, _T_3259, _T_3262, _T_3263, _T_3280, _T_3277, _T_3269 };
endmodule
