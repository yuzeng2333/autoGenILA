module SDP_Y_CORE_cfg_mul_src_rsc_triosy_obj_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:805" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:806" *)
  output outsig;
  assign outsig = in_0;
endmodule
