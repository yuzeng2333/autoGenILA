module \$paramod\SDP_X_mgc_io_sync_v1\valid=0 (ld, lz);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:77" *)
  input ld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:78" *)
  output lz;
  assign lz = ld;
endmodule
