module CDMA_chn_alu_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:358" *)
  input in_0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:359" *)
  output outsig;
  assign outsig = in_0;
endmodule
