module \$paramod\SDP_Y_CVT_mgc_in_wire_v1\rscid=7\width=2 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_cvt.v:78" *)
  output [1:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_cvt.v:79" *)
  input [1:0] z;
  assign d = z;
endmodule
