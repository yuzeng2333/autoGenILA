module FP17_ADD_leading_sign_23_0(mantissa, rtn);
  (* src = "./vmod/vlibs/HLS_fp17_add.v:110" *)
  wire _000_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *)
  wire _001_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:121" *)
  wire _002_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *)
  wire _003_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *)
  wire _004_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:123" *)
  wire _005_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *)
  wire _006_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *)
  wire _007_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _008_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _009_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _010_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _011_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _012_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *)
  wire _013_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _014_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _015_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _016_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _017_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:131" *)
  wire _018_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:131" *)
  wire _019_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:131" *)
  wire _020_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:102" *)
  wire _021_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:109" *)
  wire _022_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *)
  wire _023_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:100" *)
  wire _024_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:104" *)
  wire _025_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:105" *)
  wire _026_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:106" *)
  wire _027_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:111" *)
  wire _028_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:112" *)
  wire _029_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:113" *)
  wire _030_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *)
  wire _031_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _032_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _033_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _034_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *)
  wire _035_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:98" *)
  wire _036_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:99" *)
  wire _037_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:116" *)
  wire _038_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *)
  wire _039_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *)
  wire _040_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *)
  wire _041_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *)
  wire _042_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *)
  wire _043_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *)
  wire _044_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *)
  wire _045_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *)
  wire _046_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _047_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _048_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _049_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _050_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _051_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _052_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _053_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _054_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *)
  wire _055_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *)
  wire _056_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *)
  wire _057_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _058_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _059_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _060_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *)
  wire _061_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *)
  wire _062_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *)
  wire _063_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:120" *)
  wire _064_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *)
  wire _065_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *)
  wire _066_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *)
  wire _067_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _068_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *)
  wire _069_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *)
  wire _070_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *)
  wire _071_;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:96" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:94" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:93" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:95" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:83" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:78" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:84" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:79" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:85" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:80" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:86" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:81" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:87" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:82" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:77" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:92" *)
  wire c_h_1_10;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:88" *)
  wire c_h_1_2;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:89" *)
  wire c_h_1_5;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:90" *)
  wire c_h_1_6;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:91" *)
  wire c_h_1_9;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:74" *)
  input [22:0] mantissa;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:75" *)
  output [4:0] rtn;
  assign c_h_1_2 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp17_add.v:101" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3 = _021_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:103" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp17_add.v:107" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/vlibs/HLS_fp17_add.v:108" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _022_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:110" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:110" *) c_h_1_5;
  assign c_h_1_9 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp17_add.v:114" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  assign c_h_1_10 = c_h_1_6 & (* src = "./vmod/vlibs/HLS_fp17_add.v:115" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl = c_h_1_6 & (* src = "./vmod/vlibs/HLS_fp17_add.v:116" *) _038_;
  assign _001_ = c_h_1_2 & (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *) _062_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl = _001_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *) _063_;
  assign _002_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp17_add.v:121" *) _064_;
  assign _003_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *) _065_;
  assign _004_ = _041_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *) c_h_1_6;
  assign _005_ = _002_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:123" *) _042_;
  assign _006_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *) _066_;
  assign _007_ = _043_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *) c_h_1_10;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl = _005_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *) _044_;
  assign _008_ = _068_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) c_h_1_2;
  assign _009_ = _046_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) _048_;
  assign _010_ = _070_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) c_h_1_5;
  assign _011_ = _050_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) _052_;
  assign _012_ = _053_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) c_h_1_6;
  assign _013_ = _009_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *) _054_;
  assign _014_ = _057_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) c_h_1_9;
  assign _015_ = _056_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) _058_;
  assign _016_ = _059_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) c_h_1_10;
  assign _017_ = _013_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) _060_;
  assign _018_ = _061_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:131" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  assign _019_ = _018_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:131" *) c_h_1_9;
  assign _020_ = _019_ & (* src = "./vmod/vlibs/HLS_fp17_add.v:131" *) c_h_1_10;
  assign _021_ = ! (* src = "./vmod/vlibs/HLS_fp17_add.v:102" *) mantissa[16:15];
  assign _022_ = ! (* src = "./vmod/vlibs/HLS_fp17_add.v:109" *) mantissa[8:7];
  assign _023_ = mantissa[2:1] == (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *) 1'b1;
  assign _024_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:100" *) mantissa[18:17];
  assign _025_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:104" *) mantissa[12:11];
  assign _026_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:105" *) mantissa[14:13];
  assign _027_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:106" *) mantissa[10:9];
  assign _028_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:111" *) mantissa[4:3];
  assign _029_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:112" *) mantissa[6:5];
  assign _030_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:113" *) mantissa[2:1];
  assign _031_ = mantissa[21:20] != (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *) 1'b1;
  assign _032_ = mantissa[17:16] != (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) 1'b1;
  assign _033_ = mantissa[13:12] != (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) 1'b1;
  assign _034_ = mantissa[9:8] != (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) 1'b1;
  assign _035_ = mantissa[5:4] != (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *) 1'b1;
  assign _036_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:98" *) mantissa[20:19];
  assign _037_ = | (* src = "./vmod/vlibs/HLS_fp17_add.v:99" *) mantissa[22:21];
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:100" *) _024_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:104" *) _025_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:105" *) _026_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:106" *) _027_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:111" *) _028_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:112" *) _029_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:113" *) _030_;
  assign _038_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:116" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign _039_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign _040_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *) c_h_1_10;
  assign _041_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *) _003_;
  assign _042_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *) _004_;
  assign _043_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *) _006_;
  assign _044_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *) _007_;
  assign _045_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *) _031_;
  assign _046_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *) _067_;
  assign _047_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) _032_;
  assign _048_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) _008_;
  assign _049_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) _033_;
  assign _050_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) _069_;
  assign _051_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) _034_;
  assign _052_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) _010_;
  assign _053_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) _011_;
  assign _054_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) _012_;
  assign _055_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *) _035_;
  assign _056_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *) _071_;
  assign _057_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *) _023_;
  assign _058_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) _014_;
  assign _059_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) _015_;
  assign _060_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) _016_;
  assign _061_ = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:130" *) mantissa[0];
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:98" *) _036_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp17_add.v:99" *) _037_;
  assign _062_ = c_h_1_5 | (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *) _039_;
  assign _063_ = c_h_1_9 | (* src = "./vmod/vlibs/HLS_fp17_add.v:118" *) _040_;
  assign _064_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp17_add.v:120" *) _036_;
  assign _065_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp17_add.v:122" *) _025_;
  assign _066_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp17_add.v:124" *) _028_;
  assign _067_ = mantissa[22] | (* src = "./vmod/vlibs/HLS_fp17_add.v:126" *) _045_;
  assign _068_ = mantissa[18] | (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) _047_;
  assign _069_ = mantissa[14] | (* src = "./vmod/vlibs/HLS_fp17_add.v:127" *) _049_;
  assign _070_ = mantissa[10] | (* src = "./vmod/vlibs/HLS_fp17_add.v:128" *) _051_;
  assign _071_ = mantissa[6] | (* src = "./vmod/vlibs/HLS_fp17_add.v:129" *) _055_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl = _017_ | (* src = "./vmod/vlibs/HLS_fp17_add.v:131" *) _020_;
  assign rtn = { c_h_1_10, IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl, IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl, IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl, IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl };
endmodule
