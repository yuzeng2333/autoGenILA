module AN2D4PO4(A1, A2, Z);
  (* src = "./vmod/vlibs/AN2D4PO4.v:14" *)
  input A1;
  (* src = "./vmod/vlibs/AN2D4PO4.v:14" *)
  input A2;
  (* src = "./vmod/vlibs/AN2D4PO4.v:15" *)
  output Z;
  assign Z = A1 & (* src = "./vmod/vlibs/AN2D4PO4.v:16" *) A2;
endmodule
