module expand_key_128(clk, in, out_1, out_2, rcon);
  logic [7:0] _0000_;
  logic _0001_;
  logic _0002_;
  logic _0003_;
  logic _0004_;
  logic _0005_;
  logic _0006_;
  logic _0007_;
  logic _0008_;
  logic _0009_;
  logic _0010_;
  logic _0011_;
  logic _0012_;
  logic _0013_;
  logic _0014_;
  logic _0015_;
  logic _0016_;
  logic _0017_;
  logic _0018_;
  logic _0019_;
  logic _0020_;
  logic _0021_;
  logic _0022_;
  logic _0023_;
  logic _0024_;
  logic _0025_;
  logic _0026_;
  logic _0027_;
  logic _0028_;
  logic _0029_;
  logic _0030_;
  logic _0031_;
  logic _0032_;
  logic _0033_;
  logic _0034_;
  logic _0035_;
  logic _0036_;
  logic _0037_;
  logic _0038_;
  logic _0039_;
  logic _0040_;
  logic _0041_;
  logic _0042_;
  logic _0043_;
  logic _0044_;
  logic _0045_;
  logic _0046_;
  logic _0047_;
  logic _0048_;
  logic _0049_;
  logic _0050_;
  logic _0051_;
  logic _0052_;
  logic _0053_;
  logic _0054_;
  logic _0055_;
  logic _0056_;
  logic _0057_;
  logic _0058_;
  logic _0059_;
  logic _0060_;
  logic _0061_;
  logic _0062_;
  logic _0063_;
  logic _0064_;
  logic _0065_;
  logic _0066_;
  logic _0067_;
  logic _0068_;
  logic _0069_;
  logic _0070_;
  logic _0071_;
  logic _0072_;
  logic _0073_;
  logic _0074_;
  logic _0075_;
  logic _0076_;
  logic _0077_;
  logic _0078_;
  logic _0079_;
  logic _0080_;
  logic _0081_;
  logic _0082_;
  logic _0083_;
  logic _0084_;
  logic _0085_;
  logic _0086_;
  logic _0087_;
  logic _0088_;
  logic _0089_;
  logic _0090_;
  logic _0091_;
  logic _0092_;
  logic _0093_;
  logic _0094_;
  logic _0095_;
  logic _0096_;
  logic _0097_;
  logic _0098_;
  logic _0099_;
  logic _0100_;
  logic _0101_;
  logic _0102_;
  logic _0103_;
  logic _0104_;
  logic _0105_;
  logic _0106_;
  logic _0107_;
  logic _0108_;
  logic _0109_;
  logic _0110_;
  logic _0111_;
  logic _0112_;
  logic _0113_;
  logic _0114_;
  logic _0115_;
  logic _0116_;
  logic _0117_;
  logic _0118_;
  logic _0119_;
  logic _0120_;
  logic _0121_;
  logic _0122_;
  logic _0123_;
  logic _0124_;
  logic _0125_;
  logic _0126_;
  logic _0127_;
  logic _0128_;
  logic _0129_;
  logic _0130_;
  logic _0131_;
  logic _0132_;
  logic _0133_;
  logic _0134_;
  logic _0135_;
  logic _0136_;
  logic _0137_;
  logic _0138_;
  logic _0139_;
  logic _0140_;
  logic _0141_;
  logic _0142_;
  logic _0143_;
  logic _0144_;
  logic _0145_;
  logic _0146_;
  logic _0147_;
  logic _0148_;
  logic _0149_;
  logic _0150_;
  logic _0151_;
  logic _0152_;
  logic _0153_;
  logic _0154_;
  logic _0155_;
  logic _0156_;
  logic _0157_;
  logic _0158_;
  logic _0159_;
  logic _0160_;
  logic _0161_;
  logic _0162_;
  logic _0163_;
  logic _0164_;
  logic _0165_;
  logic _0166_;
  logic _0167_;
  logic _0168_;
  logic _0169_;
  logic _0170_;
  logic _0171_;
  logic _0172_;
  logic _0173_;
  logic _0174_;
  logic _0175_;
  logic _0176_;
  logic _0177_;
  logic _0178_;
  logic _0179_;
  logic _0180_;
  logic _0181_;
  logic _0182_;
  logic _0183_;
  logic _0184_;
  logic _0185_;
  logic _0186_;
  logic _0187_;
  logic _0188_;
  logic _0189_;
  logic _0190_;
  logic _0191_;
  logic _0192_;
  logic _0193_;
  logic _0194_;
  logic _0195_;
  logic _0196_;
  logic _0197_;
  logic _0198_;
  logic _0199_;
  logic _0200_;
  logic _0201_;
  logic _0202_;
  logic _0203_;
  logic _0204_;
  logic _0205_;
  logic _0206_;
  logic _0207_;
  logic _0208_;
  logic _0209_;
  logic _0210_;
  logic _0211_;
  logic _0212_;
  logic _0213_;
  logic _0214_;
  logic _0215_;
  logic _0216_;
  logic _0217_;
  logic _0218_;
  logic _0219_;
  logic _0220_;
  logic _0221_;
  logic _0222_;
  logic _0223_;
  logic _0224_;
  logic _0225_;
  logic _0226_;
  logic _0227_;
  logic _0228_;
  logic _0229_;
  logic _0230_;
  logic _0231_;
  logic _0232_;
  logic _0233_;
  logic _0234_;
  logic _0235_;
  logic _0236_;
  logic _0237_;
  logic _0238_;
  logic _0239_;
  logic _0240_;
  logic _0241_;
  logic _0242_;
  logic _0243_;
  logic _0244_;
  logic _0245_;
  logic _0246_;
  logic _0247_;
  logic _0248_;
  logic _0249_;
  logic _0250_;
  logic _0251_;
  logic _0252_;
  logic _0253_;
  logic _0254_;
  logic _0255_;
  logic _0256_;
  logic [7:0] _0257_;
  logic _0258_;
  logic _0259_;
  logic _0260_;
  logic _0261_;
  logic _0262_;
  logic _0263_;
  logic _0264_;
  logic _0265_;
  logic _0266_;
  logic _0267_;
  logic _0268_;
  logic _0269_;
  logic _0270_;
  logic _0271_;
  logic _0272_;
  logic _0273_;
  logic _0274_;
  logic _0275_;
  logic _0276_;
  logic _0277_;
  logic _0278_;
  logic _0279_;
  logic _0280_;
  logic _0281_;
  logic _0282_;
  logic _0283_;
  logic _0284_;
  logic _0285_;
  logic _0286_;
  logic _0287_;
  logic _0288_;
  logic _0289_;
  logic _0290_;
  logic _0291_;
  logic _0292_;
  logic _0293_;
  logic _0294_;
  logic _0295_;
  logic _0296_;
  logic _0297_;
  logic _0298_;
  logic _0299_;
  logic _0300_;
  logic _0301_;
  logic _0302_;
  logic _0303_;
  logic _0304_;
  logic _0305_;
  logic _0306_;
  logic _0307_;
  logic _0308_;
  logic _0309_;
  logic _0310_;
  logic _0311_;
  logic _0312_;
  logic _0313_;
  logic _0314_;
  logic _0315_;
  logic _0316_;
  logic _0317_;
  logic _0318_;
  logic _0319_;
  logic _0320_;
  logic _0321_;
  logic _0322_;
  logic _0323_;
  logic _0324_;
  logic _0325_;
  logic _0326_;
  logic _0327_;
  logic _0328_;
  logic _0329_;
  logic _0330_;
  logic _0331_;
  logic _0332_;
  logic _0333_;
  logic _0334_;
  logic _0335_;
  logic _0336_;
  logic _0337_;
  logic _0338_;
  logic _0339_;
  logic _0340_;
  logic _0341_;
  logic _0342_;
  logic _0343_;
  logic _0344_;
  logic _0345_;
  logic _0346_;
  logic _0347_;
  logic _0348_;
  logic _0349_;
  logic _0350_;
  logic _0351_;
  logic _0352_;
  logic _0353_;
  logic _0354_;
  logic _0355_;
  logic _0356_;
  logic _0357_;
  logic _0358_;
  logic _0359_;
  logic _0360_;
  logic _0361_;
  logic _0362_;
  logic _0363_;
  logic _0364_;
  logic _0365_;
  logic _0366_;
  logic _0367_;
  logic _0368_;
  logic _0369_;
  logic _0370_;
  logic _0371_;
  logic _0372_;
  logic _0373_;
  logic _0374_;
  logic _0375_;
  logic _0376_;
  logic _0377_;
  logic _0378_;
  logic _0379_;
  logic _0380_;
  logic _0381_;
  logic _0382_;
  logic _0383_;
  logic _0384_;
  logic _0385_;
  logic _0386_;
  logic _0387_;
  logic _0388_;
  logic _0389_;
  logic _0390_;
  logic _0391_;
  logic _0392_;
  logic _0393_;
  logic _0394_;
  logic _0395_;
  logic _0396_;
  logic _0397_;
  logic _0398_;
  logic _0399_;
  logic _0400_;
  logic _0401_;
  logic _0402_;
  logic _0403_;
  logic _0404_;
  logic _0405_;
  logic _0406_;
  logic _0407_;
  logic _0408_;
  logic _0409_;
  logic _0410_;
  logic _0411_;
  logic _0412_;
  logic _0413_;
  logic _0414_;
  logic _0415_;
  logic _0416_;
  logic _0417_;
  logic _0418_;
  logic _0419_;
  logic _0420_;
  logic _0421_;
  logic _0422_;
  logic _0423_;
  logic _0424_;
  logic _0425_;
  logic _0426_;
  logic _0427_;
  logic _0428_;
  logic _0429_;
  logic _0430_;
  logic _0431_;
  logic _0432_;
  logic _0433_;
  logic _0434_;
  logic _0435_;
  logic _0436_;
  logic _0437_;
  logic _0438_;
  logic _0439_;
  logic _0440_;
  logic _0441_;
  logic _0442_;
  logic _0443_;
  logic _0444_;
  logic _0445_;
  logic _0446_;
  logic _0447_;
  logic _0448_;
  logic _0449_;
  logic _0450_;
  logic _0451_;
  logic _0452_;
  logic _0453_;
  logic _0454_;
  logic _0455_;
  logic _0456_;
  logic _0457_;
  logic _0458_;
  logic _0459_;
  logic _0460_;
  logic _0461_;
  logic _0462_;
  logic _0463_;
  logic _0464_;
  logic _0465_;
  logic _0466_;
  logic _0467_;
  logic _0468_;
  logic _0469_;
  logic _0470_;
  logic _0471_;
  logic _0472_;
  logic _0473_;
  logic _0474_;
  logic _0475_;
  logic _0476_;
  logic _0477_;
  logic _0478_;
  logic _0479_;
  logic _0480_;
  logic _0481_;
  logic _0482_;
  logic _0483_;
  logic _0484_;
  logic _0485_;
  logic _0486_;
  logic _0487_;
  logic _0488_;
  logic _0489_;
  logic _0490_;
  logic _0491_;
  logic _0492_;
  logic _0493_;
  logic _0494_;
  logic _0495_;
  logic _0496_;
  logic _0497_;
  logic _0498_;
  logic _0499_;
  logic _0500_;
  logic _0501_;
  logic _0502_;
  logic _0503_;
  logic _0504_;
  logic _0505_;
  logic _0506_;
  logic _0507_;
  logic _0508_;
  logic _0509_;
  logic _0510_;
  logic _0511_;
  logic _0512_;
  logic _0513_;
  logic [7:0] _0514_;
  logic _0515_;
  logic _0516_;
  logic _0517_;
  logic _0518_;
  logic _0519_;
  logic _0520_;
  logic _0521_;
  logic _0522_;
  logic _0523_;
  logic _0524_;
  logic _0525_;
  logic _0526_;
  logic _0527_;
  logic _0528_;
  logic _0529_;
  logic _0530_;
  logic _0531_;
  logic _0532_;
  logic _0533_;
  logic _0534_;
  logic _0535_;
  logic _0536_;
  logic _0537_;
  logic _0538_;
  logic _0539_;
  logic _0540_;
  logic _0541_;
  logic _0542_;
  logic _0543_;
  logic _0544_;
  logic _0545_;
  logic _0546_;
  logic _0547_;
  logic _0548_;
  logic _0549_;
  logic _0550_;
  logic _0551_;
  logic _0552_;
  logic _0553_;
  logic _0554_;
  logic _0555_;
  logic _0556_;
  logic _0557_;
  logic _0558_;
  logic _0559_;
  logic _0560_;
  logic _0561_;
  logic _0562_;
  logic _0563_;
  logic _0564_;
  logic _0565_;
  logic _0566_;
  logic _0567_;
  logic _0568_;
  logic _0569_;
  logic _0570_;
  logic _0571_;
  logic _0572_;
  logic _0573_;
  logic _0574_;
  logic _0575_;
  logic _0576_;
  logic _0577_;
  logic _0578_;
  logic _0579_;
  logic _0580_;
  logic _0581_;
  logic _0582_;
  logic _0583_;
  logic _0584_;
  logic _0585_;
  logic _0586_;
  logic _0587_;
  logic _0588_;
  logic _0589_;
  logic _0590_;
  logic _0591_;
  logic _0592_;
  logic _0593_;
  logic _0594_;
  logic _0595_;
  logic _0596_;
  logic _0597_;
  logic _0598_;
  logic _0599_;
  logic _0600_;
  logic _0601_;
  logic _0602_;
  logic _0603_;
  logic _0604_;
  logic _0605_;
  logic _0606_;
  logic _0607_;
  logic _0608_;
  logic _0609_;
  logic _0610_;
  logic _0611_;
  logic _0612_;
  logic _0613_;
  logic _0614_;
  logic _0615_;
  logic _0616_;
  logic _0617_;
  logic _0618_;
  logic _0619_;
  logic _0620_;
  logic _0621_;
  logic _0622_;
  logic _0623_;
  logic _0624_;
  logic _0625_;
  logic _0626_;
  logic _0627_;
  logic _0628_;
  logic _0629_;
  logic _0630_;
  logic _0631_;
  logic _0632_;
  logic _0633_;
  logic _0634_;
  logic _0635_;
  logic _0636_;
  logic _0637_;
  logic _0638_;
  logic _0639_;
  logic _0640_;
  logic _0641_;
  logic _0642_;
  logic _0643_;
  logic _0644_;
  logic _0645_;
  logic _0646_;
  logic _0647_;
  logic _0648_;
  logic _0649_;
  logic _0650_;
  logic _0651_;
  logic _0652_;
  logic _0653_;
  logic _0654_;
  logic _0655_;
  logic _0656_;
  logic _0657_;
  logic _0658_;
  logic _0659_;
  logic _0660_;
  logic _0661_;
  logic _0662_;
  logic _0663_;
  logic _0664_;
  logic _0665_;
  logic _0666_;
  logic _0667_;
  logic _0668_;
  logic _0669_;
  logic _0670_;
  logic _0671_;
  logic _0672_;
  logic _0673_;
  logic _0674_;
  logic _0675_;
  logic _0676_;
  logic _0677_;
  logic _0678_;
  logic _0679_;
  logic _0680_;
  logic _0681_;
  logic _0682_;
  logic _0683_;
  logic _0684_;
  logic _0685_;
  logic _0686_;
  logic _0687_;
  logic _0688_;
  logic _0689_;
  logic _0690_;
  logic _0691_;
  logic _0692_;
  logic _0693_;
  logic _0694_;
  logic _0695_;
  logic _0696_;
  logic _0697_;
  logic _0698_;
  logic _0699_;
  logic _0700_;
  logic _0701_;
  logic _0702_;
  logic _0703_;
  logic _0704_;
  logic _0705_;
  logic _0706_;
  logic _0707_;
  logic _0708_;
  logic _0709_;
  logic _0710_;
  logic _0711_;
  logic _0712_;
  logic _0713_;
  logic _0714_;
  logic _0715_;
  logic _0716_;
  logic _0717_;
  logic _0718_;
  logic _0719_;
  logic _0720_;
  logic _0721_;
  logic _0722_;
  logic _0723_;
  logic _0724_;
  logic _0725_;
  logic _0726_;
  logic _0727_;
  logic _0728_;
  logic _0729_;
  logic _0730_;
  logic _0731_;
  logic _0732_;
  logic _0733_;
  logic _0734_;
  logic _0735_;
  logic _0736_;
  logic _0737_;
  logic _0738_;
  logic _0739_;
  logic _0740_;
  logic _0741_;
  logic _0742_;
  logic _0743_;
  logic _0744_;
  logic _0745_;
  logic _0746_;
  logic _0747_;
  logic _0748_;
  logic _0749_;
  logic _0750_;
  logic _0751_;
  logic _0752_;
  logic _0753_;
  logic _0754_;
  logic _0755_;
  logic _0756_;
  logic _0757_;
  logic _0758_;
  logic _0759_;
  logic _0760_;
  logic _0761_;
  logic _0762_;
  logic _0763_;
  logic _0764_;
  logic _0765_;
  logic _0766_;
  logic _0767_;
  logic _0768_;
  logic _0769_;
  logic _0770_;
  logic [7:0] _0771_;
  logic _0772_;
  logic _0773_;
  logic _0774_;
  logic _0775_;
  logic _0776_;
  logic _0777_;
  logic _0778_;
  logic _0779_;
  logic _0780_;
  logic _0781_;
  logic _0782_;
  logic _0783_;
  logic _0784_;
  logic _0785_;
  logic _0786_;
  logic _0787_;
  logic _0788_;
  logic _0789_;
  logic _0790_;
  logic _0791_;
  logic _0792_;
  logic _0793_;
  logic _0794_;
  logic _0795_;
  logic _0796_;
  logic _0797_;
  logic _0798_;
  logic _0799_;
  logic _0800_;
  logic _0801_;
  logic _0802_;
  logic _0803_;
  logic _0804_;
  logic _0805_;
  logic _0806_;
  logic _0807_;
  logic _0808_;
  logic _0809_;
  logic _0810_;
  logic _0811_;
  logic _0812_;
  logic _0813_;
  logic _0814_;
  logic _0815_;
  logic _0816_;
  logic _0817_;
  logic _0818_;
  logic _0819_;
  logic _0820_;
  logic _0821_;
  logic _0822_;
  logic _0823_;
  logic _0824_;
  logic _0825_;
  logic _0826_;
  logic _0827_;
  logic _0828_;
  logic _0829_;
  logic _0830_;
  logic _0831_;
  logic _0832_;
  logic _0833_;
  logic _0834_;
  logic _0835_;
  logic _0836_;
  logic _0837_;
  logic _0838_;
  logic _0839_;
  logic _0840_;
  logic _0841_;
  logic _0842_;
  logic _0843_;
  logic _0844_;
  logic _0845_;
  logic _0846_;
  logic _0847_;
  logic _0848_;
  logic _0849_;
  logic _0850_;
  logic _0851_;
  logic _0852_;
  logic _0853_;
  logic _0854_;
  logic _0855_;
  logic _0856_;
  logic _0857_;
  logic _0858_;
  logic _0859_;
  logic _0860_;
  logic _0861_;
  logic _0862_;
  logic _0863_;
  logic _0864_;
  logic _0865_;
  logic _0866_;
  logic _0867_;
  logic _0868_;
  logic _0869_;
  logic _0870_;
  logic _0871_;
  logic _0872_;
  logic _0873_;
  logic _0874_;
  logic _0875_;
  logic _0876_;
  logic _0877_;
  logic _0878_;
  logic _0879_;
  logic _0880_;
  logic _0881_;
  logic _0882_;
  logic _0883_;
  logic _0884_;
  logic _0885_;
  logic _0886_;
  logic _0887_;
  logic _0888_;
  logic _0889_;
  logic _0890_;
  logic _0891_;
  logic _0892_;
  logic _0893_;
  logic _0894_;
  logic _0895_;
  logic _0896_;
  logic _0897_;
  logic _0898_;
  logic _0899_;
  logic _0900_;
  logic _0901_;
  logic _0902_;
  logic _0903_;
  logic _0904_;
  logic _0905_;
  logic _0906_;
  logic _0907_;
  logic _0908_;
  logic _0909_;
  logic _0910_;
  logic _0911_;
  logic _0912_;
  logic _0913_;
  logic _0914_;
  logic _0915_;
  logic _0916_;
  logic _0917_;
  logic _0918_;
  logic _0919_;
  logic _0920_;
  logic _0921_;
  logic _0922_;
  logic _0923_;
  logic _0924_;
  logic _0925_;
  logic _0926_;
  logic _0927_;
  logic _0928_;
  logic _0929_;
  logic _0930_;
  logic _0931_;
  logic _0932_;
  logic _0933_;
  logic _0934_;
  logic _0935_;
  logic _0936_;
  logic _0937_;
  logic _0938_;
  logic _0939_;
  logic _0940_;
  logic _0941_;
  logic _0942_;
  logic _0943_;
  logic _0944_;
  logic _0945_;
  logic _0946_;
  logic _0947_;
  logic _0948_;
  logic _0949_;
  logic _0950_;
  logic _0951_;
  logic _0952_;
  logic _0953_;
  logic _0954_;
  logic _0955_;
  logic _0956_;
  logic _0957_;
  logic _0958_;
  logic _0959_;
  logic _0960_;
  logic _0961_;
  logic _0962_;
  logic _0963_;
  logic _0964_;
  logic _0965_;
  logic _0966_;
  logic _0967_;
  logic _0968_;
  logic _0969_;
  logic _0970_;
  logic _0971_;
  logic _0972_;
  logic _0973_;
  logic _0974_;
  logic _0975_;
  logic _0976_;
  logic _0977_;
  logic _0978_;
  logic _0979_;
  logic _0980_;
  logic _0981_;
  logic _0982_;
  logic _0983_;
  logic _0984_;
  logic _0985_;
  logic _0986_;
  logic _0987_;
  logic _0988_;
  logic _0989_;
  logic _0990_;
  logic _0991_;
  logic _0992_;
  logic _0993_;
  logic _0994_;
  logic _0995_;
  logic _0996_;
  logic _0997_;
  logic _0998_;
  logic _0999_;
  logic _1000_;
  logic _1001_;
  logic _1002_;
  logic _1003_;
  logic _1004_;
  logic _1005_;
  logic _1006_;
  logic _1007_;
  logic _1008_;
  logic _1009_;
  logic _1010_;
  logic _1011_;
  logic _1012_;
  logic _1013_;
  logic _1014_;
  logic _1015_;
  logic _1016_;
  logic _1017_;
  logic _1018_;
  logic _1019_;
  logic _1020_;
  logic _1021_;
  logic _1022_;
  logic _1023_;
  logic _1024_;
  logic _1025_;
  logic _1026_;
  logic _1027_;
  logic \S4_0.S_0.clk ;
  logic [7:0] \S4_0.S_0.in ;
  logic [7:0] \S4_0.S_0.out ;
  logic \S4_0.S_1.clk ;
  logic [7:0] \S4_0.S_1.in ;
  logic [7:0] \S4_0.S_1.out ;
  logic \S4_0.S_2.clk ;
  logic [7:0] \S4_0.S_2.in ;
  logic [7:0] \S4_0.S_2.out ;
  logic \S4_0.S_3.clk ;
  logic [7:0] \S4_0.S_3.in ;
  logic [7:0] \S4_0.S_3.out ;
  logic \S4_0.clk ;
  logic [31:0] \S4_0.in ;
  logic [31:0] \S4_0.out ;
  input clk;
  input [127:0] in;
  logic [31:0] k0;
  logic [31:0] k0a;
  logic [31:0] k0b;
  logic [31:0] k1;
  logic [31:0] k1a;
  logic [31:0] k1b;
  logic [31:0] k2;
  logic [31:0] k2a;
  logic [31:0] k2b;
  logic [31:0] k3;
  logic [31:0] k3a;
  logic [31:0] k3b;
  logic [31:0] k4a;
  output [127:0] out_1;
  logic [127:0] out_1;
  output [127:0] out_2;
  input [7:0] rcon;
  logic [31:0] v0;
  logic [31:0] v1;
  logic [31:0] v2;
  logic [31:0] v3;

  logic [127:0] fangyuan0;
  assign fangyuan0 = { k0b, k1b, k2b, k3b };
  always @(posedge clk)
      out_1 <= fangyuan0;

  logic [31:0] fangyuan1;
  assign fangyuan1 = { v0[31:24], in[119:96] };
  always @(posedge clk)
      k0a <= fangyuan1;
  always @(posedge clk)
      k1a <= v1;
  always @(posedge clk)
      k2a <= v2;
  always @(posedge clk)
      k3a <= v3;
  always @(posedge clk)
      \S4_0.S_0.out <= _0000_;
  assign _0001_ = in[23:16] == 8'ha8;
  assign _0002_ = in[23:16] == 8'ha7;
  assign _0003_ = in[23:16] == 8'ha6;
  assign _0004_ = in[23:16] == 8'ha5;
  assign _0005_ = in[23:16] == 8'ha4;
  assign _0006_ = in[23:16] == 8'ha3;
  assign _0007_ = in[23:16] == 8'ha2;
  assign _0008_ = in[23:16] == 8'ha1;
  assign _0009_ = in[23:16] == 8'ha0;
  assign _0010_ = in[23:16] == 8'h9f;
  assign _0011_ = in[23:16] == 8'h9e;
  assign _0012_ = in[23:16] == 8'h9d;
  assign _0013_ = in[23:16] == 8'h9c;
  assign _0014_ = in[23:16] == 8'h9b;
  assign _0015_ = in[23:16] == 8'h9a;
  assign _0016_ = in[23:16] == 8'h99;
  assign _0017_ = in[23:16] == 8'h98;
  assign _0018_ = in[23:16] == 8'h97;
  assign _0019_ = in[23:16] == 8'h96;
  assign _0020_ = in[23:16] == 8'h95;
  logic [255:0] fangyuan2;
  assign fangyuan2 = { _0182_, _0181_, _0180_, _0179_, _0178_, _0177_, _0176_, _0175_, _0174_, _0172_, _0171_, _0170_, _0169_, _0168_, _0167_, _0166_, _0165_, _0164_, _0163_, _0161_, _0160_, _0159_, _0158_, _0157_, _0156_, _0155_, _0154_, _0153_, _0152_, _0150_, _0149_, _0148_, _0147_, _0146_, _0145_, _0144_, _0143_, _0142_, _0141_, _0139_, _0138_, _0137_, _0136_, _0135_, _0134_, _0133_, _0132_, _0131_, _0130_, _0128_, _0127_, _0126_, _0125_, _0124_, _0123_, _0122_, _0121_, _0120_, _0119_, _0117_, _0116_, _0115_, _0114_, _0113_, _0112_, _0111_, _0110_, _0109_, _0108_, _0106_, _0105_, _0104_, _0103_, _0102_, _0101_, _0100_, _0099_, _0098_, _0097_, _0095_, _0094_, _0093_, _0092_, _0091_, _0090_, _0089_, _0088_, _0087_, _0086_, _0084_, _0083_, _0082_, _0081_, _0080_, _0079_, _0078_, _0077_, _0076_, _0075_, _0073_, _0072_, _0071_, _0070_, _0069_, _0068_, _0067_, _0066_, _0065_, _0064_, _0062_, _0061_, _0060_, _0059_, _0058_, _0057_, _0056_, _0055_, _0054_, _0053_, _0051_, _0050_, _0049_, _0048_, _0047_, _0046_, _0045_, _0044_, _0043_, _0042_, _0040_, _0039_, _0038_, _0037_, _0036_, _0035_, _0034_, _0033_, _0032_, _0031_, _0030_, _0029_, _0028_, _0027_, _0026_, _0025_, _0024_, _0023_, _0022_, _0021_, _0020_, _0019_, _0018_, _0017_, _0016_, _0015_, _0014_, _0013_, _0012_, _0011_, _0010_, _0009_, _0008_, _0007_, _0006_, _0005_, _0004_, _0003_, _0002_, _0001_, _0256_, _0255_, _0254_, _0253_, _0252_, _0251_, _0250_, _0249_, _0248_, _0247_, _0246_, _0245_, _0244_, _0243_, _0242_, _0241_, _0240_, _0239_, _0238_, _0237_, _0236_, _0235_, _0234_, _0233_, _0232_, _0231_, _0230_, _0229_, _0228_, _0227_, _0226_, _0225_, _0224_, _0223_, _0222_, _0221_, _0220_, _0219_, _0218_, _0217_, _0216_, _0215_, _0214_, _0213_, _0212_, _0211_, _0210_, _0209_, _0208_, _0207_, _0206_, _0205_, _0204_, _0203_, _0202_, _0201_, _0200_, _0199_, _0198_, _0197_, _0196_, _0195_, _0194_, _0193_, _0192_, _0191_, _0190_, _0189_, _0188_, _0187_, _0186_, _0185_, _0184_, _0183_, _0173_, _0162_, _0151_, _0140_, _0129_, _0118_, _0107_, _0096_, _0085_, _0074_, _0063_, _0052_, _0041_ };

  always @(\S4_0.S_0.out or fangyuan2) begin
    casez (fangyuan2)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0000_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0000_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0000_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0000_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0000_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0000_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0000_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0000_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0000_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0000_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0000_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0000_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0000_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0000_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0000_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0000_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0000_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0000_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0000_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0000_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0000_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0000_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0000_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0000_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0000_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0000_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0000_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0000_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0000_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0000_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0000_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0000_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0000_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0000_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0000_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0000_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0000_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0000_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0000_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0000_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0000_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0000_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0000_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0000_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0000_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0000_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0000_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0000_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0000_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0000_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0000_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0000_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0000_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0000_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0000_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0000_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0000_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100011 ;
      default:
        _0000_ = \S4_0.S_0.out ;
    endcase
  end
  assign _0021_ = in[23:16] == 8'h94;
  assign _0022_ = in[23:16] == 8'h93;
  assign _0023_ = in[23:16] == 8'h92;
  assign _0024_ = in[23:16] == 8'h91;
  assign _0025_ = in[23:16] == 8'h90;
  assign _0026_ = in[23:16] == 8'h8f;
  assign _0027_ = in[23:16] == 8'h8e;
  assign _0028_ = in[23:16] == 8'h8d;
  assign _0029_ = in[23:16] == 8'h8c;
  assign _0030_ = in[23:16] == 8'h8b;
  assign _0031_ = in[23:16] == 8'h8a;
  assign _0032_ = in[23:16] == 8'h89;
  assign _0033_ = in[23:16] == 8'h88;
  assign _0034_ = in[23:16] == 8'h87;
  assign _0035_ = in[23:16] == 8'h86;
  assign _0036_ = in[23:16] == 8'h85;
  assign _0037_ = in[23:16] == 8'h84;
  assign _0038_ = in[23:16] == 8'h83;
  assign _0039_ = in[23:16] == 8'h82;
  assign _0040_ = in[23:16] == 8'h81;
  assign _0041_ = in[23:16] == 8'hff;
  assign _0042_ = in[23:16] == 8'h80;
  assign _0043_ = in[23:16] == 7'h7f;
  assign _0044_ = in[23:16] == 7'h7e;
  assign _0045_ = in[23:16] == 7'h7d;
  assign _0046_ = in[23:16] == 7'h7c;
  assign _0047_ = in[23:16] == 7'h7b;
  assign _0048_ = in[23:16] == 7'h7a;
  assign _0049_ = in[23:16] == 7'h79;
  assign _0050_ = in[23:16] == 7'h78;
  assign _0051_ = in[23:16] == 7'h77;
  assign _0052_ = in[23:16] == 8'hfe;
  assign _0053_ = in[23:16] == 7'h76;
  assign _0054_ = in[23:16] == 7'h75;
  assign _0055_ = in[23:16] == 7'h74;
  assign _0056_ = in[23:16] == 7'h73;
  assign _0057_ = in[23:16] == 7'h72;
  assign _0058_ = in[23:16] == 7'h71;
  assign _0059_ = in[23:16] == 7'h70;
  assign _0060_ = in[23:16] == 7'h6f;
  assign _0061_ = in[23:16] == 7'h6e;
  assign _0062_ = in[23:16] == 7'h6d;
  assign _0063_ = in[23:16] == 8'hfd;
  assign _0064_ = in[23:16] == 7'h6c;
  assign _0065_ = in[23:16] == 7'h6b;
  assign _0066_ = in[23:16] == 7'h6a;
  assign _0067_ = in[23:16] == 7'h69;
  assign _0068_ = in[23:16] == 7'h68;
  assign _0069_ = in[23:16] == 7'h67;
  assign _0070_ = in[23:16] == 7'h66;
  assign _0071_ = in[23:16] == 7'h65;
  assign _0072_ = in[23:16] == 7'h64;
  assign _0073_ = in[23:16] == 7'h63;
  assign _0074_ = in[23:16] == 8'hfc;
  assign _0075_ = in[23:16] == 7'h62;
  assign _0076_ = in[23:16] == 7'h61;
  assign _0077_ = in[23:16] == 7'h60;
  assign _0078_ = in[23:16] == 7'h5f;
  assign _0079_ = in[23:16] == 7'h5e;
  assign _0080_ = in[23:16] == 7'h5d;
  assign _0081_ = in[23:16] == 7'h5c;
  assign _0082_ = in[23:16] == 7'h5b;
  assign _0083_ = in[23:16] == 7'h5a;
  assign _0084_ = in[23:16] == 7'h59;
  assign _0085_ = in[23:16] == 8'hfb;
  assign _0086_ = in[23:16] == 7'h58;
  assign _0087_ = in[23:16] == 7'h57;
  assign _0088_ = in[23:16] == 7'h56;
  assign _0089_ = in[23:16] == 7'h55;
  assign _0090_ = in[23:16] == 7'h54;
  assign _0091_ = in[23:16] == 7'h53;
  assign _0092_ = in[23:16] == 7'h52;
  assign _0093_ = in[23:16] == 7'h51;
  assign _0094_ = in[23:16] == 7'h50;
  assign _0095_ = in[23:16] == 7'h4f;
  assign _0096_ = in[23:16] == 8'hfa;
  assign _0097_ = in[23:16] == 7'h4e;
  assign _0098_ = in[23:16] == 7'h4d;
  assign _0099_ = in[23:16] == 7'h4c;
  assign _0100_ = in[23:16] == 7'h4b;
  assign _0101_ = in[23:16] == 7'h4a;
  assign _0102_ = in[23:16] == 7'h49;
  assign _0103_ = in[23:16] == 7'h48;
  assign _0104_ = in[23:16] == 7'h47;
  assign _0105_ = in[23:16] == 7'h46;
  assign _0106_ = in[23:16] == 7'h45;
  assign _0107_ = in[23:16] == 8'hf9;
  assign _0108_ = in[23:16] == 7'h44;
  assign _0109_ = in[23:16] == 7'h43;
  assign _0110_ = in[23:16] == 7'h42;
  assign _0111_ = in[23:16] == 7'h41;
  assign _0112_ = in[23:16] == 7'h40;
  assign _0113_ = in[23:16] == 6'h3f;
  assign _0114_ = in[23:16] == 6'h3e;
  assign _0115_ = in[23:16] == 6'h3d;
  assign _0116_ = in[23:16] == 6'h3c;
  assign _0117_ = in[23:16] == 6'h3b;
  assign _0118_ = in[23:16] == 8'hf8;
  assign _0119_ = in[23:16] == 6'h3a;
  assign _0120_ = in[23:16] == 6'h39;
  assign _0121_ = in[23:16] == 6'h38;
  assign _0122_ = in[23:16] == 6'h37;
  assign _0123_ = in[23:16] == 6'h36;
  assign _0124_ = in[23:16] == 6'h35;
  assign _0125_ = in[23:16] == 6'h34;
  assign _0126_ = in[23:16] == 6'h33;
  assign _0127_ = in[23:16] == 6'h32;
  assign _0128_ = in[23:16] == 6'h31;
  assign _0129_ = in[23:16] == 8'hf7;
  assign _0130_ = in[23:16] == 6'h30;
  assign _0131_ = in[23:16] == 6'h2f;
  assign _0132_ = in[23:16] == 6'h2e;
  assign _0133_ = in[23:16] == 6'h2d;
  assign _0134_ = in[23:16] == 6'h2c;
  assign _0135_ = in[23:16] == 6'h2b;
  assign _0136_ = in[23:16] == 6'h2a;
  assign _0137_ = in[23:16] == 6'h29;
  assign _0138_ = in[23:16] == 6'h28;
  assign _0139_ = in[23:16] == 6'h27;
  assign _0140_ = in[23:16] == 8'hf6;
  assign _0141_ = in[23:16] == 6'h26;
  assign _0142_ = in[23:16] == 6'h25;
  assign _0143_ = in[23:16] == 6'h24;
  assign _0144_ = in[23:16] == 6'h23;
  assign _0145_ = in[23:16] == 6'h22;
  assign _0146_ = in[23:16] == 6'h21;
  assign _0147_ = in[23:16] == 6'h20;
  assign _0148_ = in[23:16] == 5'h1f;
  assign _0149_ = in[23:16] == 5'h1e;
  assign _0150_ = in[23:16] == 5'h1d;
  assign _0151_ = in[23:16] == 8'hf5;
  assign _0152_ = in[23:16] == 5'h1c;
  assign _0153_ = in[23:16] == 5'h1b;
  assign _0154_ = in[23:16] == 5'h1a;
  assign _0155_ = in[23:16] == 5'h19;
  assign _0156_ = in[23:16] == 5'h18;
  assign _0157_ = in[23:16] == 5'h17;
  assign _0158_ = in[23:16] == 5'h16;
  assign _0159_ = in[23:16] == 5'h15;
  assign _0160_ = in[23:16] == 5'h14;
  assign _0161_ = in[23:16] == 5'h13;
  assign _0162_ = in[23:16] == 8'hf4;
  assign _0163_ = in[23:16] == 5'h12;
  assign _0164_ = in[23:16] == 5'h11;
  assign _0165_ = in[23:16] == 5'h10;
  assign _0166_ = in[23:16] == 4'hf;
  assign _0167_ = in[23:16] == 4'he;
  assign _0168_ = in[23:16] == 4'hd;
  assign _0169_ = in[23:16] == 4'hc;
  assign _0170_ = in[23:16] == 4'hb;
  assign _0171_ = in[23:16] == 4'ha;
  assign _0172_ = in[23:16] == 4'h9;
  assign _0173_ = in[23:16] == 8'hf3;
  assign _0174_ = in[23:16] == 4'h8;
  assign _0175_ = in[23:16] == 3'h7;
  assign _0176_ = in[23:16] == 3'h6;
  assign _0177_ = in[23:16] == 3'h5;
  assign _0178_ = in[23:16] == 3'h4;
  assign _0179_ = in[23:16] == 2'h3;
  assign _0180_ = in[23:16] == 2'h2;
  assign _0181_ = in[23:16] == 1'h1;
  assign _0182_ = ! in[23:16];
  assign _0183_ = in[23:16] == 8'hf2;
  assign _0184_ = in[23:16] == 8'hf1;
  assign _0185_ = in[23:16] == 8'hf0;
  assign _0186_ = in[23:16] == 8'hef;
  assign _0187_ = in[23:16] == 8'hee;
  assign _0188_ = in[23:16] == 8'hed;
  assign _0189_ = in[23:16] == 8'hec;
  assign _0190_ = in[23:16] == 8'heb;
  assign _0191_ = in[23:16] == 8'hea;
  assign _0192_ = in[23:16] == 8'he9;
  assign _0193_ = in[23:16] == 8'he8;
  assign _0194_ = in[23:16] == 8'he7;
  assign _0195_ = in[23:16] == 8'he6;
  assign _0196_ = in[23:16] == 8'he5;
  assign _0197_ = in[23:16] == 8'he4;
  assign _0198_ = in[23:16] == 8'he3;
  assign _0199_ = in[23:16] == 8'he2;
  assign _0200_ = in[23:16] == 8'he1;
  assign _0201_ = in[23:16] == 8'he0;
  assign _0202_ = in[23:16] == 8'hdf;
  assign _0203_ = in[23:16] == 8'hde;
  assign _0204_ = in[23:16] == 8'hdd;
  assign _0205_ = in[23:16] == 8'hdc;
  assign _0206_ = in[23:16] == 8'hdb;
  assign _0207_ = in[23:16] == 8'hda;
  assign _0208_ = in[23:16] == 8'hd9;
  assign _0209_ = in[23:16] == 8'hd8;
  assign _0210_ = in[23:16] == 8'hd7;
  assign _0211_ = in[23:16] == 8'hd6;
  assign _0212_ = in[23:16] == 8'hd5;
  assign _0213_ = in[23:16] == 8'hd4;
  assign _0214_ = in[23:16] == 8'hd3;
  assign _0215_ = in[23:16] == 8'hd2;
  assign _0216_ = in[23:16] == 8'hd1;
  assign _0217_ = in[23:16] == 8'hd0;
  assign _0218_ = in[23:16] == 8'hcf;
  assign _0219_ = in[23:16] == 8'hce;
  assign _0220_ = in[23:16] == 8'hcd;
  assign _0221_ = in[23:16] == 8'hcc;
  assign _0222_ = in[23:16] == 8'hcb;
  assign _0223_ = in[23:16] == 8'hca;
  assign _0224_ = in[23:16] == 8'hc9;
  assign _0225_ = in[23:16] == 8'hc8;
  assign _0226_ = in[23:16] == 8'hc7;
  assign _0227_ = in[23:16] == 8'hc6;
  assign _0228_ = in[23:16] == 8'hc5;
  assign _0229_ = in[23:16] == 8'hc4;
  assign _0230_ = in[23:16] == 8'hc3;
  assign _0231_ = in[23:16] == 8'hc2;
  assign _0232_ = in[23:16] == 8'hc1;
  assign _0233_ = in[23:16] == 8'hc0;
  assign _0234_ = in[23:16] == 8'hbf;
  assign _0235_ = in[23:16] == 8'hbe;
  assign _0236_ = in[23:16] == 8'hbd;
  assign _0237_ = in[23:16] == 8'hbc;
  assign _0238_ = in[23:16] == 8'hbb;
  assign _0239_ = in[23:16] == 8'hba;
  assign _0240_ = in[23:16] == 8'hb9;
  assign _0241_ = in[23:16] == 8'hb8;
  assign _0242_ = in[23:16] == 8'hb7;
  assign _0243_ = in[23:16] == 8'hb6;
  assign _0244_ = in[23:16] == 8'hb5;
  assign _0245_ = in[23:16] == 8'hb4;
  assign _0246_ = in[23:16] == 8'hb3;
  assign _0247_ = in[23:16] == 8'hb2;
  assign _0248_ = in[23:16] == 8'hb1;
  assign _0249_ = in[23:16] == 8'hb0;
  assign _0250_ = in[23:16] == 8'haf;
  assign _0251_ = in[23:16] == 8'hae;
  assign _0252_ = in[23:16] == 8'had;
  assign _0253_ = in[23:16] == 8'hac;
  assign _0254_ = in[23:16] == 8'hab;
  assign _0255_ = in[23:16] == 8'haa;
  assign _0256_ = in[23:16] == 8'ha9;
  always @(posedge clk)
      \S4_0.S_1.out <= _0257_;
  assign _0258_ = in[15:8] == 8'ha8;
  assign _0259_ = in[15:8] == 8'ha7;
  assign _0260_ = in[15:8] == 8'ha6;
  assign _0261_ = in[15:8] == 8'ha5;
  assign _0262_ = in[15:8] == 8'ha4;
  assign _0263_ = in[15:8] == 8'ha3;
  assign _0264_ = in[15:8] == 8'ha2;
  assign _0265_ = in[15:8] == 8'ha1;
  assign _0266_ = in[15:8] == 8'ha0;
  assign _0267_ = in[15:8] == 8'h9f;
  assign _0268_ = in[15:8] == 8'h9e;
  assign _0269_ = in[15:8] == 8'h9d;
  assign _0270_ = in[15:8] == 8'h9c;
  assign _0271_ = in[15:8] == 8'h9b;
  assign _0272_ = in[15:8] == 8'h9a;
  assign _0273_ = in[15:8] == 8'h99;
  assign _0274_ = in[15:8] == 8'h98;
  assign _0275_ = in[15:8] == 8'h97;
  assign _0276_ = in[15:8] == 8'h96;
  assign _0277_ = in[15:8] == 8'h95;
  logic [255:0] fangyuan3;
  assign fangyuan3 = { _0439_, _0438_, _0437_, _0436_, _0435_, _0434_, _0433_, _0432_, _0431_, _0429_, _0428_, _0427_, _0426_, _0425_, _0424_, _0423_, _0422_, _0421_, _0420_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0341_, _0340_, _0339_, _0338_, _0337_, _0336_, _0335_, _0334_, _0333_, _0332_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, _0321_, _0319_, _0318_, _0317_, _0316_, _0315_, _0314_, _0313_, _0312_, _0311_, _0310_, _0308_, _0307_, _0306_, _0305_, _0304_, _0303_, _0302_, _0301_, _0300_, _0299_, _0297_, _0296_, _0295_, _0294_, _0293_, _0292_, _0291_, _0290_, _0289_, _0288_, _0287_, _0286_, _0285_, _0284_, _0283_, _0282_, _0281_, _0280_, _0279_, _0278_, _0277_, _0276_, _0275_, _0274_, _0273_, _0272_, _0271_, _0270_, _0269_, _0268_, _0267_, _0266_, _0265_, _0264_, _0263_, _0262_, _0261_, _0260_, _0259_, _0258_, _0513_, _0512_, _0511_, _0510_, _0509_, _0508_, _0507_, _0506_, _0505_, _0504_, _0503_, _0502_, _0501_, _0500_, _0499_, _0498_, _0497_, _0496_, _0495_, _0494_, _0493_, _0492_, _0491_, _0490_, _0489_, _0488_, _0487_, _0486_, _0485_, _0484_, _0483_, _0482_, _0481_, _0480_, _0479_, _0478_, _0477_, _0476_, _0475_, _0474_, _0473_, _0472_, _0471_, _0470_, _0469_, _0468_, _0467_, _0466_, _0465_, _0464_, _0463_, _0462_, _0461_, _0460_, _0459_, _0458_, _0457_, _0456_, _0455_, _0454_, _0453_, _0452_, _0451_, _0450_, _0449_, _0448_, _0447_, _0446_, _0445_, _0444_, _0443_, _0442_, _0441_, _0440_, _0430_, _0419_, _0408_, _0397_, _0386_, _0375_, _0364_, _0353_, _0342_, _0331_, _0320_, _0309_, _0298_ };

  always @(\S4_0.S_1.out or fangyuan3) begin
    casez (fangyuan3)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0257_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0257_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0257_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0257_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0257_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0257_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0257_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0257_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0257_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0257_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0257_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0257_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0257_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0257_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0257_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0257_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0257_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0257_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0257_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0257_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0257_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0257_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0257_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0257_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0257_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0257_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0257_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0257_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0257_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0257_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0257_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0257_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0257_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0257_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0257_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0257_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0257_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0257_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0257_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0257_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0257_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0257_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0257_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0257_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0257_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0257_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0257_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0257_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0257_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0257_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0257_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0257_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0257_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0257_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0257_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0257_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0257_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100011 ;
      default:
        _0257_ = \S4_0.S_1.out ;
    endcase
  end
  assign _0278_ = in[15:8] == 8'h94;
  assign _0279_ = in[15:8] == 8'h93;
  assign _0280_ = in[15:8] == 8'h92;
  assign _0281_ = in[15:8] == 8'h91;
  assign _0282_ = in[15:8] == 8'h90;
  assign _0283_ = in[15:8] == 8'h8f;
  assign _0284_ = in[15:8] == 8'h8e;
  assign _0285_ = in[15:8] == 8'h8d;
  assign _0286_ = in[15:8] == 8'h8c;
  assign _0287_ = in[15:8] == 8'h8b;
  assign _0288_ = in[15:8] == 8'h8a;
  assign _0289_ = in[15:8] == 8'h89;
  assign _0290_ = in[15:8] == 8'h88;
  assign _0291_ = in[15:8] == 8'h87;
  assign _0292_ = in[15:8] == 8'h86;
  assign _0293_ = in[15:8] == 8'h85;
  assign _0294_ = in[15:8] == 8'h84;
  assign _0295_ = in[15:8] == 8'h83;
  assign _0296_ = in[15:8] == 8'h82;
  assign _0297_ = in[15:8] == 8'h81;
  assign _0298_ = in[15:8] == 8'hff;
  assign _0299_ = in[15:8] == 8'h80;
  assign _0300_ = in[15:8] == 7'h7f;
  assign _0301_ = in[15:8] == 7'h7e;
  assign _0302_ = in[15:8] == 7'h7d;
  assign _0303_ = in[15:8] == 7'h7c;
  assign _0304_ = in[15:8] == 7'h7b;
  assign _0305_ = in[15:8] == 7'h7a;
  assign _0306_ = in[15:8] == 7'h79;
  assign _0307_ = in[15:8] == 7'h78;
  assign _0308_ = in[15:8] == 7'h77;
  assign _0309_ = in[15:8] == 8'hfe;
  assign _0310_ = in[15:8] == 7'h76;
  assign _0311_ = in[15:8] == 7'h75;
  assign _0312_ = in[15:8] == 7'h74;
  assign _0313_ = in[15:8] == 7'h73;
  assign _0314_ = in[15:8] == 7'h72;
  assign _0315_ = in[15:8] == 7'h71;
  assign _0316_ = in[15:8] == 7'h70;
  assign _0317_ = in[15:8] == 7'h6f;
  assign _0318_ = in[15:8] == 7'h6e;
  assign _0319_ = in[15:8] == 7'h6d;
  assign _0320_ = in[15:8] == 8'hfd;
  assign _0321_ = in[15:8] == 7'h6c;
  assign _0322_ = in[15:8] == 7'h6b;
  assign _0323_ = in[15:8] == 7'h6a;
  assign _0324_ = in[15:8] == 7'h69;
  assign _0325_ = in[15:8] == 7'h68;
  assign _0326_ = in[15:8] == 7'h67;
  assign _0327_ = in[15:8] == 7'h66;
  assign _0328_ = in[15:8] == 7'h65;
  assign _0329_ = in[15:8] == 7'h64;
  assign _0330_ = in[15:8] == 7'h63;
  assign _0331_ = in[15:8] == 8'hfc;
  assign _0332_ = in[15:8] == 7'h62;
  assign _0333_ = in[15:8] == 7'h61;
  assign _0334_ = in[15:8] == 7'h60;
  assign _0335_ = in[15:8] == 7'h5f;
  assign _0336_ = in[15:8] == 7'h5e;
  assign _0337_ = in[15:8] == 7'h5d;
  assign _0338_ = in[15:8] == 7'h5c;
  assign _0339_ = in[15:8] == 7'h5b;
  assign _0340_ = in[15:8] == 7'h5a;
  assign _0341_ = in[15:8] == 7'h59;
  assign _0342_ = in[15:8] == 8'hfb;
  assign _0343_ = in[15:8] == 7'h58;
  assign _0344_ = in[15:8] == 7'h57;
  assign _0345_ = in[15:8] == 7'h56;
  assign _0346_ = in[15:8] == 7'h55;
  assign _0347_ = in[15:8] == 7'h54;
  assign _0348_ = in[15:8] == 7'h53;
  assign _0349_ = in[15:8] == 7'h52;
  assign _0350_ = in[15:8] == 7'h51;
  assign _0351_ = in[15:8] == 7'h50;
  assign _0352_ = in[15:8] == 7'h4f;
  assign _0353_ = in[15:8] == 8'hfa;
  assign _0354_ = in[15:8] == 7'h4e;
  assign _0355_ = in[15:8] == 7'h4d;
  assign _0356_ = in[15:8] == 7'h4c;
  assign _0357_ = in[15:8] == 7'h4b;
  assign _0358_ = in[15:8] == 7'h4a;
  assign _0359_ = in[15:8] == 7'h49;
  assign _0360_ = in[15:8] == 7'h48;
  assign _0361_ = in[15:8] == 7'h47;
  assign _0362_ = in[15:8] == 7'h46;
  assign _0363_ = in[15:8] == 7'h45;
  assign _0364_ = in[15:8] == 8'hf9;
  assign _0365_ = in[15:8] == 7'h44;
  assign _0366_ = in[15:8] == 7'h43;
  assign _0367_ = in[15:8] == 7'h42;
  assign _0368_ = in[15:8] == 7'h41;
  assign _0369_ = in[15:8] == 7'h40;
  assign _0370_ = in[15:8] == 6'h3f;
  assign _0371_ = in[15:8] == 6'h3e;
  assign _0372_ = in[15:8] == 6'h3d;
  assign _0373_ = in[15:8] == 6'h3c;
  assign _0374_ = in[15:8] == 6'h3b;
  assign _0375_ = in[15:8] == 8'hf8;
  assign _0376_ = in[15:8] == 6'h3a;
  assign _0377_ = in[15:8] == 6'h39;
  assign _0378_ = in[15:8] == 6'h38;
  assign _0379_ = in[15:8] == 6'h37;
  assign _0380_ = in[15:8] == 6'h36;
  assign _0381_ = in[15:8] == 6'h35;
  assign _0382_ = in[15:8] == 6'h34;
  assign _0383_ = in[15:8] == 6'h33;
  assign _0384_ = in[15:8] == 6'h32;
  assign _0385_ = in[15:8] == 6'h31;
  assign _0386_ = in[15:8] == 8'hf7;
  assign _0387_ = in[15:8] == 6'h30;
  assign _0388_ = in[15:8] == 6'h2f;
  assign _0389_ = in[15:8] == 6'h2e;
  assign _0390_ = in[15:8] == 6'h2d;
  assign _0391_ = in[15:8] == 6'h2c;
  assign _0392_ = in[15:8] == 6'h2b;
  assign _0393_ = in[15:8] == 6'h2a;
  assign _0394_ = in[15:8] == 6'h29;
  assign _0395_ = in[15:8] == 6'h28;
  assign _0396_ = in[15:8] == 6'h27;
  assign _0397_ = in[15:8] == 8'hf6;
  assign _0398_ = in[15:8] == 6'h26;
  assign _0399_ = in[15:8] == 6'h25;
  assign _0400_ = in[15:8] == 6'h24;
  assign _0401_ = in[15:8] == 6'h23;
  assign _0402_ = in[15:8] == 6'h22;
  assign _0403_ = in[15:8] == 6'h21;
  assign _0404_ = in[15:8] == 6'h20;
  assign _0405_ = in[15:8] == 5'h1f;
  assign _0406_ = in[15:8] == 5'h1e;
  assign _0407_ = in[15:8] == 5'h1d;
  assign _0408_ = in[15:8] == 8'hf5;
  assign _0409_ = in[15:8] == 5'h1c;
  assign _0410_ = in[15:8] == 5'h1b;
  assign _0411_ = in[15:8] == 5'h1a;
  assign _0412_ = in[15:8] == 5'h19;
  assign _0413_ = in[15:8] == 5'h18;
  assign _0414_ = in[15:8] == 5'h17;
  assign _0415_ = in[15:8] == 5'h16;
  assign _0416_ = in[15:8] == 5'h15;
  assign _0417_ = in[15:8] == 5'h14;
  assign _0418_ = in[15:8] == 5'h13;
  assign _0419_ = in[15:8] == 8'hf4;
  assign _0420_ = in[15:8] == 5'h12;
  assign _0421_ = in[15:8] == 5'h11;
  assign _0422_ = in[15:8] == 5'h10;
  assign _0423_ = in[15:8] == 4'hf;
  assign _0424_ = in[15:8] == 4'he;
  assign _0425_ = in[15:8] == 4'hd;
  assign _0426_ = in[15:8] == 4'hc;
  assign _0427_ = in[15:8] == 4'hb;
  assign _0428_ = in[15:8] == 4'ha;
  assign _0429_ = in[15:8] == 4'h9;
  assign _0430_ = in[15:8] == 8'hf3;
  assign _0431_ = in[15:8] == 4'h8;
  assign _0432_ = in[15:8] == 3'h7;
  assign _0433_ = in[15:8] == 3'h6;
  assign _0434_ = in[15:8] == 3'h5;
  assign _0435_ = in[15:8] == 3'h4;
  assign _0436_ = in[15:8] == 2'h3;
  assign _0437_ = in[15:8] == 2'h2;
  assign _0438_ = in[15:8] == 1'h1;
  assign _0439_ = ! in[15:8];
  assign _0440_ = in[15:8] == 8'hf2;
  assign _0441_ = in[15:8] == 8'hf1;
  assign _0442_ = in[15:8] == 8'hf0;
  assign _0443_ = in[15:8] == 8'hef;
  assign _0444_ = in[15:8] == 8'hee;
  assign _0445_ = in[15:8] == 8'hed;
  assign _0446_ = in[15:8] == 8'hec;
  assign _0447_ = in[15:8] == 8'heb;
  assign _0448_ = in[15:8] == 8'hea;
  assign _0449_ = in[15:8] == 8'he9;
  assign _0450_ = in[15:8] == 8'he8;
  assign _0451_ = in[15:8] == 8'he7;
  assign _0452_ = in[15:8] == 8'he6;
  assign _0453_ = in[15:8] == 8'he5;
  assign _0454_ = in[15:8] == 8'he4;
  assign _0455_ = in[15:8] == 8'he3;
  assign _0456_ = in[15:8] == 8'he2;
  assign _0457_ = in[15:8] == 8'he1;
  assign _0458_ = in[15:8] == 8'he0;
  assign _0459_ = in[15:8] == 8'hdf;
  assign _0460_ = in[15:8] == 8'hde;
  assign _0461_ = in[15:8] == 8'hdd;
  assign _0462_ = in[15:8] == 8'hdc;
  assign _0463_ = in[15:8] == 8'hdb;
  assign _0464_ = in[15:8] == 8'hda;
  assign _0465_ = in[15:8] == 8'hd9;
  assign _0466_ = in[15:8] == 8'hd8;
  assign _0467_ = in[15:8] == 8'hd7;
  assign _0468_ = in[15:8] == 8'hd6;
  assign _0469_ = in[15:8] == 8'hd5;
  assign _0470_ = in[15:8] == 8'hd4;
  assign _0471_ = in[15:8] == 8'hd3;
  assign _0472_ = in[15:8] == 8'hd2;
  assign _0473_ = in[15:8] == 8'hd1;
  assign _0474_ = in[15:8] == 8'hd0;
  assign _0475_ = in[15:8] == 8'hcf;
  assign _0476_ = in[15:8] == 8'hce;
  assign _0477_ = in[15:8] == 8'hcd;
  assign _0478_ = in[15:8] == 8'hcc;
  assign _0479_ = in[15:8] == 8'hcb;
  assign _0480_ = in[15:8] == 8'hca;
  assign _0481_ = in[15:8] == 8'hc9;
  assign _0482_ = in[15:8] == 8'hc8;
  assign _0483_ = in[15:8] == 8'hc7;
  assign _0484_ = in[15:8] == 8'hc6;
  assign _0485_ = in[15:8] == 8'hc5;
  assign _0486_ = in[15:8] == 8'hc4;
  assign _0487_ = in[15:8] == 8'hc3;
  assign _0488_ = in[15:8] == 8'hc2;
  assign _0489_ = in[15:8] == 8'hc1;
  assign _0490_ = in[15:8] == 8'hc0;
  assign _0491_ = in[15:8] == 8'hbf;
  assign _0492_ = in[15:8] == 8'hbe;
  assign _0493_ = in[15:8] == 8'hbd;
  assign _0494_ = in[15:8] == 8'hbc;
  assign _0495_ = in[15:8] == 8'hbb;
  assign _0496_ = in[15:8] == 8'hba;
  assign _0497_ = in[15:8] == 8'hb9;
  assign _0498_ = in[15:8] == 8'hb8;
  assign _0499_ = in[15:8] == 8'hb7;
  assign _0500_ = in[15:8] == 8'hb6;
  assign _0501_ = in[15:8] == 8'hb5;
  assign _0502_ = in[15:8] == 8'hb4;
  assign _0503_ = in[15:8] == 8'hb3;
  assign _0504_ = in[15:8] == 8'hb2;
  assign _0505_ = in[15:8] == 8'hb1;
  assign _0506_ = in[15:8] == 8'hb0;
  assign _0507_ = in[15:8] == 8'haf;
  assign _0508_ = in[15:8] == 8'hae;
  assign _0509_ = in[15:8] == 8'had;
  assign _0510_ = in[15:8] == 8'hac;
  assign _0511_ = in[15:8] == 8'hab;
  assign _0512_ = in[15:8] == 8'haa;
  assign _0513_ = in[15:8] == 8'ha9;
  always @(posedge clk)
      \S4_0.S_2.out <= _0514_;
  assign _0515_ = in[7:0] == 8'ha8;
  assign _0516_ = in[7:0] == 8'ha7;
  assign _0517_ = in[7:0] == 8'ha6;
  assign _0518_ = in[7:0] == 8'ha5;
  assign _0519_ = in[7:0] == 8'ha4;
  assign _0520_ = in[7:0] == 8'ha3;
  assign _0521_ = in[7:0] == 8'ha2;
  assign _0522_ = in[7:0] == 8'ha1;
  assign _0523_ = in[7:0] == 8'ha0;
  assign _0524_ = in[7:0] == 8'h9f;
  assign _0525_ = in[7:0] == 8'h9e;
  assign _0526_ = in[7:0] == 8'h9d;
  assign _0527_ = in[7:0] == 8'h9c;
  assign _0528_ = in[7:0] == 8'h9b;
  assign _0529_ = in[7:0] == 8'h9a;
  assign _0530_ = in[7:0] == 8'h99;
  assign _0531_ = in[7:0] == 8'h98;
  assign _0532_ = in[7:0] == 8'h97;
  assign _0533_ = in[7:0] == 8'h96;
  assign _0534_ = in[7:0] == 8'h95;
  logic [255:0] fangyuan4;
  assign fangyuan4 = { _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0686_, _0685_, _0684_, _0683_, _0682_, _0681_, _0680_, _0679_, _0678_, _0677_, _0675_, _0674_, _0673_, _0672_, _0671_, _0670_, _0669_, _0668_, _0667_, _0666_, _0664_, _0663_, _0662_, _0661_, _0660_, _0659_, _0658_, _0657_, _0656_, _0655_, _0653_, _0652_, _0651_, _0650_, _0649_, _0648_, _0647_, _0646_, _0645_, _0644_, _0642_, _0641_, _0640_, _0639_, _0638_, _0637_, _0636_, _0635_, _0634_, _0633_, _0631_, _0630_, _0629_, _0628_, _0627_, _0626_, _0625_, _0624_, _0623_, _0622_, _0620_, _0619_, _0618_, _0617_, _0616_, _0615_, _0614_, _0613_, _0612_, _0611_, _0609_, _0608_, _0607_, _0606_, _0605_, _0604_, _0603_, _0602_, _0601_, _0600_, _0598_, _0597_, _0596_, _0595_, _0594_, _0593_, _0592_, _0591_, _0590_, _0589_, _0587_, _0586_, _0585_, _0584_, _0583_, _0582_, _0581_, _0580_, _0579_, _0578_, _0576_, _0575_, _0574_, _0573_, _0572_, _0571_, _0570_, _0569_, _0568_, _0567_, _0565_, _0564_, _0563_, _0562_, _0561_, _0560_, _0559_, _0558_, _0557_, _0556_, _0554_, _0553_, _0552_, _0551_, _0550_, _0549_, _0548_, _0547_, _0546_, _0545_, _0544_, _0543_, _0542_, _0541_, _0540_, _0539_, _0538_, _0537_, _0536_, _0535_, _0534_, _0533_, _0532_, _0531_, _0530_, _0529_, _0528_, _0527_, _0526_, _0525_, _0524_, _0523_, _0522_, _0521_, _0520_, _0519_, _0518_, _0517_, _0516_, _0515_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0687_, _0676_, _0665_, _0654_, _0643_, _0632_, _0621_, _0610_, _0599_, _0588_, _0577_, _0566_, _0555_ };

  always @(\S4_0.S_2.out or fangyuan4) begin
    casez (fangyuan4)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0514_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0514_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0514_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0514_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0514_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0514_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0514_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0514_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0514_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0514_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0514_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0514_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0514_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0514_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0514_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0514_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0514_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0514_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0514_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0514_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0514_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0514_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0514_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0514_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0514_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0514_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0514_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0514_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0514_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0514_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0514_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0514_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0514_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0514_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0514_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0514_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0514_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0514_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0514_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0514_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0514_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0514_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0514_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0514_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0514_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0514_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0514_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0514_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0514_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0514_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0514_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0514_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0514_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0514_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0514_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0514_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0514_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0514_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0514_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0514_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0514_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0514_ = 8'b01100011 ;
      default:
        _0514_ = \S4_0.S_2.out ;
    endcase
  end
  assign _0535_ = in[7:0] == 8'h94;
  assign _0536_ = in[7:0] == 8'h93;
  assign _0537_ = in[7:0] == 8'h92;
  assign _0538_ = in[7:0] == 8'h91;
  assign _0539_ = in[7:0] == 8'h90;
  assign _0540_ = in[7:0] == 8'h8f;
  assign _0541_ = in[7:0] == 8'h8e;
  assign _0542_ = in[7:0] == 8'h8d;
  assign _0543_ = in[7:0] == 8'h8c;
  assign _0544_ = in[7:0] == 8'h8b;
  assign _0545_ = in[7:0] == 8'h8a;
  assign _0546_ = in[7:0] == 8'h89;
  assign _0547_ = in[7:0] == 8'h88;
  assign _0548_ = in[7:0] == 8'h87;
  assign _0549_ = in[7:0] == 8'h86;
  assign _0550_ = in[7:0] == 8'h85;
  assign _0551_ = in[7:0] == 8'h84;
  assign _0552_ = in[7:0] == 8'h83;
  assign _0553_ = in[7:0] == 8'h82;
  assign _0554_ = in[7:0] == 8'h81;
  assign _0555_ = in[7:0] == 8'hff;
  assign _0556_ = in[7:0] == 8'h80;
  assign _0557_ = in[7:0] == 7'h7f;
  assign _0558_ = in[7:0] == 7'h7e;
  assign _0559_ = in[7:0] == 7'h7d;
  assign _0560_ = in[7:0] == 7'h7c;
  assign _0561_ = in[7:0] == 7'h7b;
  assign _0562_ = in[7:0] == 7'h7a;
  assign _0563_ = in[7:0] == 7'h79;
  assign _0564_ = in[7:0] == 7'h78;
  assign _0565_ = in[7:0] == 7'h77;
  assign _0566_ = in[7:0] == 8'hfe;
  assign _0567_ = in[7:0] == 7'h76;
  assign _0568_ = in[7:0] == 7'h75;
  assign _0569_ = in[7:0] == 7'h74;
  assign _0570_ = in[7:0] == 7'h73;
  assign _0571_ = in[7:0] == 7'h72;
  assign _0572_ = in[7:0] == 7'h71;
  assign _0573_ = in[7:0] == 7'h70;
  assign _0574_ = in[7:0] == 7'h6f;
  assign _0575_ = in[7:0] == 7'h6e;
  assign _0576_ = in[7:0] == 7'h6d;
  assign _0577_ = in[7:0] == 8'hfd;
  assign _0578_ = in[7:0] == 7'h6c;
  assign _0579_ = in[7:0] == 7'h6b;
  assign _0580_ = in[7:0] == 7'h6a;
  assign _0581_ = in[7:0] == 7'h69;
  assign _0582_ = in[7:0] == 7'h68;
  assign _0583_ = in[7:0] == 7'h67;
  assign _0584_ = in[7:0] == 7'h66;
  assign _0585_ = in[7:0] == 7'h65;
  assign _0586_ = in[7:0] == 7'h64;
  assign _0587_ = in[7:0] == 7'h63;
  assign _0588_ = in[7:0] == 8'hfc;
  assign _0589_ = in[7:0] == 7'h62;
  assign _0590_ = in[7:0] == 7'h61;
  assign _0591_ = in[7:0] == 7'h60;
  assign _0592_ = in[7:0] == 7'h5f;
  assign _0593_ = in[7:0] == 7'h5e;
  assign _0594_ = in[7:0] == 7'h5d;
  assign _0595_ = in[7:0] == 7'h5c;
  assign _0596_ = in[7:0] == 7'h5b;
  assign _0597_ = in[7:0] == 7'h5a;
  assign _0598_ = in[7:0] == 7'h59;
  assign _0599_ = in[7:0] == 8'hfb;
  assign _0600_ = in[7:0] == 7'h58;
  assign _0601_ = in[7:0] == 7'h57;
  assign _0602_ = in[7:0] == 7'h56;
  assign _0603_ = in[7:0] == 7'h55;
  assign _0604_ = in[7:0] == 7'h54;
  assign _0605_ = in[7:0] == 7'h53;
  assign _0606_ = in[7:0] == 7'h52;
  assign _0607_ = in[7:0] == 7'h51;
  assign _0608_ = in[7:0] == 7'h50;
  assign _0609_ = in[7:0] == 7'h4f;
  assign _0610_ = in[7:0] == 8'hfa;
  assign _0611_ = in[7:0] == 7'h4e;
  assign _0612_ = in[7:0] == 7'h4d;
  assign _0613_ = in[7:0] == 7'h4c;
  assign _0614_ = in[7:0] == 7'h4b;
  assign _0615_ = in[7:0] == 7'h4a;
  assign _0616_ = in[7:0] == 7'h49;
  assign _0617_ = in[7:0] == 7'h48;
  assign _0618_ = in[7:0] == 7'h47;
  assign _0619_ = in[7:0] == 7'h46;
  assign _0620_ = in[7:0] == 7'h45;
  assign _0621_ = in[7:0] == 8'hf9;
  assign _0622_ = in[7:0] == 7'h44;
  assign _0623_ = in[7:0] == 7'h43;
  assign _0624_ = in[7:0] == 7'h42;
  assign _0625_ = in[7:0] == 7'h41;
  assign _0626_ = in[7:0] == 7'h40;
  assign _0627_ = in[7:0] == 6'h3f;
  assign _0628_ = in[7:0] == 6'h3e;
  assign _0629_ = in[7:0] == 6'h3d;
  assign _0630_ = in[7:0] == 6'h3c;
  assign _0631_ = in[7:0] == 6'h3b;
  assign _0632_ = in[7:0] == 8'hf8;
  assign _0633_ = in[7:0] == 6'h3a;
  assign _0634_ = in[7:0] == 6'h39;
  assign _0635_ = in[7:0] == 6'h38;
  assign _0636_ = in[7:0] == 6'h37;
  assign _0637_ = in[7:0] == 6'h36;
  assign _0638_ = in[7:0] == 6'h35;
  assign _0639_ = in[7:0] == 6'h34;
  assign _0640_ = in[7:0] == 6'h33;
  assign _0641_ = in[7:0] == 6'h32;
  assign _0642_ = in[7:0] == 6'h31;
  assign _0643_ = in[7:0] == 8'hf7;
  assign _0644_ = in[7:0] == 6'h30;
  assign _0645_ = in[7:0] == 6'h2f;
  assign _0646_ = in[7:0] == 6'h2e;
  assign _0647_ = in[7:0] == 6'h2d;
  assign _0648_ = in[7:0] == 6'h2c;
  assign _0649_ = in[7:0] == 6'h2b;
  assign _0650_ = in[7:0] == 6'h2a;
  assign _0651_ = in[7:0] == 6'h29;
  assign _0652_ = in[7:0] == 6'h28;
  assign _0653_ = in[7:0] == 6'h27;
  assign _0654_ = in[7:0] == 8'hf6;
  assign _0655_ = in[7:0] == 6'h26;
  assign _0656_ = in[7:0] == 6'h25;
  assign _0657_ = in[7:0] == 6'h24;
  assign _0658_ = in[7:0] == 6'h23;
  assign _0659_ = in[7:0] == 6'h22;
  assign _0660_ = in[7:0] == 6'h21;
  assign _0661_ = in[7:0] == 6'h20;
  assign _0662_ = in[7:0] == 5'h1f;
  assign _0663_ = in[7:0] == 5'h1e;
  assign _0664_ = in[7:0] == 5'h1d;
  assign _0665_ = in[7:0] == 8'hf5;
  assign _0666_ = in[7:0] == 5'h1c;
  assign _0667_ = in[7:0] == 5'h1b;
  assign _0668_ = in[7:0] == 5'h1a;
  assign _0669_ = in[7:0] == 5'h19;
  assign _0670_ = in[7:0] == 5'h18;
  assign _0671_ = in[7:0] == 5'h17;
  assign _0672_ = in[7:0] == 5'h16;
  assign _0673_ = in[7:0] == 5'h15;
  assign _0674_ = in[7:0] == 5'h14;
  assign _0675_ = in[7:0] == 5'h13;
  assign _0676_ = in[7:0] == 8'hf4;
  assign _0677_ = in[7:0] == 5'h12;
  assign _0678_ = in[7:0] == 5'h11;
  assign _0679_ = in[7:0] == 5'h10;
  assign _0680_ = in[7:0] == 4'hf;
  assign _0681_ = in[7:0] == 4'he;
  assign _0682_ = in[7:0] == 4'hd;
  assign _0683_ = in[7:0] == 4'hc;
  assign _0684_ = in[7:0] == 4'hb;
  assign _0685_ = in[7:0] == 4'ha;
  assign _0686_ = in[7:0] == 4'h9;
  assign _0687_ = in[7:0] == 8'hf3;
  assign _0688_ = in[7:0] == 4'h8;
  assign _0689_ = in[7:0] == 3'h7;
  assign _0690_ = in[7:0] == 3'h6;
  assign _0691_ = in[7:0] == 3'h5;
  assign _0692_ = in[7:0] == 3'h4;
  assign _0693_ = in[7:0] == 2'h3;
  assign _0694_ = in[7:0] == 2'h2;
  assign _0695_ = in[7:0] == 1'h1;
  assign _0696_ = ! in[7:0];
  assign _0697_ = in[7:0] == 8'hf2;
  assign _0698_ = in[7:0] == 8'hf1;
  assign _0699_ = in[7:0] == 8'hf0;
  assign _0700_ = in[7:0] == 8'hef;
  assign _0701_ = in[7:0] == 8'hee;
  assign _0702_ = in[7:0] == 8'hed;
  assign _0703_ = in[7:0] == 8'hec;
  assign _0704_ = in[7:0] == 8'heb;
  assign _0705_ = in[7:0] == 8'hea;
  assign _0706_ = in[7:0] == 8'he9;
  assign _0707_ = in[7:0] == 8'he8;
  assign _0708_ = in[7:0] == 8'he7;
  assign _0709_ = in[7:0] == 8'he6;
  assign _0710_ = in[7:0] == 8'he5;
  assign _0711_ = in[7:0] == 8'he4;
  assign _0712_ = in[7:0] == 8'he3;
  assign _0713_ = in[7:0] == 8'he2;
  assign _0714_ = in[7:0] == 8'he1;
  assign _0715_ = in[7:0] == 8'he0;
  assign _0716_ = in[7:0] == 8'hdf;
  assign _0717_ = in[7:0] == 8'hde;
  assign _0718_ = in[7:0] == 8'hdd;
  assign _0719_ = in[7:0] == 8'hdc;
  assign _0720_ = in[7:0] == 8'hdb;
  assign _0721_ = in[7:0] == 8'hda;
  assign _0722_ = in[7:0] == 8'hd9;
  assign _0723_ = in[7:0] == 8'hd8;
  assign _0724_ = in[7:0] == 8'hd7;
  assign _0725_ = in[7:0] == 8'hd6;
  assign _0726_ = in[7:0] == 8'hd5;
  assign _0727_ = in[7:0] == 8'hd4;
  assign _0728_ = in[7:0] == 8'hd3;
  assign _0729_ = in[7:0] == 8'hd2;
  assign _0730_ = in[7:0] == 8'hd1;
  assign _0731_ = in[7:0] == 8'hd0;
  assign _0732_ = in[7:0] == 8'hcf;
  assign _0733_ = in[7:0] == 8'hce;
  assign _0734_ = in[7:0] == 8'hcd;
  assign _0735_ = in[7:0] == 8'hcc;
  assign _0736_ = in[7:0] == 8'hcb;
  assign _0737_ = in[7:0] == 8'hca;
  assign _0738_ = in[7:0] == 8'hc9;
  assign _0739_ = in[7:0] == 8'hc8;
  assign _0740_ = in[7:0] == 8'hc7;
  assign _0741_ = in[7:0] == 8'hc6;
  assign _0742_ = in[7:0] == 8'hc5;
  assign _0743_ = in[7:0] == 8'hc4;
  assign _0744_ = in[7:0] == 8'hc3;
  assign _0745_ = in[7:0] == 8'hc2;
  assign _0746_ = in[7:0] == 8'hc1;
  assign _0747_ = in[7:0] == 8'hc0;
  assign _0748_ = in[7:0] == 8'hbf;
  assign _0749_ = in[7:0] == 8'hbe;
  assign _0750_ = in[7:0] == 8'hbd;
  assign _0751_ = in[7:0] == 8'hbc;
  assign _0752_ = in[7:0] == 8'hbb;
  assign _0753_ = in[7:0] == 8'hba;
  assign _0754_ = in[7:0] == 8'hb9;
  assign _0755_ = in[7:0] == 8'hb8;
  assign _0756_ = in[7:0] == 8'hb7;
  assign _0757_ = in[7:0] == 8'hb6;
  assign _0758_ = in[7:0] == 8'hb5;
  assign _0759_ = in[7:0] == 8'hb4;
  assign _0760_ = in[7:0] == 8'hb3;
  assign _0761_ = in[7:0] == 8'hb2;
  assign _0762_ = in[7:0] == 8'hb1;
  assign _0763_ = in[7:0] == 8'hb0;
  assign _0764_ = in[7:0] == 8'haf;
  assign _0765_ = in[7:0] == 8'hae;
  assign _0766_ = in[7:0] == 8'had;
  assign _0767_ = in[7:0] == 8'hac;
  assign _0768_ = in[7:0] == 8'hab;
  assign _0769_ = in[7:0] == 8'haa;
  assign _0770_ = in[7:0] == 8'ha9;
  always @(posedge clk)
      \S4_0.S_3.out <= _0771_;
  assign _0772_ = in[31:24] == 8'ha8;
  assign _0773_ = in[31:24] == 8'ha7;
  assign _0774_ = in[31:24] == 8'ha6;
  assign _0775_ = in[31:24] == 8'ha5;
  assign _0776_ = in[31:24] == 8'ha4;
  assign _0777_ = in[31:24] == 8'ha3;
  assign _0778_ = in[31:24] == 8'ha2;
  assign _0779_ = in[31:24] == 8'ha1;
  assign _0780_ = in[31:24] == 8'ha0;
  assign _0781_ = in[31:24] == 8'h9f;
  assign _0782_ = in[31:24] == 8'h9e;
  assign _0783_ = in[31:24] == 8'h9d;
  assign _0784_ = in[31:24] == 8'h9c;
  assign _0785_ = in[31:24] == 8'h9b;
  assign _0786_ = in[31:24] == 8'h9a;
  assign _0787_ = in[31:24] == 8'h99;
  assign _0788_ = in[31:24] == 8'h98;
  assign _0789_ = in[31:24] == 8'h97;
  assign _0790_ = in[31:24] == 8'h96;
  assign _0791_ = in[31:24] == 8'h95;
  logic [255:0] fangyuan5;
  assign fangyuan5 = { _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_, _0943_, _0942_, _0941_, _0940_, _0939_, _0938_, _0937_, _0936_, _0935_, _0934_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_, _0774_, _0773_, _0772_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0944_, _0933_, _0922_, _0911_, _0900_, _0889_, _0878_, _0867_, _0856_, _0845_, _0834_, _0823_, _0812_ };

  always @(\S4_0.S_3.out or fangyuan5) begin
    casez (fangyuan5)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0771_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0771_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0771_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0771_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0771_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0771_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0771_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0771_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0771_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0771_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0771_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0771_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0771_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0771_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0771_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0771_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0771_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0771_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0771_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0771_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0771_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0771_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0771_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0771_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0771_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0771_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0771_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0771_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0771_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0771_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0771_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0771_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0771_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0771_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0771_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0771_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0771_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0771_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0771_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0771_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0771_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0771_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0771_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0771_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0771_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0771_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0771_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0771_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0771_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0771_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0771_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0771_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0771_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0771_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0771_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0771_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0771_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0771_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0771_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0771_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0771_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0771_ = 8'b01100011 ;
      default:
        _0771_ = \S4_0.S_3.out ;
    endcase
  end
  assign _0792_ = in[31:24] == 8'h94;
  assign _0793_ = in[31:24] == 8'h93;
  assign _0794_ = in[31:24] == 8'h92;
  assign _0795_ = in[31:24] == 8'h91;
  assign _0796_ = in[31:24] == 8'h90;
  assign _0797_ = in[31:24] == 8'h8f;
  assign _0798_ = in[31:24] == 8'h8e;
  assign _0799_ = in[31:24] == 8'h8d;
  assign _0800_ = in[31:24] == 8'h8c;
  assign _0801_ = in[31:24] == 8'h8b;
  assign _0802_ = in[31:24] == 8'h8a;
  assign _0803_ = in[31:24] == 8'h89;
  assign _0804_ = in[31:24] == 8'h88;
  assign _0805_ = in[31:24] == 8'h87;
  assign _0806_ = in[31:24] == 8'h86;
  assign _0807_ = in[31:24] == 8'h85;
  assign _0808_ = in[31:24] == 8'h84;
  assign _0809_ = in[31:24] == 8'h83;
  assign _0810_ = in[31:24] == 8'h82;
  assign _0811_ = in[31:24] == 8'h81;
  assign _0812_ = in[31:24] == 8'hff;
  assign _0813_ = in[31:24] == 8'h80;
  assign _0814_ = in[31:24] == 7'h7f;
  assign _0815_ = in[31:24] == 7'h7e;
  assign _0816_ = in[31:24] == 7'h7d;
  assign _0817_ = in[31:24] == 7'h7c;
  assign _0818_ = in[31:24] == 7'h7b;
  assign _0819_ = in[31:24] == 7'h7a;
  assign _0820_ = in[31:24] == 7'h79;
  assign _0821_ = in[31:24] == 7'h78;
  assign _0822_ = in[31:24] == 7'h77;
  assign _0823_ = in[31:24] == 8'hfe;
  assign _0824_ = in[31:24] == 7'h76;
  assign _0825_ = in[31:24] == 7'h75;
  assign _0826_ = in[31:24] == 7'h74;
  assign _0827_ = in[31:24] == 7'h73;
  assign _0828_ = in[31:24] == 7'h72;
  assign _0829_ = in[31:24] == 7'h71;
  assign _0830_ = in[31:24] == 7'h70;
  assign _0831_ = in[31:24] == 7'h6f;
  assign _0832_ = in[31:24] == 7'h6e;
  assign _0833_ = in[31:24] == 7'h6d;
  assign _0834_ = in[31:24] == 8'hfd;
  assign _0835_ = in[31:24] == 7'h6c;
  assign _0836_ = in[31:24] == 7'h6b;
  assign _0837_ = in[31:24] == 7'h6a;
  assign _0838_ = in[31:24] == 7'h69;
  assign _0839_ = in[31:24] == 7'h68;
  assign _0840_ = in[31:24] == 7'h67;
  assign _0841_ = in[31:24] == 7'h66;
  assign _0842_ = in[31:24] == 7'h65;
  assign _0843_ = in[31:24] == 7'h64;
  assign _0844_ = in[31:24] == 7'h63;
  assign _0845_ = in[31:24] == 8'hfc;
  assign _0846_ = in[31:24] == 7'h62;
  assign _0847_ = in[31:24] == 7'h61;
  assign _0848_ = in[31:24] == 7'h60;
  assign _0849_ = in[31:24] == 7'h5f;
  assign _0850_ = in[31:24] == 7'h5e;
  assign _0851_ = in[31:24] == 7'h5d;
  assign _0852_ = in[31:24] == 7'h5c;
  assign _0853_ = in[31:24] == 7'h5b;
  assign _0854_ = in[31:24] == 7'h5a;
  assign _0855_ = in[31:24] == 7'h59;
  assign _0856_ = in[31:24] == 8'hfb;
  assign _0857_ = in[31:24] == 7'h58;
  assign _0858_ = in[31:24] == 7'h57;
  assign _0859_ = in[31:24] == 7'h56;
  assign _0860_ = in[31:24] == 7'h55;
  assign _0861_ = in[31:24] == 7'h54;
  assign _0862_ = in[31:24] == 7'h53;
  assign _0863_ = in[31:24] == 7'h52;
  assign _0864_ = in[31:24] == 7'h51;
  assign _0865_ = in[31:24] == 7'h50;
  assign _0866_ = in[31:24] == 7'h4f;
  assign _0867_ = in[31:24] == 8'hfa;
  assign _0868_ = in[31:24] == 7'h4e;
  assign _0869_ = in[31:24] == 7'h4d;
  assign _0870_ = in[31:24] == 7'h4c;
  assign _0871_ = in[31:24] == 7'h4b;
  assign _0872_ = in[31:24] == 7'h4a;
  assign _0873_ = in[31:24] == 7'h49;
  assign _0874_ = in[31:24] == 7'h48;
  assign _0875_ = in[31:24] == 7'h47;
  assign _0876_ = in[31:24] == 7'h46;
  assign _0877_ = in[31:24] == 7'h45;
  assign _0878_ = in[31:24] == 8'hf9;
  assign _0879_ = in[31:24] == 7'h44;
  assign _0880_ = in[31:24] == 7'h43;
  assign _0881_ = in[31:24] == 7'h42;
  assign _0882_ = in[31:24] == 7'h41;
  assign _0883_ = in[31:24] == 7'h40;
  assign _0884_ = in[31:24] == 6'h3f;
  assign _0885_ = in[31:24] == 6'h3e;
  assign _0886_ = in[31:24] == 6'h3d;
  assign _0887_ = in[31:24] == 6'h3c;
  assign _0888_ = in[31:24] == 6'h3b;
  assign _0889_ = in[31:24] == 8'hf8;
  assign _0890_ = in[31:24] == 6'h3a;
  assign _0891_ = in[31:24] == 6'h39;
  assign _0892_ = in[31:24] == 6'h38;
  assign _0893_ = in[31:24] == 6'h37;
  assign _0894_ = in[31:24] == 6'h36;
  assign _0895_ = in[31:24] == 6'h35;
  assign _0896_ = in[31:24] == 6'h34;
  assign _0897_ = in[31:24] == 6'h33;
  assign _0898_ = in[31:24] == 6'h32;
  assign _0899_ = in[31:24] == 6'h31;
  assign _0900_ = in[31:24] == 8'hf7;
  assign _0901_ = in[31:24] == 6'h30;
  assign _0902_ = in[31:24] == 6'h2f;
  assign _0903_ = in[31:24] == 6'h2e;
  assign _0904_ = in[31:24] == 6'h2d;
  assign _0905_ = in[31:24] == 6'h2c;
  assign _0906_ = in[31:24] == 6'h2b;
  assign _0907_ = in[31:24] == 6'h2a;
  assign _0908_ = in[31:24] == 6'h29;
  assign _0909_ = in[31:24] == 6'h28;
  assign _0910_ = in[31:24] == 6'h27;
  assign _0911_ = in[31:24] == 8'hf6;
  assign _0912_ = in[31:24] == 6'h26;
  assign _0913_ = in[31:24] == 6'h25;
  assign _0914_ = in[31:24] == 6'h24;
  assign _0915_ = in[31:24] == 6'h23;
  assign _0916_ = in[31:24] == 6'h22;
  assign _0917_ = in[31:24] == 6'h21;
  assign _0918_ = in[31:24] == 6'h20;
  assign _0919_ = in[31:24] == 5'h1f;
  assign _0920_ = in[31:24] == 5'h1e;
  assign _0921_ = in[31:24] == 5'h1d;
  assign _0922_ = in[31:24] == 8'hf5;
  assign _0923_ = in[31:24] == 5'h1c;
  assign _0924_ = in[31:24] == 5'h1b;
  assign _0925_ = in[31:24] == 5'h1a;
  assign _0926_ = in[31:24] == 5'h19;
  assign _0927_ = in[31:24] == 5'h18;
  assign _0928_ = in[31:24] == 5'h17;
  assign _0929_ = in[31:24] == 5'h16;
  assign _0930_ = in[31:24] == 5'h15;
  assign _0931_ = in[31:24] == 5'h14;
  assign _0932_ = in[31:24] == 5'h13;
  assign _0933_ = in[31:24] == 8'hf4;
  assign _0934_ = in[31:24] == 5'h12;
  assign _0935_ = in[31:24] == 5'h11;
  assign _0936_ = in[31:24] == 5'h10;
  assign _0937_ = in[31:24] == 4'hf;
  assign _0938_ = in[31:24] == 4'he;
  assign _0939_ = in[31:24] == 4'hd;
  assign _0940_ = in[31:24] == 4'hc;
  assign _0941_ = in[31:24] == 4'hb;
  assign _0942_ = in[31:24] == 4'ha;
  assign _0943_ = in[31:24] == 4'h9;
  assign _0944_ = in[31:24] == 8'hf3;
  assign _0945_ = in[31:24] == 4'h8;
  assign _0946_ = in[31:24] == 3'h7;
  assign _0947_ = in[31:24] == 3'h6;
  assign _0948_ = in[31:24] == 3'h5;
  assign _0949_ = in[31:24] == 3'h4;
  assign _0950_ = in[31:24] == 2'h3;
  assign _0951_ = in[31:24] == 2'h2;
  assign _0952_ = in[31:24] == 1'h1;
  assign _0953_ = ! in[31:24];
  assign _0954_ = in[31:24] == 8'hf2;
  assign _0955_ = in[31:24] == 8'hf1;
  assign _0956_ = in[31:24] == 8'hf0;
  assign _0957_ = in[31:24] == 8'hef;
  assign _0958_ = in[31:24] == 8'hee;
  assign _0959_ = in[31:24] == 8'hed;
  assign _0960_ = in[31:24] == 8'hec;
  assign _0961_ = in[31:24] == 8'heb;
  assign _0962_ = in[31:24] == 8'hea;
  assign _0963_ = in[31:24] == 8'he9;
  assign _0964_ = in[31:24] == 8'he8;
  assign _0965_ = in[31:24] == 8'he7;
  assign _0966_ = in[31:24] == 8'he6;
  assign _0967_ = in[31:24] == 8'he5;
  assign _0968_ = in[31:24] == 8'he4;
  assign _0969_ = in[31:24] == 8'he3;
  assign _0970_ = in[31:24] == 8'he2;
  assign _0971_ = in[31:24] == 8'he1;
  assign _0972_ = in[31:24] == 8'he0;
  assign _0973_ = in[31:24] == 8'hdf;
  assign _0974_ = in[31:24] == 8'hde;
  assign _0975_ = in[31:24] == 8'hdd;
  assign _0976_ = in[31:24] == 8'hdc;
  assign _0977_ = in[31:24] == 8'hdb;
  assign _0978_ = in[31:24] == 8'hda;
  assign _0979_ = in[31:24] == 8'hd9;
  assign _0980_ = in[31:24] == 8'hd8;
  assign _0981_ = in[31:24] == 8'hd7;
  assign _0982_ = in[31:24] == 8'hd6;
  assign _0983_ = in[31:24] == 8'hd5;
  assign _0984_ = in[31:24] == 8'hd4;
  assign _0985_ = in[31:24] == 8'hd3;
  assign _0986_ = in[31:24] == 8'hd2;
  assign _0987_ = in[31:24] == 8'hd1;
  assign _0988_ = in[31:24] == 8'hd0;
  assign _0989_ = in[31:24] == 8'hcf;
  assign _0990_ = in[31:24] == 8'hce;
  assign _0991_ = in[31:24] == 8'hcd;
  assign _0992_ = in[31:24] == 8'hcc;
  assign _0993_ = in[31:24] == 8'hcb;
  assign _0994_ = in[31:24] == 8'hca;
  assign _0995_ = in[31:24] == 8'hc9;
  assign _0996_ = in[31:24] == 8'hc8;
  assign _0997_ = in[31:24] == 8'hc7;
  assign _0998_ = in[31:24] == 8'hc6;
  assign _0999_ = in[31:24] == 8'hc5;
  assign _1000_ = in[31:24] == 8'hc4;
  assign _1001_ = in[31:24] == 8'hc3;
  assign _1002_ = in[31:24] == 8'hc2;
  assign _1003_ = in[31:24] == 8'hc1;
  assign _1004_ = in[31:24] == 8'hc0;
  assign _1005_ = in[31:24] == 8'hbf;
  assign _1006_ = in[31:24] == 8'hbe;
  assign _1007_ = in[31:24] == 8'hbd;
  assign _1008_ = in[31:24] == 8'hbc;
  assign _1009_ = in[31:24] == 8'hbb;
  assign _1010_ = in[31:24] == 8'hba;
  assign _1011_ = in[31:24] == 8'hb9;
  assign _1012_ = in[31:24] == 8'hb8;
  assign _1013_ = in[31:24] == 8'hb7;
  assign _1014_ = in[31:24] == 8'hb6;
  assign _1015_ = in[31:24] == 8'hb5;
  assign _1016_ = in[31:24] == 8'hb4;
  assign _1017_ = in[31:24] == 8'hb3;
  assign _1018_ = in[31:24] == 8'hb2;
  assign _1019_ = in[31:24] == 8'hb1;
  assign _1020_ = in[31:24] == 8'hb0;
  assign _1021_ = in[31:24] == 8'haf;
  assign _1022_ = in[31:24] == 8'hae;
  assign _1023_ = in[31:24] == 8'had;
  assign _1024_ = in[31:24] == 8'hac;
  assign _1025_ = in[31:24] == 8'hab;
  assign _1026_ = in[31:24] == 8'haa;
  assign _1027_ = in[31:24] == 8'ha9;
  assign v0[31:24] = in[127:120] ^ rcon;
  logic [31:0] fangyuan6;
  assign fangyuan6 = { v0[31:24], in[119:96] };

  assign v1 = fangyuan6 ^ in[95:64];
  assign v2 = v1 ^ in[63:32];
  assign v3 = v2 ^ in[31:0];
  logic [31:0] fangyuan7;
  assign fangyuan7 = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out };

  assign k0b = k0a ^ fangyuan7;
  logic [31:0] fangyuan8;
  assign fangyuan8 = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out };

  assign k1b = k1a ^ fangyuan8;
  logic [31:0] fangyuan9;
  assign fangyuan9 = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out };

  assign k2b = k2a ^ fangyuan9;
  logic [31:0] fangyuan10;
  assign fangyuan10 = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out };

  assign k3b = k3a ^ fangyuan10;
  assign \S4_0.S_0.clk = clk;
  assign \S4_0.S_0.in = in[23:16];
  assign \S4_0.S_1.clk = clk;
  assign \S4_0.S_1.in = in[15:8];
  assign \S4_0.S_2.clk = clk;
  assign \S4_0.S_2.in = in[7:0];
  assign \S4_0.S_3.clk = clk;
  assign \S4_0.S_3.in = in[31:24];
  assign \S4_0.clk = clk;
  assign \S4_0.in = { in[23:0], in[31:24] };
  assign \S4_0.out = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out };
  assign k0 = in[127:96];
  assign k1 = in[95:64];
  assign k2 = in[63:32];
  assign k3 = in[31:0];
  assign k4a = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out };
  assign out_2 = { k0b, k1b, k2b, k3b };
  assign v0[23:0] = in[119:96];
endmodule
