module bar__DOT__i1(
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
i_wb_data,
kp,
ki,
kd,
sp,
pv,
RS,
un,
__COUNTER_start__n0
);
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg     [31:0] i_wb_data;
output reg     [15:0] kp;
output reg     [15:0] ki;
output reg     [15:0] kd;
output reg     [15:0] sp;
output reg     [15:0] pv;
output reg            RS;
output reg     [31:0] un;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire            bv_1_0_n2;
wire            bv_1_1_n5;
wire            clk;
wire            n1;
wire            n10;
wire            n100;
wire            n1000;
wire            n10000;
wire            n10001;
wire            n10002;
wire            n10003;
wire            n10004;
wire            n10005;
wire            n10006;
wire            n10007;
wire            n10008;
wire            n10009;
wire            n1001;
wire            n10010;
wire            n10011;
wire            n10012;
wire            n10013;
wire            n10014;
wire            n10015;
wire            n10016;
wire            n10017;
wire            n10018;
wire            n10019;
wire            n1002;
wire            n10020;
wire            n10021;
wire            n10022;
wire            n10023;
wire            n10024;
wire            n10025;
wire            n10026;
wire            n10027;
wire            n10028;
wire            n10029;
wire            n1003;
wire            n10030;
wire            n10031;
wire            n10032;
wire            n10033;
wire            n10034;
wire            n10035;
wire            n10036;
wire            n10037;
wire            n10038;
wire            n10039;
wire            n1004;
wire            n10040;
wire            n10041;
wire            n10042;
wire            n10043;
wire            n10044;
wire            n10045;
wire            n10046;
wire            n10047;
wire            n10048;
wire            n10049;
wire            n1005;
wire            n10050;
wire            n10051;
wire            n10052;
wire            n10053;
wire            n10054;
wire            n10055;
wire            n10056;
wire            n10057;
wire            n10058;
wire            n10059;
wire            n1006;
wire            n10060;
wire            n10061;
wire            n10062;
wire            n10063;
wire            n10064;
wire            n10065;
wire            n10066;
wire            n10067;
wire            n10068;
wire            n10069;
wire            n1007;
wire            n10070;
wire            n10071;
wire            n10072;
wire            n10073;
wire            n10074;
wire            n10075;
wire            n10076;
wire            n10077;
wire            n10078;
wire            n10079;
wire            n1008;
wire            n10080;
wire            n10081;
wire            n10082;
wire            n10083;
wire            n10084;
wire            n10085;
wire            n10086;
wire            n10087;
wire            n10088;
wire            n10089;
wire            n1009;
wire            n10090;
wire            n10091;
wire            n10092;
wire            n10093;
wire            n10094;
wire            n10095;
wire            n10096;
wire            n10097;
wire            n10098;
wire            n10099;
wire            n101;
wire            n1010;
wire            n10100;
wire            n10101;
wire            n10102;
wire            n10103;
wire            n10104;
wire            n10105;
wire            n10106;
wire            n10107;
wire            n10108;
wire            n10109;
wire            n1011;
wire            n10110;
wire            n10111;
wire            n10112;
wire            n10113;
wire            n10114;
wire            n10115;
wire            n10116;
wire            n10117;
wire            n10118;
wire            n10119;
wire            n1012;
wire            n10120;
wire            n10121;
wire            n10122;
wire            n10123;
wire            n10124;
wire            n10125;
wire            n10126;
wire            n10127;
wire            n10128;
wire            n10129;
wire            n1013;
wire            n10130;
wire            n10131;
wire            n10132;
wire            n10133;
wire            n10134;
wire            n10135;
wire            n10136;
wire            n10137;
wire            n10138;
wire            n10139;
wire            n1014;
wire            n10140;
wire            n10141;
wire            n10142;
wire            n10143;
wire            n10144;
wire            n10145;
wire            n10146;
wire            n10147;
wire            n10148;
wire            n10149;
wire            n1015;
wire            n10150;
wire            n10151;
wire            n10152;
wire            n10153;
wire            n10154;
wire            n10155;
wire            n10156;
wire            n10157;
wire            n10158;
wire            n10159;
wire            n1016;
wire            n10160;
wire            n10161;
wire            n10162;
wire            n10163;
wire            n10164;
wire            n10165;
wire            n10166;
wire            n10167;
wire            n10168;
wire            n10169;
wire            n1017;
wire            n10170;
wire            n10171;
wire            n10172;
wire            n10173;
wire            n10174;
wire            n10175;
wire            n10176;
wire            n10177;
wire            n10178;
wire            n10179;
wire            n1018;
wire            n10180;
wire            n10181;
wire            n10182;
wire            n10183;
wire            n10184;
wire            n10185;
wire            n10186;
wire            n10187;
wire            n10188;
wire            n10189;
wire            n1019;
wire            n10190;
wire            n10191;
wire            n10192;
wire            n10193;
wire            n10194;
wire            n10195;
wire            n10196;
wire            n10197;
wire            n10198;
wire            n10199;
wire            n102;
wire            n1020;
wire            n10200;
wire            n10201;
wire            n10202;
wire            n10203;
wire            n10204;
wire            n10205;
wire            n10206;
wire            n10207;
wire            n10208;
wire            n10209;
wire            n1021;
wire            n10210;
wire            n10211;
wire            n10212;
wire            n10213;
wire            n10214;
wire            n10215;
wire            n10216;
wire            n10217;
wire            n10218;
wire            n10219;
wire            n1022;
wire            n10220;
wire            n10221;
wire            n10222;
wire            n10223;
wire            n10224;
wire            n10225;
wire            n10226;
wire            n10227;
wire            n10228;
wire            n10229;
wire            n1023;
wire            n10230;
wire            n10231;
wire            n10232;
wire            n10233;
wire            n10234;
wire            n10235;
wire            n10236;
wire            n10237;
wire            n10238;
wire            n10239;
wire            n1024;
wire            n10240;
wire            n10241;
wire            n10242;
wire            n10243;
wire            n10244;
wire            n10245;
wire            n10246;
wire            n10247;
wire            n10248;
wire            n10249;
wire            n1025;
wire            n10250;
wire            n10251;
wire            n10252;
wire            n10253;
wire            n10254;
wire            n10255;
wire            n10256;
wire            n10257;
wire            n10258;
wire            n10259;
wire            n1026;
wire            n10260;
wire            n10261;
wire            n10262;
wire            n10263;
wire            n10264;
wire            n10265;
wire            n10266;
wire            n10267;
wire            n10268;
wire            n10269;
wire            n1027;
wire            n10270;
wire            n10271;
wire            n10272;
wire            n10273;
wire            n10274;
wire            n10275;
wire            n10276;
wire            n10277;
wire            n10278;
wire            n10279;
wire            n1028;
wire            n10280;
wire            n10281;
wire            n10282;
wire            n10283;
wire            n10284;
wire            n10285;
wire            n10286;
wire            n10287;
wire            n10288;
wire            n10289;
wire            n1029;
wire            n10290;
wire            n10291;
wire            n10292;
wire            n10293;
wire            n10294;
wire            n10295;
wire            n10296;
wire            n10297;
wire            n10298;
wire            n10299;
wire            n103;
wire            n1030;
wire            n10300;
wire            n10301;
wire            n10302;
wire            n10303;
wire            n10304;
wire            n10305;
wire            n10306;
wire            n10307;
wire            n10308;
wire            n10309;
wire            n1031;
wire            n10310;
wire            n10311;
wire            n10312;
wire            n10313;
wire            n10314;
wire            n10315;
wire            n10316;
wire            n10317;
wire            n10318;
wire            n10319;
wire            n1032;
wire            n10320;
wire            n10321;
wire            n10322;
wire            n10323;
wire            n10324;
wire            n10325;
wire            n10326;
wire            n10327;
wire            n10328;
wire            n10329;
wire            n1033;
wire            n10330;
wire            n10331;
wire            n10332;
wire            n10333;
wire            n10334;
wire            n10335;
wire            n10336;
wire            n10337;
wire            n10338;
wire            n10339;
wire            n1034;
wire            n10340;
wire            n10341;
wire            n10342;
wire            n10343;
wire            n10344;
wire            n10345;
wire            n10346;
wire            n10347;
wire            n10348;
wire            n10349;
wire            n1035;
wire            n10350;
wire            n10351;
wire            n10352;
wire            n10353;
wire            n10354;
wire            n10355;
wire            n10356;
wire            n10357;
wire            n10358;
wire            n10359;
wire            n1036;
wire            n10360;
wire            n10361;
wire            n10362;
wire            n10363;
wire            n10364;
wire            n10365;
wire            n10366;
wire            n10367;
wire            n10368;
wire            n10369;
wire            n1037;
wire            n10370;
wire            n10371;
wire            n10372;
wire            n10373;
wire            n10374;
wire            n10375;
wire            n10376;
wire            n10377;
wire            n10378;
wire            n10379;
wire            n1038;
wire            n10380;
wire            n10381;
wire            n10382;
wire            n10383;
wire            n10384;
wire            n10385;
wire            n10386;
wire            n10387;
wire            n10388;
wire            n10389;
wire            n1039;
wire            n10390;
wire            n10391;
wire            n10392;
wire            n10393;
wire            n10394;
wire            n10395;
wire            n10396;
wire            n10397;
wire            n10398;
wire            n10399;
wire            n104;
wire            n1040;
wire            n10400;
wire            n10401;
wire            n10402;
wire            n10403;
wire            n10404;
wire            n10405;
wire            n10406;
wire            n10407;
wire            n10408;
wire            n10409;
wire            n1041;
wire            n10410;
wire            n10411;
wire            n10412;
wire            n10413;
wire            n10414;
wire            n10415;
wire            n10416;
wire            n10417;
wire            n10418;
wire            n10419;
wire            n1042;
wire            n10420;
wire            n10421;
wire            n10422;
wire            n10423;
wire            n10424;
wire            n10425;
wire            n10426;
wire            n10427;
wire            n10428;
wire            n10429;
wire            n1043;
wire            n10430;
wire            n10431;
wire            n10432;
wire            n10433;
wire            n10434;
wire            n10435;
wire            n10436;
wire            n10437;
wire            n10438;
wire            n10439;
wire            n1044;
wire            n10440;
wire            n10441;
wire            n10442;
wire            n10443;
wire            n10444;
wire            n10445;
wire            n10446;
wire            n10447;
wire            n10448;
wire            n10449;
wire            n1045;
wire            n10450;
wire            n10451;
wire            n10452;
wire            n10453;
wire            n10454;
wire            n10455;
wire            n10456;
wire            n10457;
wire            n10458;
wire            n10459;
wire            n1046;
wire            n10460;
wire            n10461;
wire            n10462;
wire            n10463;
wire            n10464;
wire            n10465;
wire            n10466;
wire            n10467;
wire            n10468;
wire            n10469;
wire            n1047;
wire            n10470;
wire            n10471;
wire            n10472;
wire            n10473;
wire            n10474;
wire            n10475;
wire            n10476;
wire            n10477;
wire            n10478;
wire            n10479;
wire            n1048;
wire            n10480;
wire            n10481;
wire            n10482;
wire            n10483;
wire            n10484;
wire            n10485;
wire            n10486;
wire            n10487;
wire            n10488;
wire            n10489;
wire            n1049;
wire            n10490;
wire            n10491;
wire            n10492;
wire            n10493;
wire            n10494;
wire            n10495;
wire            n10496;
wire            n10497;
wire            n10498;
wire            n10499;
wire            n105;
wire            n1050;
wire            n10500;
wire            n10501;
wire            n10502;
wire            n10503;
wire            n10504;
wire            n10505;
wire            n10506;
wire            n10507;
wire            n10508;
wire            n10509;
wire            n1051;
wire            n10510;
wire            n10511;
wire            n10512;
wire            n10513;
wire            n10514;
wire            n10515;
wire            n10516;
wire            n10517;
wire            n10518;
wire            n10519;
wire            n1052;
wire            n10520;
wire            n10521;
wire            n10522;
wire            n10523;
wire            n10524;
wire            n10525;
wire            n10526;
wire            n10527;
wire            n10528;
wire            n10529;
wire            n1053;
wire            n10530;
wire            n10531;
wire            n10532;
wire            n10533;
wire            n10534;
wire            n10535;
wire            n10536;
wire            n10537;
wire            n10538;
wire            n10539;
wire            n1054;
wire            n10540;
wire            n10541;
wire            n10542;
wire            n10543;
wire            n10544;
wire            n10545;
wire            n10546;
wire            n10547;
wire            n10548;
wire            n10549;
wire            n1055;
wire            n10550;
wire            n10551;
wire            n10552;
wire            n10553;
wire            n10554;
wire            n10555;
wire            n10556;
wire            n10557;
wire            n10558;
wire            n10559;
wire            n1056;
wire            n10560;
wire            n10561;
wire            n10562;
wire            n10563;
wire            n10564;
wire            n10565;
wire            n10566;
wire            n10567;
wire            n10568;
wire            n10569;
wire            n1057;
wire            n10570;
wire            n10571;
wire            n10572;
wire            n10573;
wire            n10574;
wire            n10575;
wire            n10576;
wire            n10577;
wire            n10578;
wire            n10579;
wire            n1058;
wire            n10580;
wire            n10581;
wire            n10582;
wire            n10583;
wire            n10584;
wire            n10585;
wire            n10586;
wire            n10587;
wire            n10588;
wire            n10589;
wire            n1059;
wire            n10590;
wire            n10591;
wire            n10592;
wire            n10593;
wire            n10594;
wire            n10595;
wire            n10596;
wire            n10597;
wire            n10598;
wire            n10599;
wire            n106;
wire            n1060;
wire            n10600;
wire            n10601;
wire            n10602;
wire            n10603;
wire            n10604;
wire            n10605;
wire            n10606;
wire            n10607;
wire            n10608;
wire            n10609;
wire            n1061;
wire            n10610;
wire            n10611;
wire            n10612;
wire            n10613;
wire            n10614;
wire            n10615;
wire            n10616;
wire            n10617;
wire            n10618;
wire            n10619;
wire            n1062;
wire            n10620;
wire            n10621;
wire            n10622;
wire            n10623;
wire            n10624;
wire            n10625;
wire            n10626;
wire            n10627;
wire            n10628;
wire            n10629;
wire            n1063;
wire            n10630;
wire            n10631;
wire            n10632;
wire            n10633;
wire            n10634;
wire            n10635;
wire            n10636;
wire            n10637;
wire            n10638;
wire            n10639;
wire            n1064;
wire            n10640;
wire            n10641;
wire            n10642;
wire            n10643;
wire            n10644;
wire            n10645;
wire            n10646;
wire            n10647;
wire            n10648;
wire            n10649;
wire            n1065;
wire            n10650;
wire            n10651;
wire            n10652;
wire            n10653;
wire            n10654;
wire            n10655;
wire            n10656;
wire            n10657;
wire            n10658;
wire            n10659;
wire            n1066;
wire            n10660;
wire            n10661;
wire            n10662;
wire            n10663;
wire            n10664;
wire            n10665;
wire            n10666;
wire            n10667;
wire            n10668;
wire            n10669;
wire            n1067;
wire            n10670;
wire            n10671;
wire            n10672;
wire            n10673;
wire            n10674;
wire            n10675;
wire            n10676;
wire            n10677;
wire            n10678;
wire            n10679;
wire            n1068;
wire            n10680;
wire            n10681;
wire            n10682;
wire            n10683;
wire            n10684;
wire            n10685;
wire            n10686;
wire            n10687;
wire            n10688;
wire            n10689;
wire            n1069;
wire            n10690;
wire            n10691;
wire            n10692;
wire            n10693;
wire            n10694;
wire            n10695;
wire            n10696;
wire            n10697;
wire            n10698;
wire            n10699;
wire            n107;
wire            n1070;
wire            n10700;
wire            n10701;
wire            n10702;
wire            n10703;
wire            n10704;
wire            n10705;
wire            n10706;
wire            n10707;
wire            n10708;
wire            n10709;
wire            n1071;
wire            n10710;
wire            n10711;
wire            n10712;
wire            n10713;
wire            n10714;
wire            n10715;
wire            n10716;
wire            n10717;
wire            n10718;
wire            n10719;
wire            n1072;
wire            n10720;
wire            n10721;
wire            n10722;
wire            n10723;
wire            n10724;
wire            n10725;
wire            n10726;
wire            n10727;
wire            n10728;
wire            n10729;
wire            n1073;
wire            n10730;
wire            n10731;
wire            n10732;
wire            n10733;
wire            n10734;
wire            n10735;
wire            n10736;
wire            n10737;
wire            n10738;
wire            n10739;
wire            n1074;
wire            n10740;
wire            n10741;
wire            n10742;
wire            n10743;
wire            n10744;
wire            n10745;
wire            n10746;
wire            n10747;
wire            n10748;
wire            n10749;
wire            n1075;
wire            n10750;
wire            n10751;
wire            n10752;
wire            n10753;
wire            n10754;
wire            n10755;
wire            n10756;
wire            n10757;
wire            n10758;
wire            n10759;
wire            n1076;
wire            n10760;
wire            n10761;
wire            n10762;
wire            n10763;
wire            n10764;
wire            n10765;
wire            n10766;
wire            n10767;
wire            n10768;
wire            n10769;
wire            n1077;
wire            n10770;
wire            n10771;
wire            n10772;
wire            n10773;
wire            n10774;
wire            n10775;
wire            n10776;
wire            n10777;
wire            n10778;
wire            n10779;
wire            n1078;
wire            n10780;
wire            n10781;
wire            n10782;
wire            n10783;
wire            n10784;
wire            n10785;
wire            n10786;
wire            n10787;
wire            n10788;
wire            n10789;
wire            n1079;
wire            n10790;
wire            n10791;
wire            n10792;
wire            n10793;
wire            n10794;
wire            n10795;
wire            n10796;
wire            n10797;
wire            n10798;
wire            n10799;
wire            n108;
wire            n1080;
wire            n10800;
wire            n10801;
wire            n10802;
wire            n10803;
wire            n10804;
wire            n10805;
wire            n10806;
wire            n10807;
wire            n10808;
wire            n10809;
wire            n1081;
wire            n10810;
wire            n10811;
wire            n10812;
wire            n10813;
wire            n10814;
wire            n10815;
wire            n10816;
wire            n10817;
wire            n10818;
wire            n10819;
wire            n1082;
wire            n10820;
wire            n10821;
wire            n10822;
wire            n10823;
wire            n10824;
wire            n10825;
wire            n10826;
wire            n10827;
wire            n10828;
wire            n10829;
wire            n1083;
wire            n10830;
wire            n10831;
wire            n10832;
wire            n10833;
wire            n10834;
wire            n10835;
wire            n10836;
wire            n10837;
wire            n10838;
wire            n10839;
wire            n1084;
wire            n10840;
wire            n10841;
wire            n10842;
wire            n10843;
wire            n10844;
wire            n10845;
wire            n10846;
wire            n10847;
wire            n10848;
wire            n10849;
wire            n1085;
wire            n10850;
wire            n10851;
wire            n10852;
wire            n10853;
wire            n10854;
wire            n10855;
wire            n10856;
wire            n10857;
wire            n10858;
wire            n10859;
wire            n1086;
wire            n10860;
wire            n10861;
wire            n10862;
wire            n10863;
wire            n10864;
wire            n10865;
wire            n10866;
wire            n10867;
wire            n10868;
wire            n10869;
wire            n1087;
wire            n10870;
wire            n10871;
wire            n10872;
wire            n10873;
wire            n10874;
wire            n10875;
wire            n10876;
wire            n10877;
wire            n10878;
wire            n10879;
wire            n1088;
wire            n10880;
wire            n10881;
wire            n10882;
wire            n10883;
wire            n10884;
wire            n10885;
wire            n10886;
wire            n10887;
wire            n10888;
wire            n10889;
wire            n1089;
wire            n10890;
wire            n10891;
wire            n10892;
wire            n10893;
wire            n10894;
wire            n10895;
wire            n10896;
wire            n10897;
wire            n10898;
wire            n10899;
wire            n109;
wire            n1090;
wire            n10900;
wire            n10901;
wire            n10902;
wire            n10903;
wire            n10904;
wire            n10905;
wire            n10906;
wire            n10907;
wire            n10908;
wire            n10909;
wire            n1091;
wire            n10910;
wire            n10911;
wire            n10912;
wire            n10913;
wire            n10914;
wire            n10915;
wire            n10916;
wire            n10917;
wire            n10918;
wire            n10919;
wire            n1092;
wire            n10920;
wire            n10921;
wire            n10922;
wire            n10923;
wire            n10924;
wire            n10925;
wire            n10926;
wire            n10927;
wire            n10928;
wire            n10929;
wire            n1093;
wire            n10930;
wire            n10931;
wire            n10932;
wire            n10933;
wire            n10934;
wire            n10935;
wire            n10936;
wire            n10937;
wire            n10938;
wire            n10939;
wire            n1094;
wire            n10940;
wire            n10941;
wire            n10942;
wire            n10943;
wire            n10944;
wire            n10945;
wire            n10946;
wire            n10947;
wire            n10948;
wire            n10949;
wire            n1095;
wire            n10950;
wire            n10951;
wire            n10952;
wire            n10953;
wire            n10954;
wire            n10955;
wire            n10956;
wire            n10957;
wire            n10958;
wire            n10959;
wire            n1096;
wire            n10960;
wire            n10961;
wire            n10962;
wire            n10963;
wire            n10964;
wire            n10965;
wire            n10966;
wire            n10967;
wire            n10968;
wire            n10969;
wire            n1097;
wire            n10970;
wire            n10971;
wire            n10972;
wire            n10973;
wire            n10974;
wire            n10975;
wire            n10976;
wire            n10977;
wire            n10978;
wire            n10979;
wire            n1098;
wire            n10980;
wire            n10981;
wire            n10982;
wire            n10983;
wire            n10984;
wire            n10985;
wire            n10986;
wire            n10987;
wire            n10988;
wire            n10989;
wire            n1099;
wire            n10990;
wire            n10991;
wire            n10992;
wire            n10993;
wire            n10994;
wire            n10995;
wire            n10996;
wire            n10997;
wire            n10998;
wire            n10999;
wire            n11;
wire            n110;
wire            n1100;
wire            n11000;
wire            n11001;
wire            n11002;
wire            n11003;
wire            n11004;
wire            n11005;
wire            n11006;
wire            n11007;
wire            n11008;
wire            n11009;
wire            n1101;
wire            n11010;
wire            n11011;
wire            n11012;
wire            n11013;
wire            n11014;
wire            n11015;
wire            n11016;
wire            n11017;
wire            n11018;
wire            n11019;
wire            n1102;
wire            n11020;
wire            n11021;
wire            n11022;
wire            n11023;
wire            n11024;
wire            n11025;
wire            n11026;
wire            n11027;
wire            n11028;
wire            n11029;
wire            n1103;
wire            n11030;
wire            n11031;
wire            n11032;
wire            n11033;
wire            n11034;
wire            n11035;
wire            n11036;
wire            n11037;
wire            n11038;
wire            n11039;
wire            n1104;
wire            n11040;
wire            n11041;
wire            n11042;
wire            n11043;
wire            n11044;
wire            n11045;
wire            n11046;
wire            n11047;
wire            n11048;
wire            n11049;
wire            n1105;
wire            n11050;
wire            n11051;
wire            n11052;
wire            n11053;
wire            n11054;
wire            n11055;
wire            n11056;
wire            n11057;
wire            n11058;
wire            n11059;
wire            n1106;
wire            n11060;
wire            n11061;
wire            n11062;
wire            n11063;
wire            n11064;
wire            n11065;
wire            n11066;
wire            n11067;
wire            n11068;
wire            n11069;
wire            n1107;
wire            n11070;
wire            n11071;
wire            n11072;
wire            n11073;
wire            n11074;
wire            n11075;
wire            n11076;
wire            n11077;
wire            n11078;
wire            n11079;
wire            n1108;
wire            n11080;
wire            n11081;
wire            n11082;
wire            n11083;
wire            n11084;
wire            n11085;
wire            n11086;
wire            n11087;
wire            n11088;
wire            n11089;
wire            n1109;
wire            n11090;
wire            n11091;
wire            n11092;
wire            n11093;
wire            n11094;
wire            n11095;
wire            n11096;
wire            n11097;
wire            n11098;
wire            n11099;
wire            n111;
wire            n1110;
wire            n11100;
wire            n11101;
wire            n11102;
wire            n11103;
wire            n11104;
wire            n11105;
wire            n11106;
wire            n11107;
wire            n11108;
wire            n11109;
wire            n1111;
wire            n11110;
wire            n11111;
wire            n11112;
wire            n11113;
wire            n11114;
wire            n11115;
wire            n11116;
wire            n11117;
wire            n11118;
wire            n11119;
wire            n1112;
wire            n11120;
wire            n11121;
wire            n11122;
wire            n11123;
wire            n11124;
wire            n11125;
wire            n11126;
wire            n11127;
wire            n11128;
wire            n11129;
wire            n1113;
wire            n11130;
wire            n11131;
wire            n11132;
wire            n11133;
wire            n11134;
wire            n11135;
wire            n11136;
wire            n11137;
wire            n11138;
wire            n11139;
wire            n1114;
wire            n11140;
wire            n11141;
wire            n11142;
wire            n11143;
wire            n11144;
wire            n11145;
wire            n11146;
wire            n11147;
wire            n11148;
wire            n11149;
wire            n1115;
wire            n11150;
wire            n11151;
wire            n11152;
wire            n11153;
wire            n11154;
wire            n11155;
wire            n11156;
wire            n11157;
wire            n11158;
wire            n11159;
wire            n1116;
wire            n11160;
wire            n11161;
wire            n11162;
wire            n11163;
wire            n11164;
wire            n11165;
wire            n11166;
wire            n11167;
wire            n11168;
wire            n11169;
wire            n1117;
wire            n11170;
wire            n11171;
wire            n11172;
wire            n11173;
wire            n11174;
wire            n11175;
wire            n11176;
wire            n11177;
wire            n11178;
wire            n11179;
wire            n1118;
wire            n11180;
wire            n11181;
wire            n11182;
wire            n11183;
wire            n11184;
wire            n11185;
wire            n11186;
wire            n11187;
wire            n11188;
wire            n11189;
wire            n1119;
wire            n11190;
wire            n11191;
wire            n11192;
wire            n11193;
wire            n11194;
wire            n11195;
wire            n11196;
wire            n11197;
wire            n11198;
wire            n11199;
wire            n112;
wire            n1120;
wire            n11200;
wire            n11201;
wire            n11202;
wire            n11203;
wire            n11204;
wire            n11205;
wire            n11206;
wire            n11207;
wire            n11208;
wire            n11209;
wire            n1121;
wire            n11210;
wire            n11211;
wire            n11212;
wire            n11213;
wire            n11214;
wire            n11215;
wire            n11216;
wire            n11217;
wire            n11218;
wire            n11219;
wire            n1122;
wire            n11220;
wire            n11221;
wire            n11222;
wire            n11223;
wire            n11224;
wire            n11225;
wire            n11226;
wire            n11227;
wire            n11228;
wire            n11229;
wire            n1123;
wire            n11230;
wire            n11231;
wire            n11232;
wire            n11233;
wire            n11234;
wire            n11235;
wire            n11236;
wire            n11237;
wire            n11238;
wire            n11239;
wire            n1124;
wire            n11240;
wire            n11241;
wire            n11242;
wire            n11243;
wire            n11244;
wire            n11245;
wire            n11246;
wire            n11247;
wire            n11248;
wire            n11249;
wire            n1125;
wire            n11250;
wire            n11251;
wire            n11252;
wire            n11253;
wire            n11254;
wire            n11255;
wire            n11256;
wire            n11257;
wire            n11258;
wire            n11259;
wire            n1126;
wire            n11260;
wire            n11261;
wire            n11262;
wire            n11263;
wire            n11264;
wire            n11265;
wire            n11266;
wire            n11267;
wire            n11268;
wire            n11269;
wire            n1127;
wire            n11270;
wire            n11271;
wire            n11272;
wire            n11273;
wire            n11274;
wire            n11275;
wire            n11276;
wire            n11277;
wire            n11278;
wire            n11279;
wire            n1128;
wire            n11280;
wire            n11281;
wire            n11282;
wire            n11283;
wire            n11284;
wire            n11285;
wire            n11286;
wire            n11287;
wire            n11288;
wire            n11289;
wire            n1129;
wire            n11290;
wire            n11291;
wire            n11292;
wire            n11293;
wire            n11294;
wire            n11295;
wire            n11296;
wire            n11297;
wire            n11298;
wire            n11299;
wire            n113;
wire            n1130;
wire            n11300;
wire            n11301;
wire            n11302;
wire            n11303;
wire            n11304;
wire            n11305;
wire            n11306;
wire            n11307;
wire            n11308;
wire            n11309;
wire            n1131;
wire            n11310;
wire            n11311;
wire            n11312;
wire            n11313;
wire            n11314;
wire            n11315;
wire            n11316;
wire            n11317;
wire            n11318;
wire            n11319;
wire            n1132;
wire            n11320;
wire            n11321;
wire            n11322;
wire            n11323;
wire            n11324;
wire            n11325;
wire            n11326;
wire            n11327;
wire            n11328;
wire            n11329;
wire            n1133;
wire            n11330;
wire            n11331;
wire            n11332;
wire            n11333;
wire            n11334;
wire            n11335;
wire            n11336;
wire            n11337;
wire            n11338;
wire            n11339;
wire            n1134;
wire            n11340;
wire            n11341;
wire            n11342;
wire            n11343;
wire            n11344;
wire            n11345;
wire            n11346;
wire            n11347;
wire            n11348;
wire            n11349;
wire            n1135;
wire            n11350;
wire            n11351;
wire            n11352;
wire            n11353;
wire            n11354;
wire            n11355;
wire            n11356;
wire            n11357;
wire            n11358;
wire            n11359;
wire            n1136;
wire            n11360;
wire            n11361;
wire            n11362;
wire            n11363;
wire            n11364;
wire            n11365;
wire            n11366;
wire            n11367;
wire            n11368;
wire            n11369;
wire            n1137;
wire            n11370;
wire            n11371;
wire            n11372;
wire            n11373;
wire            n11374;
wire            n11375;
wire            n11376;
wire            n11377;
wire            n11378;
wire            n11379;
wire            n1138;
wire            n11380;
wire            n11381;
wire            n11382;
wire            n11383;
wire            n11384;
wire            n11385;
wire            n11386;
wire            n11387;
wire            n11388;
wire            n11389;
wire            n1139;
wire            n11390;
wire            n11391;
wire            n11392;
wire            n11393;
wire            n11394;
wire            n11395;
wire            n11396;
wire            n11397;
wire            n11398;
wire            n11399;
wire            n114;
wire            n1140;
wire            n11400;
wire            n11401;
wire            n11402;
wire            n11403;
wire            n11404;
wire            n11405;
wire            n11406;
wire            n11407;
wire            n11408;
wire            n11409;
wire            n1141;
wire            n11410;
wire            n11411;
wire            n11412;
wire            n11413;
wire            n11414;
wire            n11415;
wire            n11416;
wire            n11417;
wire            n11418;
wire            n11419;
wire            n1142;
wire            n11420;
wire            n11421;
wire            n11422;
wire            n11423;
wire            n11424;
wire            n11425;
wire            n11426;
wire            n11427;
wire            n11428;
wire            n11429;
wire            n1143;
wire            n11430;
wire            n11431;
wire            n11432;
wire            n11433;
wire            n11434;
wire            n11435;
wire            n11436;
wire            n11437;
wire            n11438;
wire            n11439;
wire            n1144;
wire            n11440;
wire            n11441;
wire            n11442;
wire            n11443;
wire            n11444;
wire            n11445;
wire            n11446;
wire            n11447;
wire            n11448;
wire            n11449;
wire            n1145;
wire            n11450;
wire            n11451;
wire            n11452;
wire            n11453;
wire            n11454;
wire            n11455;
wire            n11456;
wire            n11457;
wire            n11458;
wire            n11459;
wire            n1146;
wire            n11460;
wire            n11461;
wire            n11462;
wire            n11463;
wire            n11464;
wire            n11465;
wire            n11466;
wire            n11467;
wire            n11468;
wire            n11469;
wire            n1147;
wire            n11470;
wire            n11471;
wire            n11472;
wire            n11473;
wire            n11474;
wire            n11475;
wire            n11476;
wire            n11477;
wire            n11478;
wire            n11479;
wire            n1148;
wire            n11480;
wire            n11481;
wire            n11482;
wire            n11483;
wire            n11484;
wire            n11485;
wire            n11486;
wire            n11487;
wire            n11488;
wire            n11489;
wire            n1149;
wire            n11490;
wire            n11491;
wire            n11492;
wire            n11493;
wire            n11494;
wire            n11495;
wire            n11496;
wire            n11497;
wire            n11498;
wire            n11499;
wire            n115;
wire            n1150;
wire            n11500;
wire            n11501;
wire            n11502;
wire            n11503;
wire            n11504;
wire            n11505;
wire            n11506;
wire            n11507;
wire            n11508;
wire            n11509;
wire            n1151;
wire            n11510;
wire            n11511;
wire            n11512;
wire            n11513;
wire            n11514;
wire            n11515;
wire            n11516;
wire            n11517;
wire            n11518;
wire            n11519;
wire            n1152;
wire            n11520;
wire            n11521;
wire            n11522;
wire            n11523;
wire            n11524;
wire            n11525;
wire            n11526;
wire            n11527;
wire            n11528;
wire            n11529;
wire            n1153;
wire            n11530;
wire            n11531;
wire            n11532;
wire            n11533;
wire            n11534;
wire            n11535;
wire            n11536;
wire            n11537;
wire            n11538;
wire            n11539;
wire            n1154;
wire            n11540;
wire            n11541;
wire            n11542;
wire            n11543;
wire            n11544;
wire            n11545;
wire            n11546;
wire            n11547;
wire            n11548;
wire            n11549;
wire            n1155;
wire            n11550;
wire            n11551;
wire            n11552;
wire            n11553;
wire            n11554;
wire            n11555;
wire            n11556;
wire            n11557;
wire            n11558;
wire            n11559;
wire            n1156;
wire            n11560;
wire            n11561;
wire            n11562;
wire            n11563;
wire            n11564;
wire            n11565;
wire            n11566;
wire            n11567;
wire            n11568;
wire            n11569;
wire            n1157;
wire            n11570;
wire            n11571;
wire            n11572;
wire            n11573;
wire            n11574;
wire            n11575;
wire            n11576;
wire            n11577;
wire            n11578;
wire            n11579;
wire            n1158;
wire            n11580;
wire            n11581;
wire            n11582;
wire            n11583;
wire            n11584;
wire            n11585;
wire            n11586;
wire            n11587;
wire            n11588;
wire            n11589;
wire            n1159;
wire            n11590;
wire            n11591;
wire            n11592;
wire            n11593;
wire            n11594;
wire            n11595;
wire            n11596;
wire            n11597;
wire            n11598;
wire            n11599;
wire            n116;
wire            n1160;
wire            n11600;
wire            n11601;
wire            n11602;
wire            n11603;
wire            n11604;
wire            n11605;
wire            n11606;
wire            n11607;
wire            n11608;
wire            n11609;
wire            n1161;
wire            n11610;
wire            n11611;
wire            n11612;
wire            n11613;
wire            n11614;
wire            n11615;
wire            n11616;
wire            n11617;
wire            n11618;
wire            n11619;
wire            n1162;
wire            n11620;
wire            n11621;
wire            n11622;
wire            n11623;
wire            n11624;
wire            n11625;
wire            n11626;
wire            n11627;
wire            n11628;
wire            n11629;
wire            n1163;
wire            n11630;
wire            n11631;
wire            n11632;
wire            n11633;
wire            n11634;
wire            n11635;
wire            n11636;
wire            n11637;
wire            n11638;
wire            n11639;
wire            n1164;
wire            n11640;
wire            n11641;
wire            n11642;
wire            n11643;
wire            n11644;
wire            n11645;
wire            n11646;
wire            n11647;
wire            n11648;
wire            n11649;
wire            n1165;
wire            n11650;
wire            n11651;
wire            n11652;
wire            n11653;
wire            n11654;
wire            n11655;
wire            n11656;
wire            n11657;
wire            n11658;
wire            n11659;
wire            n1166;
wire            n11660;
wire            n11661;
wire            n11662;
wire            n11663;
wire            n11664;
wire            n11665;
wire            n11666;
wire            n11667;
wire            n11668;
wire            n11669;
wire            n1167;
wire            n11670;
wire            n11671;
wire            n11672;
wire            n11673;
wire            n11674;
wire            n11675;
wire            n11676;
wire            n11677;
wire            n11678;
wire            n11679;
wire            n1168;
wire            n11680;
wire            n11681;
wire            n11682;
wire            n11683;
wire            n11684;
wire            n11685;
wire            n11686;
wire            n11687;
wire            n11688;
wire            n11689;
wire            n1169;
wire            n11690;
wire            n11691;
wire            n11692;
wire            n11693;
wire            n11694;
wire            n11695;
wire            n11696;
wire            n11697;
wire            n11698;
wire            n11699;
wire            n117;
wire            n1170;
wire            n11700;
wire            n11701;
wire            n11702;
wire            n11703;
wire            n11704;
wire            n11705;
wire            n11706;
wire            n11707;
wire            n11708;
wire            n11709;
wire            n1171;
wire            n11710;
wire            n11711;
wire            n11712;
wire            n11713;
wire            n11714;
wire            n11715;
wire            n11716;
wire            n11717;
wire            n11718;
wire            n11719;
wire            n1172;
wire            n11720;
wire            n11721;
wire            n11722;
wire            n11723;
wire            n11724;
wire            n11725;
wire            n11726;
wire            n11727;
wire            n11728;
wire            n11729;
wire            n1173;
wire            n11730;
wire            n11731;
wire            n11732;
wire            n11733;
wire            n11734;
wire            n11735;
wire            n11736;
wire            n11737;
wire            n11738;
wire            n11739;
wire            n1174;
wire            n11740;
wire            n11741;
wire            n11742;
wire            n11743;
wire            n11744;
wire            n11745;
wire            n11746;
wire            n11747;
wire            n11748;
wire            n11749;
wire            n1175;
wire            n11750;
wire            n11751;
wire            n11752;
wire            n11753;
wire            n11754;
wire            n11755;
wire            n11756;
wire            n11757;
wire            n11758;
wire            n11759;
wire            n1176;
wire            n11760;
wire            n11761;
wire            n11762;
wire            n11763;
wire            n11764;
wire            n11765;
wire            n11766;
wire            n11767;
wire            n11768;
wire            n11769;
wire            n1177;
wire            n11770;
wire            n11771;
wire            n11772;
wire            n11773;
wire            n11774;
wire            n11775;
wire            n11776;
wire            n11777;
wire            n11778;
wire            n11779;
wire            n1178;
wire            n11780;
wire            n11781;
wire            n11782;
wire            n11783;
wire            n11784;
wire            n11785;
wire            n11786;
wire            n11787;
wire            n11788;
wire            n11789;
wire            n1179;
wire            n11790;
wire            n11791;
wire            n11792;
wire            n11793;
wire            n11794;
wire            n11795;
wire            n11796;
wire            n11797;
wire            n11798;
wire            n11799;
wire            n118;
wire            n1180;
wire            n11800;
wire            n11801;
wire            n11802;
wire            n11803;
wire            n11804;
wire            n11805;
wire            n11806;
wire            n11807;
wire            n11808;
wire            n11809;
wire            n1181;
wire            n11810;
wire            n11811;
wire            n11812;
wire            n11813;
wire            n11814;
wire            n11815;
wire            n11816;
wire            n11817;
wire            n11818;
wire            n11819;
wire            n1182;
wire            n11820;
wire            n11821;
wire            n11822;
wire            n11823;
wire            n11824;
wire            n11825;
wire            n11826;
wire            n11827;
wire            n11828;
wire            n11829;
wire            n1183;
wire            n11830;
wire            n11831;
wire            n11832;
wire            n11833;
wire            n11834;
wire            n11835;
wire            n11836;
wire            n11837;
wire            n11838;
wire            n11839;
wire            n1184;
wire            n11840;
wire            n11841;
wire            n11842;
wire            n11843;
wire            n11844;
wire            n11845;
wire            n11846;
wire            n11847;
wire            n11848;
wire            n11849;
wire            n1185;
wire            n11850;
wire            n11851;
wire            n11852;
wire            n11853;
wire            n11854;
wire            n11855;
wire            n11856;
wire            n11857;
wire            n11858;
wire            n11859;
wire            n1186;
wire            n11860;
wire            n11861;
wire            n11862;
wire            n11863;
wire            n11864;
wire            n11865;
wire            n11866;
wire            n11867;
wire            n11868;
wire            n11869;
wire            n1187;
wire            n11870;
wire            n11871;
wire            n11872;
wire            n11873;
wire            n11874;
wire            n11875;
wire            n11876;
wire            n11877;
wire            n11878;
wire            n11879;
wire            n1188;
wire            n11880;
wire            n11881;
wire            n11882;
wire            n11883;
wire            n11884;
wire            n11885;
wire            n11886;
wire            n11887;
wire            n11888;
wire            n11889;
wire            n1189;
wire            n11890;
wire            n11891;
wire            n11892;
wire            n11893;
wire            n11894;
wire            n11895;
wire            n11896;
wire            n11897;
wire            n11898;
wire            n11899;
wire            n119;
wire            n1190;
wire            n11900;
wire            n11901;
wire            n11902;
wire            n11903;
wire            n11904;
wire            n11905;
wire            n11906;
wire            n11907;
wire            n11908;
wire            n11909;
wire            n1191;
wire            n11910;
wire            n11911;
wire            n11912;
wire            n11913;
wire            n11914;
wire            n11915;
wire            n11916;
wire            n11917;
wire            n11918;
wire            n11919;
wire            n1192;
wire            n11920;
wire            n11921;
wire            n11922;
wire            n11923;
wire            n11924;
wire            n11925;
wire            n11926;
wire            n11927;
wire            n11928;
wire            n11929;
wire            n1193;
wire            n11930;
wire            n11931;
wire            n11932;
wire            n11933;
wire            n11934;
wire            n11935;
wire            n11936;
wire            n11937;
wire            n11938;
wire            n11939;
wire            n1194;
wire            n11940;
wire            n11941;
wire            n11942;
wire            n11943;
wire            n11944;
wire            n11945;
wire            n11946;
wire            n11947;
wire            n11948;
wire            n11949;
wire            n1195;
wire            n11950;
wire            n11951;
wire            n11952;
wire            n11953;
wire            n11954;
wire            n11955;
wire            n11956;
wire            n11957;
wire            n11958;
wire            n11959;
wire            n1196;
wire            n11960;
wire            n11961;
wire            n11962;
wire            n11963;
wire            n11964;
wire            n11965;
wire            n11966;
wire            n11967;
wire            n11968;
wire            n11969;
wire            n1197;
wire            n11970;
wire            n11971;
wire            n11972;
wire            n11973;
wire            n11974;
wire            n11975;
wire            n11976;
wire            n11977;
wire            n11978;
wire            n11979;
wire            n1198;
wire            n11980;
wire            n11981;
wire            n11982;
wire            n11983;
wire            n11984;
wire            n11985;
wire            n11986;
wire            n11987;
wire            n11988;
wire            n11989;
wire            n1199;
wire            n11990;
wire            n11991;
wire            n11992;
wire            n11993;
wire            n11994;
wire            n11995;
wire            n11996;
wire            n11997;
wire            n11998;
wire            n11999;
wire            n12;
wire            n120;
wire            n1200;
wire            n12000;
wire            n12001;
wire            n12002;
wire            n12003;
wire            n12004;
wire            n12005;
wire            n12006;
wire            n12007;
wire            n12008;
wire            n12009;
wire            n1201;
wire            n12010;
wire            n12011;
wire            n12012;
wire            n12013;
wire            n12014;
wire            n12015;
wire            n12016;
wire            n12017;
wire            n12018;
wire            n12019;
wire            n1202;
wire            n12020;
wire            n12021;
wire            n12022;
wire            n12023;
wire            n12024;
wire            n12025;
wire            n12026;
wire            n12027;
wire            n12028;
wire            n12029;
wire            n1203;
wire            n12030;
wire            n12031;
wire            n12032;
wire            n12033;
wire            n12034;
wire            n12035;
wire            n12036;
wire            n12037;
wire            n12038;
wire            n12039;
wire            n1204;
wire            n12040;
wire            n12041;
wire            n12042;
wire            n12043;
wire            n12044;
wire            n12045;
wire            n12046;
wire            n12047;
wire            n12048;
wire            n12049;
wire            n1205;
wire            n12050;
wire            n12051;
wire            n12052;
wire            n12053;
wire            n12054;
wire            n12055;
wire            n12056;
wire            n12057;
wire            n12058;
wire            n12059;
wire            n1206;
wire            n12060;
wire            n12061;
wire            n12062;
wire            n12063;
wire            n12064;
wire            n12065;
wire            n12066;
wire            n12067;
wire            n12068;
wire            n12069;
wire            n1207;
wire            n12070;
wire            n12071;
wire            n12072;
wire            n12073;
wire            n12074;
wire            n12075;
wire            n12076;
wire            n12077;
wire            n12078;
wire            n12079;
wire            n1208;
wire            n12080;
wire            n12081;
wire            n12082;
wire            n12083;
wire            n12084;
wire            n12085;
wire            n12086;
wire            n12087;
wire            n12088;
wire            n12089;
wire            n1209;
wire            n12090;
wire            n12091;
wire            n12092;
wire            n12093;
wire            n12094;
wire            n12095;
wire            n12096;
wire            n12097;
wire            n12098;
wire            n12099;
wire            n121;
wire            n1210;
wire            n12100;
wire            n12101;
wire            n12102;
wire            n12103;
wire            n12104;
wire            n12105;
wire            n12106;
wire            n12107;
wire            n12108;
wire            n12109;
wire            n1211;
wire            n12110;
wire            n12111;
wire            n12112;
wire            n12113;
wire            n12114;
wire            n12115;
wire            n12116;
wire            n12117;
wire            n12118;
wire            n12119;
wire            n1212;
wire            n12120;
wire            n12121;
wire            n12122;
wire            n12123;
wire            n12124;
wire            n12125;
wire            n12126;
wire            n12127;
wire            n12128;
wire            n12129;
wire            n1213;
wire            n12130;
wire            n12131;
wire            n12132;
wire            n12133;
wire            n12134;
wire            n12135;
wire            n12136;
wire            n12137;
wire            n12138;
wire            n12139;
wire            n1214;
wire            n12140;
wire            n12141;
wire            n12142;
wire            n12143;
wire            n12144;
wire            n12145;
wire            n12146;
wire            n12147;
wire            n12148;
wire            n12149;
wire            n1215;
wire            n12150;
wire            n12151;
wire            n12152;
wire            n12153;
wire            n12154;
wire            n12155;
wire            n12156;
wire            n12157;
wire            n12158;
wire            n12159;
wire            n1216;
wire            n12160;
wire            n12161;
wire            n12162;
wire            n12163;
wire            n12164;
wire            n12165;
wire            n12166;
wire            n12167;
wire            n12168;
wire            n12169;
wire            n1217;
wire            n12170;
wire            n12171;
wire            n12172;
wire            n12173;
wire            n12174;
wire            n12175;
wire            n12176;
wire            n12177;
wire            n12178;
wire            n12179;
wire            n1218;
wire            n12180;
wire            n12181;
wire            n12182;
wire            n12183;
wire            n12184;
wire            n12185;
wire            n12186;
wire            n12187;
wire            n12188;
wire            n12189;
wire            n1219;
wire            n12190;
wire            n12191;
wire            n12192;
wire            n12193;
wire            n12194;
wire            n12195;
wire            n12196;
wire            n12197;
wire            n12198;
wire            n12199;
wire            n122;
wire            n1220;
wire            n12200;
wire            n12201;
wire            n12202;
wire            n12203;
wire            n12204;
wire            n12205;
wire            n12206;
wire            n12207;
wire            n12208;
wire            n12209;
wire            n1221;
wire            n12210;
wire            n12211;
wire            n12212;
wire            n12213;
wire            n12214;
wire            n12215;
wire            n12216;
wire            n12217;
wire            n12218;
wire            n12219;
wire            n1222;
wire            n12220;
wire            n12221;
wire            n12222;
wire            n12223;
wire            n12224;
wire            n12225;
wire            n12226;
wire            n12227;
wire            n12228;
wire            n12229;
wire            n1223;
wire            n12230;
wire            n12231;
wire            n12232;
wire            n12233;
wire            n12234;
wire            n12235;
wire            n12236;
wire            n12237;
wire            n12238;
wire            n12239;
wire            n1224;
wire            n12240;
wire            n12241;
wire            n12242;
wire            n12243;
wire            n12244;
wire            n12245;
wire            n12246;
wire            n12247;
wire            n12248;
wire            n12249;
wire            n1225;
wire            n12250;
wire            n12251;
wire            n12252;
wire            n12253;
wire            n12254;
wire            n12255;
wire            n12256;
wire            n12257;
wire            n12258;
wire            n12259;
wire            n1226;
wire            n12260;
wire            n12261;
wire            n12262;
wire            n12263;
wire            n12264;
wire            n12265;
wire            n12266;
wire            n12267;
wire            n12268;
wire            n12269;
wire            n1227;
wire            n12270;
wire            n12271;
wire            n12272;
wire            n12273;
wire            n12274;
wire            n12275;
wire            n12276;
wire            n12277;
wire            n12278;
wire            n12279;
wire            n1228;
wire            n12280;
wire            n12281;
wire            n12282;
wire            n12283;
wire            n12284;
wire            n12285;
wire            n12286;
wire            n12287;
wire            n12288;
wire            n12289;
wire            n1229;
wire            n12290;
wire            n12291;
wire            n12292;
wire            n12293;
wire            n12294;
wire            n12295;
wire            n12296;
wire            n12297;
wire            n12298;
wire            n12299;
wire            n123;
wire            n1230;
wire            n12300;
wire            n12301;
wire            n12302;
wire            n12303;
wire            n12304;
wire            n12305;
wire            n12306;
wire            n12307;
wire            n12308;
wire            n12309;
wire            n1231;
wire            n12310;
wire            n12311;
wire            n12312;
wire            n12313;
wire            n12314;
wire            n12315;
wire            n12316;
wire            n12317;
wire            n12318;
wire            n12319;
wire            n1232;
wire            n12320;
wire            n12321;
wire            n12322;
wire            n12323;
wire            n12324;
wire            n12325;
wire            n12326;
wire            n12327;
wire            n12328;
wire            n12329;
wire            n1233;
wire            n12330;
wire            n12331;
wire            n12332;
wire            n12333;
wire            n12334;
wire            n12335;
wire            n12336;
wire            n12337;
wire            n12338;
wire            n12339;
wire            n1234;
wire            n12340;
wire            n12341;
wire            n12342;
wire            n12343;
wire            n12344;
wire            n12345;
wire            n12346;
wire            n12347;
wire            n12348;
wire            n12349;
wire            n1235;
wire            n12350;
wire            n12351;
wire            n12352;
wire            n12353;
wire            n12354;
wire            n12355;
wire            n12356;
wire            n12357;
wire            n12358;
wire            n12359;
wire            n1236;
wire            n12360;
wire            n12361;
wire            n12362;
wire            n12363;
wire            n12364;
wire            n12365;
wire            n12366;
wire            n12367;
wire            n12368;
wire            n12369;
wire            n1237;
wire            n12370;
wire            n12371;
wire            n12372;
wire            n12373;
wire            n12374;
wire            n12375;
wire            n12376;
wire            n12377;
wire            n12378;
wire            n12379;
wire            n1238;
wire            n12380;
wire            n12381;
wire            n12382;
wire            n12383;
wire            n12384;
wire            n12385;
wire            n12386;
wire            n12387;
wire            n12388;
wire            n12389;
wire            n1239;
wire            n12390;
wire            n12391;
wire            n12392;
wire            n12393;
wire            n12394;
wire            n12395;
wire            n12396;
wire            n12397;
wire            n12398;
wire            n12399;
wire            n124;
wire            n1240;
wire            n12400;
wire            n12401;
wire            n12402;
wire            n12403;
wire            n12404;
wire            n12405;
wire            n12406;
wire            n12407;
wire            n12408;
wire            n12409;
wire            n1241;
wire            n12410;
wire            n12411;
wire            n12412;
wire            n12413;
wire            n12414;
wire            n12415;
wire            n12416;
wire            n12417;
wire            n12418;
wire            n12419;
wire            n1242;
wire            n12420;
wire            n12421;
wire            n12422;
wire            n12423;
wire            n12424;
wire            n12425;
wire            n12426;
wire            n12427;
wire            n12428;
wire            n12429;
wire            n1243;
wire            n12430;
wire            n12431;
wire            n12432;
wire            n12433;
wire            n12434;
wire            n12435;
wire            n12436;
wire            n12437;
wire            n12438;
wire            n12439;
wire            n1244;
wire            n12440;
wire            n12441;
wire            n12442;
wire            n12443;
wire            n12444;
wire            n12445;
wire            n12446;
wire            n12447;
wire            n12448;
wire            n12449;
wire            n1245;
wire            n12450;
wire            n12451;
wire            n12452;
wire            n12453;
wire            n12454;
wire            n12455;
wire            n12456;
wire            n12457;
wire            n12458;
wire            n12459;
wire            n1246;
wire            n12460;
wire            n12461;
wire            n12462;
wire            n12463;
wire            n12464;
wire            n12465;
wire            n12466;
wire            n12467;
wire            n12468;
wire            n12469;
wire            n1247;
wire            n12470;
wire            n12471;
wire            n12472;
wire            n12473;
wire            n12474;
wire            n12475;
wire            n12476;
wire            n12477;
wire            n12478;
wire            n12479;
wire            n1248;
wire            n12480;
wire            n12481;
wire            n12482;
wire            n12483;
wire            n12484;
wire            n12485;
wire            n12486;
wire            n12487;
wire            n12488;
wire            n12489;
wire            n1249;
wire            n12490;
wire            n12491;
wire            n12492;
wire            n12493;
wire            n12494;
wire            n12495;
wire            n12496;
wire            n12497;
wire            n12498;
wire            n12499;
wire            n125;
wire            n1250;
wire            n12500;
wire            n12501;
wire            n12502;
wire            n12503;
wire            n12504;
wire            n12505;
wire            n12506;
wire            n12507;
wire            n12508;
wire            n12509;
wire            n1251;
wire            n12510;
wire            n12511;
wire            n12512;
wire            n12513;
wire            n12514;
wire            n12515;
wire            n12516;
wire            n12517;
wire            n12518;
wire            n12519;
wire            n1252;
wire            n12520;
wire            n12521;
wire            n12522;
wire            n12523;
wire            n12524;
wire            n12525;
wire            n12526;
wire            n12527;
wire            n12528;
wire            n12529;
wire            n1253;
wire            n12530;
wire            n12531;
wire            n12532;
wire            n12533;
wire            n12534;
wire            n12535;
wire            n12536;
wire            n12537;
wire            n12538;
wire            n12539;
wire            n1254;
wire            n12540;
wire            n12541;
wire            n12542;
wire            n12543;
wire            n12544;
wire            n12545;
wire            n12546;
wire            n12547;
wire            n12548;
wire            n12549;
wire            n1255;
wire            n12550;
wire            n12551;
wire            n12552;
wire            n12553;
wire            n12554;
wire            n12555;
wire            n12556;
wire            n12557;
wire            n12558;
wire            n12559;
wire            n1256;
wire            n12560;
wire            n12561;
wire            n12562;
wire            n12563;
wire            n12564;
wire            n12565;
wire            n12566;
wire            n12567;
wire            n12568;
wire            n12569;
wire            n1257;
wire            n12570;
wire            n12571;
wire            n12572;
wire            n12573;
wire            n12574;
wire            n12575;
wire            n12576;
wire            n12577;
wire            n12578;
wire            n12579;
wire            n1258;
wire            n12580;
wire            n12581;
wire            n12582;
wire            n12583;
wire            n12584;
wire            n12585;
wire            n12586;
wire            n12587;
wire            n12588;
wire            n12589;
wire            n1259;
wire            n12590;
wire            n12591;
wire            n12592;
wire            n12593;
wire            n12594;
wire            n12595;
wire            n12596;
wire            n12597;
wire            n12598;
wire            n12599;
wire            n126;
wire            n1260;
wire            n12600;
wire            n12601;
wire            n12602;
wire            n12603;
wire            n12604;
wire            n12605;
wire            n12606;
wire            n12607;
wire            n12608;
wire            n12609;
wire            n1261;
wire            n12610;
wire            n12611;
wire            n12612;
wire            n12613;
wire            n12614;
wire            n12615;
wire            n12616;
wire            n12617;
wire            n12618;
wire            n12619;
wire            n1262;
wire            n12620;
wire            n12621;
wire            n12622;
wire            n12623;
wire            n12624;
wire            n12625;
wire            n12626;
wire            n12627;
wire            n12628;
wire            n12629;
wire            n1263;
wire            n12630;
wire            n12631;
wire            n12632;
wire            n12633;
wire            n12634;
wire            n12635;
wire            n12636;
wire            n12637;
wire            n12638;
wire            n12639;
wire            n1264;
wire            n12640;
wire            n12641;
wire            n12642;
wire            n12643;
wire            n12644;
wire            n12645;
wire            n12646;
wire            n12647;
wire            n12648;
wire            n12649;
wire            n1265;
wire            n12650;
wire            n12651;
wire            n12652;
wire            n12653;
wire            n12654;
wire            n12655;
wire            n12656;
wire            n12657;
wire            n12658;
wire            n12659;
wire            n1266;
wire            n12660;
wire            n12661;
wire            n12662;
wire            n12663;
wire            n12664;
wire            n12665;
wire            n12666;
wire            n12667;
wire            n12668;
wire            n12669;
wire            n1267;
wire            n12670;
wire            n12671;
wire            n12672;
wire            n12673;
wire            n12674;
wire            n12675;
wire            n12676;
wire            n12677;
wire            n12678;
wire            n12679;
wire            n1268;
wire            n12680;
wire            n12681;
wire            n12682;
wire            n12683;
wire            n12684;
wire            n12685;
wire            n12686;
wire            n12687;
wire            n12688;
wire            n12689;
wire            n1269;
wire            n12690;
wire            n12691;
wire            n12692;
wire            n12693;
wire            n12694;
wire            n12695;
wire            n12696;
wire            n12697;
wire            n12698;
wire            n12699;
wire            n127;
wire            n1270;
wire            n12700;
wire            n12701;
wire            n12702;
wire            n12703;
wire            n12704;
wire            n12705;
wire            n12706;
wire            n12707;
wire            n12708;
wire            n12709;
wire            n1271;
wire            n12710;
wire            n12711;
wire            n12712;
wire            n12713;
wire            n12714;
wire            n12715;
wire            n12716;
wire            n12717;
wire            n12718;
wire            n12719;
wire            n1272;
wire            n12720;
wire            n12721;
wire            n12722;
wire            n12723;
wire            n12724;
wire            n12725;
wire            n12726;
wire            n12727;
wire            n12728;
wire            n12729;
wire            n1273;
wire            n12730;
wire            n12731;
wire            n12732;
wire            n12733;
wire            n12734;
wire            n12735;
wire            n12736;
wire            n12737;
wire            n12738;
wire            n12739;
wire            n1274;
wire            n12740;
wire            n12741;
wire            n12742;
wire            n12743;
wire            n12744;
wire            n12745;
wire            n12746;
wire            n12747;
wire            n12748;
wire            n12749;
wire            n1275;
wire            n12750;
wire            n12751;
wire            n12752;
wire            n12753;
wire            n12754;
wire            n12755;
wire            n12756;
wire            n12757;
wire            n12758;
wire            n12759;
wire            n1276;
wire            n12760;
wire            n12761;
wire            n12762;
wire            n12763;
wire            n12764;
wire            n12765;
wire            n12766;
wire            n12767;
wire            n12768;
wire            n12769;
wire            n1277;
wire            n12770;
wire            n12771;
wire            n12772;
wire            n12773;
wire            n12774;
wire            n12775;
wire            n12776;
wire            n12777;
wire            n12778;
wire            n12779;
wire            n1278;
wire            n12780;
wire            n12781;
wire            n12782;
wire            n12783;
wire            n12784;
wire            n12785;
wire            n12786;
wire            n12787;
wire            n12788;
wire            n12789;
wire            n1279;
wire            n12790;
wire            n12791;
wire            n12792;
wire            n12793;
wire            n12794;
wire            n12795;
wire            n12796;
wire            n12797;
wire            n12798;
wire            n12799;
wire            n128;
wire            n1280;
wire            n12800;
wire            n12801;
wire            n12802;
wire            n12803;
wire            n12804;
wire            n12805;
wire            n12806;
wire            n12807;
wire            n12808;
wire            n12809;
wire            n1281;
wire            n12810;
wire            n12811;
wire            n12812;
wire            n12813;
wire            n12814;
wire            n12815;
wire            n12816;
wire            n12817;
wire            n12818;
wire            n12819;
wire            n1282;
wire            n12820;
wire            n12821;
wire            n12822;
wire            n12823;
wire            n12824;
wire            n12825;
wire            n12826;
wire            n12827;
wire            n12828;
wire            n12829;
wire            n1283;
wire            n12830;
wire            n12831;
wire            n12832;
wire            n12833;
wire            n12834;
wire            n12835;
wire            n12836;
wire            n12837;
wire            n12838;
wire            n12839;
wire            n1284;
wire            n12840;
wire            n12841;
wire            n12842;
wire            n12843;
wire            n12844;
wire            n12845;
wire            n12846;
wire            n12847;
wire            n12848;
wire            n12849;
wire            n1285;
wire            n12850;
wire            n12851;
wire            n12852;
wire            n12853;
wire            n12854;
wire            n12855;
wire            n12856;
wire            n12857;
wire            n12858;
wire            n12859;
wire            n1286;
wire            n12860;
wire            n12861;
wire            n12862;
wire            n12863;
wire            n12864;
wire            n12865;
wire            n12866;
wire            n12867;
wire            n12868;
wire            n12869;
wire            n1287;
wire            n12870;
wire            n12871;
wire            n12872;
wire            n12873;
wire            n12874;
wire            n12875;
wire            n12876;
wire            n12877;
wire            n12878;
wire            n12879;
wire            n1288;
wire            n12880;
wire            n12881;
wire            n12882;
wire            n12883;
wire            n12884;
wire            n12885;
wire            n12886;
wire            n12887;
wire            n12888;
wire            n12889;
wire            n1289;
wire            n12890;
wire            n12891;
wire            n12892;
wire            n12893;
wire            n12894;
wire            n12895;
wire            n12896;
wire            n12897;
wire            n12898;
wire            n12899;
wire            n129;
wire            n1290;
wire            n12900;
wire            n12901;
wire            n12902;
wire            n12903;
wire            n12904;
wire            n12905;
wire            n12906;
wire            n12907;
wire            n12908;
wire            n12909;
wire            n1291;
wire            n12910;
wire            n12911;
wire            n12912;
wire            n12913;
wire            n12914;
wire            n12915;
wire            n12916;
wire            n12917;
wire            n12918;
wire            n12919;
wire            n1292;
wire            n12920;
wire            n12921;
wire            n12922;
wire            n12923;
wire            n12924;
wire            n12925;
wire            n12926;
wire            n12927;
wire            n12928;
wire            n12929;
wire            n1293;
wire            n12930;
wire            n12931;
wire            n12932;
wire            n12933;
wire            n12934;
wire            n12935;
wire            n12936;
wire            n12937;
wire            n12938;
wire            n12939;
wire            n1294;
wire            n12940;
wire            n12941;
wire            n12942;
wire            n12943;
wire            n12944;
wire            n12945;
wire            n12946;
wire            n12947;
wire            n12948;
wire            n12949;
wire            n1295;
wire            n12950;
wire            n12951;
wire            n12952;
wire            n12953;
wire            n12954;
wire            n12955;
wire            n12956;
wire            n12957;
wire            n12958;
wire            n12959;
wire            n1296;
wire            n12960;
wire            n12961;
wire            n12962;
wire            n12963;
wire            n12964;
wire            n12965;
wire            n12966;
wire            n12967;
wire            n12968;
wire            n12969;
wire            n1297;
wire            n12970;
wire            n12971;
wire            n12972;
wire            n12973;
wire            n12974;
wire            n12975;
wire            n12976;
wire            n12977;
wire            n12978;
wire            n12979;
wire            n1298;
wire            n12980;
wire            n12981;
wire            n12982;
wire            n12983;
wire            n12984;
wire            n12985;
wire            n12986;
wire            n12987;
wire            n12988;
wire            n12989;
wire            n1299;
wire            n12990;
wire            n12991;
wire            n12992;
wire            n12993;
wire            n12994;
wire            n12995;
wire            n12996;
wire            n12997;
wire            n12998;
wire            n12999;
wire            n13;
wire            n130;
wire            n1300;
wire            n13000;
wire            n13001;
wire            n13002;
wire            n13003;
wire            n13004;
wire            n13005;
wire            n13006;
wire            n13007;
wire            n13008;
wire            n13009;
wire            n1301;
wire            n13010;
wire            n13011;
wire            n13012;
wire            n13013;
wire            n13014;
wire            n13015;
wire            n13016;
wire            n13017;
wire            n13018;
wire            n13019;
wire            n1302;
wire            n13020;
wire            n13021;
wire            n13022;
wire            n13023;
wire            n13024;
wire            n13025;
wire            n13026;
wire            n13027;
wire            n13028;
wire            n13029;
wire            n1303;
wire            n13030;
wire            n13031;
wire            n13032;
wire            n13033;
wire            n13034;
wire            n13035;
wire            n13036;
wire            n13037;
wire            n13038;
wire            n13039;
wire            n1304;
wire            n13040;
wire            n13041;
wire            n13042;
wire            n13043;
wire            n13044;
wire            n13045;
wire            n13046;
wire            n13047;
wire            n13048;
wire            n13049;
wire            n1305;
wire            n13050;
wire            n13051;
wire            n13052;
wire            n13053;
wire            n13054;
wire            n13055;
wire            n13056;
wire            n13057;
wire            n13058;
wire            n13059;
wire            n1306;
wire            n13060;
wire            n13061;
wire            n13062;
wire            n13063;
wire            n13064;
wire            n13065;
wire            n13066;
wire            n13067;
wire            n13068;
wire            n13069;
wire            n1307;
wire            n13070;
wire            n13071;
wire            n13072;
wire            n13073;
wire            n13074;
wire            n13075;
wire            n13076;
wire            n13077;
wire            n13078;
wire            n13079;
wire            n1308;
wire            n13080;
wire            n13081;
wire            n13082;
wire            n13083;
wire            n13084;
wire            n13085;
wire            n13086;
wire            n13087;
wire            n13088;
wire            n13089;
wire            n1309;
wire            n13090;
wire            n13091;
wire            n13092;
wire            n13093;
wire            n13094;
wire            n13095;
wire            n13096;
wire            n13097;
wire            n13098;
wire            n13099;
wire            n131;
wire            n1310;
wire            n13100;
wire            n13101;
wire            n13102;
wire            n13103;
wire            n13104;
wire            n13105;
wire            n13106;
wire            n13107;
wire            n13108;
wire            n13109;
wire            n1311;
wire            n13110;
wire            n13111;
wire            n13112;
wire            n13113;
wire            n13114;
wire            n13115;
wire            n13116;
wire            n13117;
wire            n13118;
wire            n13119;
wire            n1312;
wire            n13120;
wire            n13121;
wire            n13122;
wire            n13123;
wire            n13124;
wire            n13125;
wire            n13126;
wire            n13127;
wire            n13128;
wire            n13129;
wire            n1313;
wire            n13130;
wire            n13131;
wire            n13132;
wire            n13133;
wire            n13134;
wire            n13135;
wire            n13136;
wire            n13137;
wire            n13138;
wire            n13139;
wire            n1314;
wire            n13140;
wire            n13141;
wire            n13142;
wire            n13143;
wire            n13144;
wire            n13145;
wire            n13146;
wire            n13147;
wire            n13148;
wire            n13149;
wire            n1315;
wire            n13150;
wire            n13151;
wire            n13152;
wire            n13153;
wire            n13154;
wire            n13155;
wire            n13156;
wire            n13157;
wire            n13158;
wire            n13159;
wire            n1316;
wire            n13160;
wire            n13161;
wire            n13162;
wire            n13163;
wire            n13164;
wire            n13165;
wire            n13166;
wire            n13167;
wire            n13168;
wire            n13169;
wire            n1317;
wire            n13170;
wire            n13171;
wire            n13172;
wire            n13173;
wire            n13174;
wire            n13175;
wire            n13176;
wire            n13177;
wire            n13178;
wire            n13179;
wire            n1318;
wire            n13180;
wire            n13181;
wire            n13182;
wire            n13183;
wire            n13184;
wire            n13185;
wire            n13186;
wire            n13187;
wire            n13188;
wire            n13189;
wire            n1319;
wire            n13190;
wire            n13191;
wire            n13192;
wire            n13193;
wire            n13194;
wire            n13195;
wire            n13196;
wire            n13197;
wire            n13198;
wire            n13199;
wire            n132;
wire            n1320;
wire            n13200;
wire            n13201;
wire            n13202;
wire            n13203;
wire            n13204;
wire            n13205;
wire            n13206;
wire            n13207;
wire            n13208;
wire            n13209;
wire            n1321;
wire            n13210;
wire            n13211;
wire            n13212;
wire            n13213;
wire            n13214;
wire            n13215;
wire            n13216;
wire            n13217;
wire            n13218;
wire            n13219;
wire            n1322;
wire            n13220;
wire            n13221;
wire            n13222;
wire            n13223;
wire            n13224;
wire            n13225;
wire            n13226;
wire            n13227;
wire            n13228;
wire            n13229;
wire            n1323;
wire            n13230;
wire            n13231;
wire            n13232;
wire            n13233;
wire            n13234;
wire            n13235;
wire            n13236;
wire            n13237;
wire            n13238;
wire            n13239;
wire            n1324;
wire            n13240;
wire            n13241;
wire            n13242;
wire            n13243;
wire            n13244;
wire            n13245;
wire            n13246;
wire            n13247;
wire            n13248;
wire            n13249;
wire            n1325;
wire            n13250;
wire            n13251;
wire            n13252;
wire            n13253;
wire            n13254;
wire            n13255;
wire            n13256;
wire            n13257;
wire            n13258;
wire            n13259;
wire            n1326;
wire            n13260;
wire            n13261;
wire            n13262;
wire            n13263;
wire            n13264;
wire            n13265;
wire            n13266;
wire            n13267;
wire            n13268;
wire            n13269;
wire            n1327;
wire            n13270;
wire            n13271;
wire            n13272;
wire            n13273;
wire            n13274;
wire            n13275;
wire            n13276;
wire            n13277;
wire            n13278;
wire            n13279;
wire            n1328;
wire            n13280;
wire            n13281;
wire            n13282;
wire            n13283;
wire            n13284;
wire            n13285;
wire            n13286;
wire            n13287;
wire            n13288;
wire            n13289;
wire            n1329;
wire            n13290;
wire            n13291;
wire            n13292;
wire            n13293;
wire            n13294;
wire            n13295;
wire            n13296;
wire            n13297;
wire            n13298;
wire            n13299;
wire            n133;
wire            n1330;
wire            n13300;
wire            n13301;
wire            n13302;
wire            n13303;
wire            n13304;
wire            n13305;
wire            n13306;
wire            n13307;
wire            n13308;
wire            n13309;
wire            n1331;
wire            n13310;
wire            n13311;
wire            n13312;
wire            n13313;
wire            n13314;
wire            n13315;
wire            n13316;
wire            n13317;
wire            n13318;
wire            n13319;
wire            n1332;
wire            n13320;
wire            n13321;
wire            n13322;
wire            n13323;
wire            n13324;
wire            n13325;
wire            n13326;
wire            n13327;
wire            n13328;
wire            n13329;
wire            n1333;
wire            n13330;
wire            n13331;
wire            n13332;
wire            n13333;
wire            n13334;
wire            n13335;
wire            n13336;
wire            n13337;
wire            n13338;
wire            n13339;
wire            n1334;
wire            n13340;
wire            n13341;
wire            n13342;
wire            n13343;
wire            n13344;
wire            n13345;
wire            n13346;
wire            n13347;
wire            n13348;
wire            n13349;
wire            n1335;
wire            n13350;
wire            n13351;
wire            n13352;
wire            n13353;
wire            n13354;
wire            n13355;
wire            n13356;
wire            n13357;
wire            n13358;
wire            n13359;
wire            n1336;
wire            n13360;
wire            n13361;
wire            n13362;
wire            n13363;
wire            n13364;
wire            n13365;
wire            n13366;
wire            n13367;
wire            n13368;
wire            n13369;
wire            n1337;
wire            n13370;
wire            n13371;
wire            n13372;
wire            n13373;
wire            n13374;
wire            n13375;
wire            n13376;
wire            n13377;
wire            n13378;
wire            n13379;
wire            n1338;
wire            n13380;
wire            n13381;
wire            n13382;
wire            n13383;
wire            n13384;
wire            n13385;
wire            n13386;
wire            n13387;
wire            n13388;
wire            n13389;
wire            n1339;
wire            n13390;
wire            n13391;
wire            n13392;
wire            n13393;
wire            n13394;
wire            n13395;
wire            n13396;
wire            n13397;
wire            n13398;
wire            n13399;
wire            n134;
wire            n1340;
wire            n13400;
wire            n13401;
wire            n13402;
wire            n13403;
wire            n13404;
wire            n13405;
wire            n13406;
wire            n13407;
wire            n13408;
wire            n13409;
wire            n1341;
wire            n13410;
wire            n13411;
wire            n13412;
wire            n13413;
wire            n13414;
wire            n13415;
wire            n13416;
wire            n13417;
wire            n13418;
wire            n13419;
wire            n1342;
wire            n13420;
wire            n13421;
wire            n13422;
wire            n13423;
wire            n13424;
wire            n13425;
wire            n13426;
wire            n13427;
wire            n13428;
wire            n13429;
wire            n1343;
wire            n13430;
wire            n13431;
wire            n13432;
wire            n13433;
wire            n13434;
wire            n13435;
wire            n13436;
wire            n13437;
wire            n13438;
wire            n13439;
wire            n1344;
wire            n13440;
wire            n13441;
wire            n13442;
wire            n13443;
wire            n13444;
wire            n13445;
wire            n13446;
wire            n13447;
wire            n13448;
wire            n13449;
wire            n1345;
wire            n13450;
wire            n13451;
wire            n13452;
wire            n13453;
wire            n13454;
wire            n13455;
wire            n13456;
wire            n13457;
wire            n13458;
wire            n13459;
wire            n1346;
wire            n13460;
wire            n13461;
wire            n13462;
wire            n13463;
wire            n13464;
wire            n13465;
wire            n13466;
wire            n13467;
wire            n13468;
wire            n13469;
wire            n1347;
wire            n13470;
wire            n13471;
wire            n13472;
wire            n13473;
wire            n13474;
wire            n13475;
wire            n13476;
wire            n13477;
wire            n13478;
wire            n13479;
wire            n1348;
wire            n13480;
wire            n13481;
wire            n13482;
wire            n13483;
wire            n13484;
wire            n13485;
wire            n13486;
wire            n13487;
wire            n13488;
wire            n13489;
wire            n1349;
wire            n13490;
wire            n13491;
wire            n13492;
wire            n13493;
wire            n13494;
wire            n13495;
wire            n13496;
wire            n13497;
wire            n13498;
wire            n13499;
wire            n135;
wire            n1350;
wire            n13500;
wire            n13501;
wire            n13502;
wire            n13503;
wire            n13504;
wire            n13505;
wire            n13506;
wire            n13507;
wire            n13508;
wire            n13509;
wire            n1351;
wire            n13510;
wire            n13511;
wire            n13512;
wire            n13513;
wire            n13514;
wire            n13515;
wire            n13516;
wire            n13517;
wire            n13518;
wire            n13519;
wire            n1352;
wire            n13520;
wire            n13521;
wire            n13522;
wire            n13523;
wire            n13524;
wire            n13525;
wire            n13526;
wire            n13527;
wire            n13528;
wire            n13529;
wire            n1353;
wire            n13530;
wire            n13531;
wire            n13532;
wire            n13533;
wire            n13534;
wire            n13535;
wire            n13536;
wire            n13537;
wire            n13538;
wire            n13539;
wire            n1354;
wire            n13540;
wire            n13541;
wire            n13542;
wire            n13543;
wire            n13544;
wire            n13545;
wire            n13546;
wire            n13547;
wire            n13548;
wire            n13549;
wire            n1355;
wire            n13550;
wire            n13551;
wire            n13552;
wire            n13553;
wire            n13554;
wire            n13555;
wire            n13556;
wire            n13557;
wire            n13558;
wire            n13559;
wire            n1356;
wire            n13560;
wire            n13561;
wire            n13562;
wire            n13563;
wire            n13564;
wire            n13565;
wire            n13566;
wire            n13567;
wire            n13568;
wire            n13569;
wire            n1357;
wire            n13570;
wire            n13571;
wire            n13572;
wire            n13573;
wire            n13574;
wire            n13575;
wire            n13576;
wire            n13577;
wire            n13578;
wire            n13579;
wire            n1358;
wire            n13580;
wire            n13581;
wire            n13582;
wire            n13583;
wire            n13584;
wire            n13585;
wire            n13586;
wire            n13587;
wire            n13588;
wire            n13589;
wire            n1359;
wire            n13590;
wire            n13591;
wire            n13592;
wire            n13593;
wire            n13594;
wire            n13595;
wire            n13596;
wire            n13597;
wire            n13598;
wire            n13599;
wire            n136;
wire            n1360;
wire            n13600;
wire            n13601;
wire            n13602;
wire            n13603;
wire            n13604;
wire            n13605;
wire            n13606;
wire            n13607;
wire            n13608;
wire            n13609;
wire            n1361;
wire            n13610;
wire            n13611;
wire            n13612;
wire            n13613;
wire            n13614;
wire            n13615;
wire            n13616;
wire            n13617;
wire            n13618;
wire            n13619;
wire            n1362;
wire            n13620;
wire            n13621;
wire            n13622;
wire            n13623;
wire            n13624;
wire            n13625;
wire            n13626;
wire            n13627;
wire            n13628;
wire            n13629;
wire            n1363;
wire            n13630;
wire            n13631;
wire            n13632;
wire            n13633;
wire            n13634;
wire            n13635;
wire            n13636;
wire            n13637;
wire            n13638;
wire            n13639;
wire            n1364;
wire            n13640;
wire            n13641;
wire            n13642;
wire            n13643;
wire            n13644;
wire            n13645;
wire            n13646;
wire            n13647;
wire            n13648;
wire            n13649;
wire            n1365;
wire            n13650;
wire            n13651;
wire            n13652;
wire            n13653;
wire            n13654;
wire            n13655;
wire            n13656;
wire            n13657;
wire            n13658;
wire            n13659;
wire            n1366;
wire            n13660;
wire            n13661;
wire            n13662;
wire            n13663;
wire            n13664;
wire            n13665;
wire            n13666;
wire            n13667;
wire            n13668;
wire            n13669;
wire            n1367;
wire            n13670;
wire            n13671;
wire            n13672;
wire            n13673;
wire            n13674;
wire            n13675;
wire            n13676;
wire            n13677;
wire            n13678;
wire            n13679;
wire            n1368;
wire            n13680;
wire            n13681;
wire            n13682;
wire            n13683;
wire            n13684;
wire            n13685;
wire            n13686;
wire            n13687;
wire            n13688;
wire            n13689;
wire            n1369;
wire            n13690;
wire            n13691;
wire            n13692;
wire            n13693;
wire            n13694;
wire            n13695;
wire            n13696;
wire            n13697;
wire            n13698;
wire            n13699;
wire            n137;
wire            n1370;
wire            n13700;
wire            n13701;
wire            n13702;
wire            n13703;
wire            n13704;
wire            n13705;
wire            n13706;
wire            n13707;
wire            n13708;
wire            n13709;
wire            n1371;
wire            n13710;
wire            n13711;
wire            n13712;
wire            n13713;
wire            n13714;
wire            n13715;
wire            n13716;
wire            n13717;
wire            n13718;
wire            n13719;
wire            n1372;
wire            n13720;
wire            n13721;
wire            n13722;
wire            n13723;
wire            n13724;
wire            n13725;
wire            n13726;
wire            n13727;
wire            n13728;
wire            n13729;
wire            n1373;
wire            n13730;
wire            n13731;
wire            n13732;
wire            n13733;
wire            n13734;
wire            n13735;
wire            n13736;
wire            n13737;
wire            n13738;
wire            n13739;
wire            n1374;
wire            n13740;
wire            n13741;
wire            n13742;
wire            n13743;
wire            n13744;
wire            n13745;
wire            n13746;
wire            n13747;
wire            n13748;
wire            n13749;
wire            n1375;
wire            n13750;
wire            n13751;
wire            n13752;
wire            n13753;
wire            n13754;
wire            n13755;
wire            n13756;
wire            n13757;
wire            n13758;
wire            n13759;
wire            n1376;
wire            n13760;
wire            n13761;
wire            n13762;
wire            n13763;
wire            n13764;
wire            n13765;
wire            n13766;
wire            n13767;
wire            n13768;
wire            n13769;
wire            n1377;
wire            n13770;
wire            n13771;
wire            n13772;
wire            n13773;
wire            n13774;
wire            n13775;
wire            n13776;
wire            n13777;
wire            n13778;
wire            n13779;
wire            n1378;
wire            n13780;
wire            n13781;
wire            n13782;
wire            n13783;
wire            n13784;
wire            n13785;
wire            n13786;
wire            n13787;
wire            n13788;
wire            n13789;
wire            n1379;
wire            n13790;
wire            n13791;
wire            n13792;
wire            n13793;
wire            n13794;
wire            n13795;
wire            n13796;
wire            n13797;
wire            n13798;
wire            n13799;
wire            n138;
wire            n1380;
wire            n13800;
wire            n13801;
wire            n13802;
wire            n13803;
wire            n13804;
wire            n13805;
wire            n13806;
wire            n13807;
wire            n13808;
wire            n13809;
wire            n1381;
wire            n13810;
wire            n13811;
wire            n13812;
wire            n13813;
wire            n13814;
wire            n13815;
wire            n13816;
wire            n13817;
wire            n13818;
wire            n13819;
wire            n1382;
wire            n13820;
wire            n13821;
wire            n13822;
wire            n13823;
wire            n13824;
wire            n13825;
wire            n13826;
wire            n13827;
wire            n13828;
wire            n13829;
wire            n1383;
wire            n13830;
wire            n13831;
wire            n13832;
wire            n13833;
wire            n13834;
wire            n13835;
wire            n13836;
wire            n13837;
wire            n13838;
wire            n13839;
wire            n1384;
wire            n13840;
wire            n13841;
wire            n13842;
wire            n13843;
wire            n13844;
wire            n13845;
wire            n13846;
wire            n13847;
wire            n13848;
wire            n13849;
wire            n1385;
wire            n13850;
wire            n13851;
wire            n13852;
wire            n13853;
wire            n13854;
wire            n13855;
wire            n13856;
wire            n13857;
wire            n13858;
wire            n13859;
wire            n1386;
wire            n13860;
wire            n13861;
wire            n13862;
wire            n13863;
wire            n13864;
wire            n13865;
wire            n13866;
wire            n13867;
wire            n13868;
wire            n13869;
wire            n1387;
wire            n13870;
wire            n13871;
wire            n13872;
wire            n13873;
wire            n13874;
wire            n13875;
wire            n13876;
wire            n13877;
wire            n13878;
wire            n13879;
wire            n1388;
wire            n13880;
wire            n13881;
wire            n13882;
wire            n13883;
wire            n13884;
wire            n13885;
wire            n13886;
wire            n13887;
wire            n13888;
wire            n13889;
wire            n1389;
wire            n13890;
wire            n13891;
wire            n13892;
wire            n13893;
wire            n13894;
wire            n13895;
wire            n13896;
wire            n13897;
wire            n13898;
wire            n13899;
wire            n139;
wire            n1390;
wire            n13900;
wire            n13901;
wire            n13902;
wire            n13903;
wire            n13904;
wire            n13905;
wire            n13906;
wire            n13907;
wire            n13908;
wire            n13909;
wire            n1391;
wire            n13910;
wire            n13911;
wire            n13912;
wire            n13913;
wire            n13914;
wire            n13915;
wire            n13916;
wire            n13917;
wire            n13918;
wire            n13919;
wire            n1392;
wire            n13920;
wire            n13921;
wire            n13922;
wire            n13923;
wire            n13924;
wire            n13925;
wire            n13926;
wire            n13927;
wire            n13928;
wire            n13929;
wire            n1393;
wire            n13930;
wire            n13931;
wire            n13932;
wire            n13933;
wire            n13934;
wire            n13935;
wire            n13936;
wire            n13937;
wire            n13938;
wire            n13939;
wire            n1394;
wire            n13940;
wire            n13941;
wire            n13942;
wire            n13943;
wire            n13944;
wire            n13945;
wire            n13946;
wire            n13947;
wire            n13948;
wire            n13949;
wire            n1395;
wire            n13950;
wire            n13951;
wire            n13952;
wire            n13953;
wire            n13954;
wire            n13955;
wire            n13956;
wire            n13957;
wire            n13958;
wire            n13959;
wire            n1396;
wire            n13960;
wire            n13961;
wire            n13962;
wire            n13963;
wire            n13964;
wire            n13965;
wire            n13966;
wire            n13967;
wire            n13968;
wire            n13969;
wire            n1397;
wire            n13970;
wire            n13971;
wire            n13972;
wire            n13973;
wire            n13974;
wire            n13975;
wire            n13976;
wire            n13977;
wire            n13978;
wire            n13979;
wire            n1398;
wire            n13980;
wire            n13981;
wire            n13982;
wire            n13983;
wire            n13984;
wire            n13985;
wire            n13986;
wire            n13987;
wire            n13988;
wire            n13989;
wire            n1399;
wire            n13990;
wire            n13991;
wire            n13992;
wire            n13993;
wire            n13994;
wire            n13995;
wire            n13996;
wire            n13997;
wire            n13998;
wire            n13999;
wire            n14;
wire            n140;
wire            n1400;
wire            n14000;
wire            n14001;
wire            n14002;
wire            n14003;
wire            n14004;
wire            n14005;
wire            n14006;
wire            n14007;
wire            n14008;
wire            n14009;
wire            n1401;
wire            n14010;
wire            n14011;
wire            n14012;
wire            n14013;
wire            n14014;
wire            n14015;
wire            n14016;
wire            n14017;
wire            n14018;
wire            n14019;
wire            n1402;
wire            n14020;
wire            n14021;
wire            n14022;
wire            n14023;
wire            n14024;
wire            n14025;
wire            n14026;
wire            n14027;
wire            n14028;
wire            n14029;
wire            n1403;
wire            n14030;
wire            n14031;
wire            n14032;
wire            n14033;
wire            n14034;
wire            n14035;
wire            n14036;
wire            n14037;
wire            n14038;
wire            n14039;
wire            n1404;
wire            n14040;
wire            n14041;
wire            n14042;
wire            n14043;
wire            n14044;
wire            n14045;
wire            n14046;
wire            n14047;
wire            n14048;
wire            n14049;
wire            n1405;
wire            n14050;
wire            n14051;
wire            n14052;
wire            n14053;
wire            n14054;
wire            n14055;
wire            n14056;
wire            n14057;
wire            n14058;
wire            n14059;
wire            n1406;
wire            n14060;
wire            n14061;
wire            n14062;
wire            n14063;
wire            n14064;
wire            n14065;
wire            n14066;
wire            n14067;
wire            n14068;
wire            n14069;
wire            n1407;
wire            n14070;
wire            n14071;
wire            n14072;
wire            n14073;
wire            n14074;
wire            n14075;
wire            n14076;
wire            n14077;
wire            n14078;
wire            n14079;
wire            n1408;
wire            n14080;
wire            n14081;
wire            n14082;
wire            n14083;
wire            n14084;
wire            n14085;
wire            n14086;
wire            n14087;
wire            n14088;
wire            n14089;
wire            n1409;
wire            n14090;
wire            n14091;
wire            n14092;
wire            n14093;
wire            n14094;
wire            n14095;
wire            n14096;
wire            n14097;
wire            n14098;
wire            n14099;
wire            n141;
wire            n1410;
wire            n14100;
wire            n14101;
wire            n14102;
wire            n14103;
wire            n14104;
wire            n14105;
wire            n14106;
wire            n14107;
wire            n14108;
wire            n14109;
wire            n1411;
wire            n14110;
wire            n14111;
wire            n14112;
wire            n14113;
wire            n14114;
wire            n14115;
wire            n14116;
wire            n14117;
wire            n14118;
wire            n14119;
wire            n1412;
wire            n14120;
wire            n14121;
wire            n14122;
wire            n14123;
wire            n14124;
wire            n14125;
wire            n14126;
wire            n14127;
wire            n14128;
wire            n14129;
wire            n1413;
wire            n14130;
wire            n14131;
wire            n14132;
wire            n14133;
wire            n14134;
wire            n14135;
wire            n14136;
wire            n14137;
wire            n14138;
wire            n14139;
wire            n1414;
wire            n14140;
wire            n14141;
wire            n14142;
wire            n14143;
wire            n14144;
wire            n14145;
wire            n14146;
wire            n14147;
wire            n14148;
wire            n14149;
wire            n1415;
wire            n14150;
wire            n14151;
wire            n14152;
wire            n14153;
wire            n14154;
wire            n14155;
wire            n14156;
wire            n14157;
wire            n14158;
wire            n14159;
wire            n1416;
wire            n14160;
wire            n14161;
wire            n14162;
wire            n14163;
wire            n14164;
wire            n14165;
wire            n14166;
wire            n14167;
wire            n14168;
wire            n14169;
wire            n1417;
wire            n14170;
wire            n14171;
wire            n14172;
wire            n14173;
wire            n14174;
wire            n14175;
wire            n14176;
wire            n14177;
wire            n14178;
wire            n14179;
wire            n1418;
wire            n14180;
wire            n14181;
wire            n14182;
wire            n14183;
wire            n14184;
wire            n14185;
wire            n14186;
wire            n14187;
wire            n14188;
wire            n14189;
wire            n1419;
wire            n14190;
wire            n14191;
wire            n14192;
wire            n14193;
wire            n14194;
wire            n14195;
wire            n14196;
wire            n14197;
wire            n14198;
wire            n14199;
wire            n142;
wire            n1420;
wire            n14200;
wire            n14201;
wire            n14202;
wire            n14203;
wire            n14204;
wire            n14205;
wire            n14206;
wire            n14207;
wire            n14208;
wire            n14209;
wire            n1421;
wire            n14210;
wire            n14211;
wire            n14212;
wire            n14213;
wire            n14214;
wire            n14215;
wire            n14216;
wire            n14217;
wire            n14218;
wire            n14219;
wire            n1422;
wire            n14220;
wire            n14221;
wire            n14222;
wire            n14223;
wire            n14224;
wire            n14225;
wire            n14226;
wire            n14227;
wire            n14228;
wire            n14229;
wire            n1423;
wire            n14230;
wire            n14231;
wire            n14232;
wire            n14233;
wire            n14234;
wire            n14235;
wire            n14236;
wire            n14237;
wire            n14238;
wire            n14239;
wire            n1424;
wire            n14240;
wire            n14241;
wire            n14242;
wire            n14243;
wire            n14244;
wire            n14245;
wire            n14246;
wire            n14247;
wire            n14248;
wire            n14249;
wire            n1425;
wire            n14250;
wire            n14251;
wire            n14252;
wire            n14253;
wire            n14254;
wire            n14255;
wire            n14256;
wire            n14257;
wire            n14258;
wire            n14259;
wire            n1426;
wire            n14260;
wire            n14261;
wire            n14262;
wire            n14263;
wire            n14264;
wire            n14265;
wire            n14266;
wire            n14267;
wire            n14268;
wire            n14269;
wire            n1427;
wire            n14270;
wire            n14271;
wire            n14272;
wire            n14273;
wire            n14274;
wire            n14275;
wire            n14276;
wire            n14277;
wire            n14278;
wire            n14279;
wire            n1428;
wire            n14280;
wire            n14281;
wire            n14282;
wire            n14283;
wire            n14284;
wire            n14285;
wire            n14286;
wire            n14287;
wire            n14288;
wire            n14289;
wire            n1429;
wire            n14290;
wire            n14291;
wire            n14292;
wire            n14293;
wire            n14294;
wire            n14295;
wire            n14296;
wire            n14297;
wire            n14298;
wire            n14299;
wire            n143;
wire            n1430;
wire            n14300;
wire            n14301;
wire            n14302;
wire            n14303;
wire            n14304;
wire            n14305;
wire            n14306;
wire            n14307;
wire            n14308;
wire            n14309;
wire            n1431;
wire            n14310;
wire            n14311;
wire            n14312;
wire            n14313;
wire            n14314;
wire            n14315;
wire            n14316;
wire            n14317;
wire            n14318;
wire            n14319;
wire            n1432;
wire            n14320;
wire            n14321;
wire            n14322;
wire            n14323;
wire            n14324;
wire            n14325;
wire            n14326;
wire            n14327;
wire            n14328;
wire            n14329;
wire            n1433;
wire            n14330;
wire            n14331;
wire            n14332;
wire            n14333;
wire            n14334;
wire            n14335;
wire            n14336;
wire            n14337;
wire            n14338;
wire            n14339;
wire            n1434;
wire            n14340;
wire            n14341;
wire            n14342;
wire            n14343;
wire            n14344;
wire            n14345;
wire            n14346;
wire            n14347;
wire            n14348;
wire            n14349;
wire            n1435;
wire            n14350;
wire            n14351;
wire            n14352;
wire            n14353;
wire            n14354;
wire            n14355;
wire            n14356;
wire            n14357;
wire            n14358;
wire            n14359;
wire            n1436;
wire            n14360;
wire            n14361;
wire            n14362;
wire            n14363;
wire            n14364;
wire            n14365;
wire            n14366;
wire            n14367;
wire            n14368;
wire            n14369;
wire            n1437;
wire            n14370;
wire            n14371;
wire            n14372;
wire            n14373;
wire            n14374;
wire            n14375;
wire            n14376;
wire            n14377;
wire            n14378;
wire            n14379;
wire            n1438;
wire            n14380;
wire            n14381;
wire            n14382;
wire            n14383;
wire            n14384;
wire            n14385;
wire            n14386;
wire            n14387;
wire            n14388;
wire            n14389;
wire            n1439;
wire            n14390;
wire            n14391;
wire            n14392;
wire            n14393;
wire            n14394;
wire            n14395;
wire            n14396;
wire            n14397;
wire            n14398;
wire            n14399;
wire            n144;
wire            n1440;
wire            n14400;
wire            n14401;
wire            n14402;
wire            n14403;
wire            n14404;
wire            n14405;
wire            n14406;
wire            n14407;
wire            n14408;
wire            n14409;
wire            n1441;
wire            n14410;
wire            n14411;
wire            n14412;
wire            n14413;
wire            n14414;
wire            n14415;
wire            n14416;
wire            n14417;
wire            n14418;
wire            n14419;
wire            n1442;
wire            n14420;
wire            n14421;
wire            n14422;
wire            n14423;
wire            n14424;
wire            n14425;
wire            n14426;
wire            n14427;
wire            n14428;
wire            n14429;
wire            n1443;
wire            n14430;
wire            n14431;
wire            n14432;
wire            n14433;
wire            n14434;
wire            n14435;
wire            n14436;
wire            n14437;
wire            n14438;
wire            n14439;
wire            n1444;
wire            n14440;
wire            n14441;
wire            n14442;
wire            n14443;
wire            n14444;
wire            n14445;
wire            n14446;
wire            n14447;
wire            n14448;
wire            n14449;
wire            n1445;
wire            n14450;
wire            n14451;
wire            n14452;
wire            n14453;
wire            n14454;
wire            n14455;
wire            n14456;
wire            n14457;
wire            n14458;
wire            n14459;
wire            n1446;
wire            n14460;
wire            n14461;
wire            n14462;
wire            n14463;
wire            n14464;
wire            n14465;
wire            n14466;
wire            n14467;
wire            n14468;
wire            n14469;
wire            n1447;
wire            n14470;
wire            n14471;
wire            n14472;
wire            n14473;
wire            n14474;
wire            n14475;
wire            n14476;
wire            n14477;
wire            n14478;
wire            n14479;
wire            n1448;
wire            n14480;
wire            n14481;
wire            n14482;
wire            n14483;
wire            n14484;
wire            n14485;
wire            n14486;
wire            n14487;
wire            n14488;
wire            n14489;
wire            n1449;
wire            n14490;
wire            n14491;
wire            n14492;
wire            n14493;
wire            n14494;
wire            n14495;
wire            n14496;
wire            n14497;
wire            n14498;
wire            n14499;
wire            n145;
wire            n1450;
wire            n14500;
wire            n14501;
wire            n14502;
wire            n14503;
wire            n14504;
wire            n14505;
wire            n14506;
wire            n14507;
wire            n14508;
wire            n14509;
wire            n1451;
wire            n14510;
wire            n14511;
wire            n14512;
wire            n14513;
wire            n14514;
wire            n14515;
wire            n14516;
wire            n14517;
wire            n14518;
wire            n14519;
wire            n1452;
wire            n14520;
wire            n14521;
wire            n14522;
wire            n14523;
wire            n14524;
wire            n14525;
wire            n14526;
wire            n14527;
wire            n14528;
wire            n14529;
wire            n1453;
wire            n14530;
wire            n14531;
wire            n14532;
wire            n14533;
wire            n14534;
wire            n14535;
wire            n14536;
wire            n14537;
wire            n14538;
wire            n14539;
wire            n1454;
wire            n14540;
wire            n14541;
wire            n14542;
wire            n14543;
wire            n14544;
wire            n14545;
wire            n14546;
wire            n14547;
wire            n14548;
wire            n14549;
wire            n1455;
wire            n14550;
wire            n14551;
wire            n14552;
wire            n14553;
wire            n14554;
wire            n14555;
wire            n14556;
wire            n14557;
wire            n14558;
wire            n14559;
wire            n1456;
wire            n14560;
wire            n14561;
wire            n14562;
wire            n14563;
wire            n14564;
wire            n14565;
wire            n14566;
wire            n14567;
wire            n14568;
wire            n14569;
wire            n1457;
wire            n14570;
wire            n14571;
wire            n14572;
wire            n14573;
wire            n14574;
wire            n14575;
wire            n14576;
wire            n14577;
wire            n14578;
wire            n14579;
wire            n1458;
wire            n14580;
wire            n14581;
wire            n14582;
wire            n14583;
wire            n14584;
wire            n14585;
wire            n14586;
wire            n14587;
wire            n14588;
wire            n14589;
wire            n1459;
wire            n14590;
wire            n14591;
wire            n14592;
wire            n14593;
wire            n14594;
wire            n14595;
wire            n14596;
wire            n14597;
wire            n14598;
wire            n14599;
wire            n146;
wire            n1460;
wire            n14600;
wire            n14601;
wire            n14602;
wire            n14603;
wire            n14604;
wire            n14605;
wire            n14606;
wire            n14607;
wire            n14608;
wire            n14609;
wire            n1461;
wire            n14610;
wire            n14611;
wire            n14612;
wire            n14613;
wire            n14614;
wire            n14615;
wire            n14616;
wire            n14617;
wire            n14618;
wire            n14619;
wire            n1462;
wire            n14620;
wire            n14621;
wire            n14622;
wire            n14623;
wire            n14624;
wire            n14625;
wire            n14626;
wire            n14627;
wire            n14628;
wire            n14629;
wire            n1463;
wire            n14630;
wire            n14631;
wire            n14632;
wire            n14633;
wire            n14634;
wire            n14635;
wire            n14636;
wire            n14637;
wire            n14638;
wire            n14639;
wire            n1464;
wire            n14640;
wire            n14641;
wire            n14642;
wire            n14643;
wire            n14644;
wire            n14645;
wire            n14646;
wire            n14647;
wire            n14648;
wire            n14649;
wire            n1465;
wire            n14650;
wire            n14651;
wire            n14652;
wire            n14653;
wire            n14654;
wire            n14655;
wire            n14656;
wire            n14657;
wire            n14658;
wire            n14659;
wire            n1466;
wire            n14660;
wire            n14661;
wire            n14662;
wire            n14663;
wire            n14664;
wire            n14665;
wire            n14666;
wire            n14667;
wire            n14668;
wire            n14669;
wire            n1467;
wire            n14670;
wire            n14671;
wire            n14672;
wire            n14673;
wire            n14674;
wire            n14675;
wire            n14676;
wire            n14677;
wire            n14678;
wire            n14679;
wire            n1468;
wire            n14680;
wire            n14681;
wire            n14682;
wire            n14683;
wire            n14684;
wire            n14685;
wire            n14686;
wire            n14687;
wire            n14688;
wire            n14689;
wire            n1469;
wire            n14690;
wire            n14691;
wire            n14692;
wire            n14693;
wire            n14694;
wire            n14695;
wire            n14696;
wire            n14697;
wire            n14698;
wire            n14699;
wire            n147;
wire            n1470;
wire            n14700;
wire            n14701;
wire            n14702;
wire            n14703;
wire            n14704;
wire            n14705;
wire            n14706;
wire            n14707;
wire            n14708;
wire            n14709;
wire            n1471;
wire            n14710;
wire            n14711;
wire            n14712;
wire            n14713;
wire            n14714;
wire            n14715;
wire            n14716;
wire            n14717;
wire            n14718;
wire            n14719;
wire            n1472;
wire            n14720;
wire            n14721;
wire            n14722;
wire            n14723;
wire            n14724;
wire            n14725;
wire            n14726;
wire            n14727;
wire            n14728;
wire            n14729;
wire            n1473;
wire            n14730;
wire            n14731;
wire            n14732;
wire            n14733;
wire            n14734;
wire            n14735;
wire            n14736;
wire            n14737;
wire            n14738;
wire            n14739;
wire            n1474;
wire            n14740;
wire            n14741;
wire            n14742;
wire            n14743;
wire            n14744;
wire            n14745;
wire            n14746;
wire            n14747;
wire            n14748;
wire            n14749;
wire            n1475;
wire            n14750;
wire            n14751;
wire            n14752;
wire            n14753;
wire            n14754;
wire            n14755;
wire            n14756;
wire            n14757;
wire            n14758;
wire            n14759;
wire            n1476;
wire            n14760;
wire            n14761;
wire            n14762;
wire            n14763;
wire            n14764;
wire            n14765;
wire            n14766;
wire            n14767;
wire            n14768;
wire            n14769;
wire            n1477;
wire            n14770;
wire            n14771;
wire            n14772;
wire            n14773;
wire            n14774;
wire            n14775;
wire            n14776;
wire            n14777;
wire            n14778;
wire            n14779;
wire            n1478;
wire            n14780;
wire            n14781;
wire            n14782;
wire            n14783;
wire            n14784;
wire            n14785;
wire            n14786;
wire            n14787;
wire            n14788;
wire            n14789;
wire            n1479;
wire            n14790;
wire            n14791;
wire            n14792;
wire            n14793;
wire            n14794;
wire            n14795;
wire            n14796;
wire            n14797;
wire            n14798;
wire            n14799;
wire            n148;
wire            n1480;
wire            n14800;
wire            n14801;
wire            n14802;
wire            n14803;
wire            n14804;
wire            n14805;
wire            n14806;
wire            n14807;
wire            n14808;
wire            n14809;
wire            n1481;
wire            n14810;
wire            n14811;
wire            n14812;
wire            n14813;
wire            n14814;
wire            n14815;
wire            n14816;
wire            n14817;
wire            n14818;
wire            n14819;
wire            n1482;
wire            n14820;
wire            n14821;
wire            n14822;
wire            n14823;
wire            n14824;
wire            n14825;
wire            n14826;
wire            n14827;
wire            n14828;
wire            n14829;
wire            n1483;
wire            n14830;
wire            n14831;
wire            n14832;
wire            n14833;
wire            n14834;
wire            n14835;
wire            n14836;
wire            n14837;
wire            n14838;
wire            n14839;
wire            n1484;
wire            n14840;
wire            n14841;
wire            n14842;
wire            n14843;
wire            n14844;
wire            n14845;
wire            n14846;
wire            n14847;
wire            n14848;
wire            n14849;
wire            n1485;
wire            n14850;
wire            n14851;
wire            n14852;
wire            n14853;
wire            n14854;
wire            n14855;
wire            n14856;
wire            n14857;
wire            n14858;
wire            n14859;
wire            n1486;
wire            n14860;
wire            n14861;
wire            n14862;
wire            n14863;
wire            n14864;
wire            n14865;
wire            n14866;
wire            n14867;
wire            n14868;
wire            n14869;
wire            n1487;
wire            n14870;
wire            n14871;
wire            n14872;
wire            n14873;
wire            n14874;
wire            n14875;
wire            n14876;
wire            n14877;
wire            n14878;
wire            n14879;
wire            n1488;
wire            n14880;
wire            n14881;
wire            n14882;
wire            n14883;
wire            n14884;
wire            n14885;
wire            n14886;
wire            n14887;
wire            n14888;
wire            n14889;
wire            n1489;
wire            n14890;
wire            n14891;
wire            n14892;
wire            n14893;
wire            n14894;
wire            n14895;
wire            n14896;
wire            n14897;
wire            n14898;
wire            n14899;
wire            n149;
wire            n1490;
wire            n14900;
wire            n14901;
wire            n14902;
wire            n14903;
wire            n14904;
wire            n14905;
wire            n14906;
wire            n14907;
wire            n14908;
wire            n14909;
wire            n1491;
wire            n14910;
wire            n14911;
wire            n14912;
wire            n14913;
wire            n14914;
wire            n14915;
wire            n14916;
wire            n14917;
wire            n14918;
wire            n14919;
wire            n1492;
wire            n14920;
wire            n14921;
wire            n14922;
wire            n14923;
wire            n14924;
wire            n14925;
wire            n14926;
wire            n14927;
wire            n14928;
wire            n14929;
wire            n1493;
wire            n14930;
wire            n14931;
wire            n14932;
wire            n14933;
wire            n14934;
wire            n14935;
wire            n14936;
wire            n14937;
wire            n14938;
wire            n14939;
wire            n1494;
wire            n14940;
wire            n14941;
wire            n14942;
wire            n14943;
wire            n14944;
wire            n14945;
wire            n14946;
wire            n14947;
wire            n14948;
wire            n14949;
wire            n1495;
wire            n14950;
wire            n14951;
wire            n14952;
wire            n14953;
wire            n14954;
wire            n14955;
wire            n14956;
wire            n14957;
wire            n14958;
wire            n14959;
wire            n1496;
wire            n14960;
wire            n14961;
wire            n14962;
wire            n14963;
wire            n14964;
wire            n14965;
wire            n14966;
wire            n14967;
wire            n14968;
wire            n14969;
wire            n1497;
wire            n14970;
wire            n14971;
wire            n14972;
wire            n14973;
wire            n14974;
wire            n14975;
wire            n14976;
wire            n14977;
wire            n14978;
wire            n14979;
wire            n1498;
wire            n14980;
wire            n14981;
wire            n14982;
wire            n14983;
wire            n14984;
wire            n14985;
wire            n14986;
wire            n14987;
wire            n14988;
wire            n14989;
wire            n1499;
wire            n14990;
wire            n14991;
wire            n14992;
wire            n14993;
wire            n14994;
wire            n14995;
wire            n14996;
wire            n14997;
wire            n14998;
wire            n14999;
wire            n15;
wire            n150;
wire            n1500;
wire            n15000;
wire            n15001;
wire            n15002;
wire            n15003;
wire            n15004;
wire            n15005;
wire            n15006;
wire            n15007;
wire            n15008;
wire            n15009;
wire            n1501;
wire            n15010;
wire            n15011;
wire            n15012;
wire            n15013;
wire            n15014;
wire            n15015;
wire            n15016;
wire            n15017;
wire            n15018;
wire            n15019;
wire            n1502;
wire            n15020;
wire            n15021;
wire            n15022;
wire            n15023;
wire            n15024;
wire            n15025;
wire            n15026;
wire            n15027;
wire            n15028;
wire            n15029;
wire            n1503;
wire            n15030;
wire            n15031;
wire            n15032;
wire            n15033;
wire            n15034;
wire            n15035;
wire            n15036;
wire            n15037;
wire            n15038;
wire            n15039;
wire            n1504;
wire            n15040;
wire            n15041;
wire            n15042;
wire            n15043;
wire            n15044;
wire            n15045;
wire            n15046;
wire            n15047;
wire            n15048;
wire            n15049;
wire            n1505;
wire            n15050;
wire            n15051;
wire            n15052;
wire            n15053;
wire            n15054;
wire            n15055;
wire            n15056;
wire            n15057;
wire            n15058;
wire            n15059;
wire            n1506;
wire            n15060;
wire            n15061;
wire            n15062;
wire            n15063;
wire            n15064;
wire            n15065;
wire            n15066;
wire            n15067;
wire            n15068;
wire            n15069;
wire            n1507;
wire            n15070;
wire            n15071;
wire            n15072;
wire            n15073;
wire            n15074;
wire            n15075;
wire            n15076;
wire            n15077;
wire            n15078;
wire            n15079;
wire            n1508;
wire            n15080;
wire            n15081;
wire            n15082;
wire            n15083;
wire            n15084;
wire            n15085;
wire            n15086;
wire            n15087;
wire            n15088;
wire            n15089;
wire            n1509;
wire            n15090;
wire            n15091;
wire            n15092;
wire            n15093;
wire            n15094;
wire            n15095;
wire            n15096;
wire            n15097;
wire            n15098;
wire            n15099;
wire            n151;
wire            n1510;
wire            n15100;
wire            n15101;
wire            n15102;
wire            n15103;
wire            n15104;
wire            n15105;
wire            n15106;
wire            n15107;
wire            n15108;
wire            n15109;
wire            n1511;
wire            n15110;
wire            n15111;
wire            n15112;
wire            n15113;
wire            n15114;
wire            n15115;
wire            n15116;
wire            n15117;
wire            n15118;
wire            n15119;
wire            n1512;
wire            n15120;
wire            n15121;
wire            n15122;
wire            n15123;
wire            n15124;
wire            n15125;
wire            n15126;
wire            n15127;
wire            n15128;
wire            n15129;
wire            n1513;
wire            n15130;
wire            n15131;
wire            n15132;
wire            n15133;
wire            n15134;
wire            n15135;
wire            n15136;
wire            n15137;
wire            n15138;
wire            n15139;
wire            n1514;
wire            n15140;
wire            n15141;
wire            n15142;
wire            n15143;
wire            n15144;
wire            n15145;
wire            n15146;
wire            n15147;
wire            n15148;
wire            n15149;
wire            n1515;
wire            n15150;
wire            n15151;
wire            n15152;
wire            n15153;
wire            n15154;
wire            n15155;
wire            n15156;
wire            n15157;
wire            n15158;
wire            n15159;
wire            n1516;
wire            n15160;
wire            n15161;
wire            n15162;
wire            n15163;
wire            n15164;
wire            n15165;
wire            n15166;
wire            n15167;
wire            n15168;
wire            n15169;
wire            n1517;
wire            n15170;
wire            n15171;
wire            n15172;
wire            n15173;
wire            n15174;
wire            n15175;
wire            n15176;
wire            n15177;
wire            n15178;
wire            n15179;
wire            n1518;
wire            n15180;
wire            n15181;
wire            n15182;
wire            n15183;
wire            n15184;
wire            n15185;
wire            n15186;
wire            n15187;
wire            n15188;
wire            n15189;
wire            n1519;
wire            n15190;
wire            n15191;
wire            n15192;
wire            n15193;
wire            n15194;
wire            n15195;
wire            n15196;
wire            n15197;
wire            n15198;
wire            n15199;
wire            n152;
wire            n1520;
wire            n15200;
wire            n15201;
wire            n15202;
wire            n15203;
wire            n15204;
wire            n15205;
wire            n15206;
wire            n15207;
wire            n15208;
wire            n15209;
wire            n1521;
wire            n15210;
wire            n15211;
wire            n15212;
wire            n15213;
wire            n15214;
wire            n15215;
wire            n15216;
wire            n15217;
wire            n15218;
wire            n15219;
wire            n1522;
wire            n15220;
wire            n15221;
wire            n15222;
wire            n15223;
wire            n15224;
wire            n15225;
wire            n15226;
wire            n15227;
wire            n15228;
wire            n15229;
wire            n1523;
wire            n15230;
wire            n15231;
wire            n15232;
wire            n15233;
wire            n15234;
wire            n15235;
wire            n15236;
wire            n15237;
wire            n15238;
wire            n15239;
wire            n1524;
wire            n15240;
wire            n15241;
wire            n15242;
wire            n15243;
wire            n15244;
wire            n15245;
wire            n15246;
wire            n15247;
wire            n15248;
wire            n15249;
wire            n1525;
wire            n15250;
wire            n15251;
wire            n15252;
wire            n15253;
wire            n15254;
wire            n15255;
wire            n15256;
wire            n15257;
wire            n15258;
wire            n15259;
wire            n1526;
wire            n15260;
wire            n15261;
wire            n15262;
wire            n15263;
wire            n15264;
wire            n15265;
wire            n15266;
wire            n15267;
wire            n15268;
wire            n15269;
wire            n1527;
wire            n15270;
wire            n15271;
wire            n15272;
wire            n15273;
wire            n15274;
wire            n15275;
wire            n15276;
wire            n15277;
wire            n15278;
wire            n15279;
wire            n1528;
wire            n15280;
wire            n15281;
wire            n15282;
wire            n15283;
wire            n15284;
wire            n15285;
wire            n15286;
wire            n15287;
wire            n15288;
wire            n15289;
wire            n1529;
wire            n15290;
wire            n15291;
wire            n15292;
wire            n15293;
wire            n15294;
wire            n15295;
wire            n15296;
wire            n15297;
wire            n15298;
wire            n15299;
wire            n153;
wire            n1530;
wire            n15300;
wire            n15301;
wire            n15302;
wire            n15303;
wire            n15304;
wire            n15305;
wire            n15306;
wire            n15307;
wire            n15308;
wire            n15309;
wire            n1531;
wire            n15310;
wire            n15311;
wire            n15312;
wire            n15313;
wire            n15314;
wire            n15315;
wire            n15316;
wire            n15317;
wire            n15318;
wire            n15319;
wire            n1532;
wire            n15320;
wire            n15321;
wire            n15322;
wire            n15323;
wire            n15324;
wire            n15325;
wire            n15326;
wire            n15327;
wire            n15328;
wire            n15329;
wire            n1533;
wire            n15330;
wire            n15331;
wire            n15332;
wire            n15333;
wire            n15334;
wire            n15335;
wire            n15336;
wire            n15337;
wire            n15338;
wire            n15339;
wire            n1534;
wire            n15340;
wire            n15341;
wire            n15342;
wire            n15343;
wire            n15344;
wire            n15345;
wire            n15346;
wire            n15347;
wire            n15348;
wire            n15349;
wire            n1535;
wire            n15350;
wire            n15351;
wire            n15352;
wire            n15353;
wire            n15354;
wire            n15355;
wire            n15356;
wire            n15357;
wire            n15358;
wire            n15359;
wire            n1536;
wire            n15360;
wire            n15361;
wire            n15362;
wire            n15363;
wire            n15364;
wire            n15365;
wire            n15366;
wire            n15367;
wire            n15368;
wire            n15369;
wire            n1537;
wire            n15370;
wire            n15371;
wire            n15372;
wire            n15373;
wire            n15374;
wire            n15375;
wire            n15376;
wire            n15377;
wire            n15378;
wire            n15379;
wire            n1538;
wire            n15380;
wire            n15381;
wire            n15382;
wire            n15383;
wire            n15384;
wire            n15385;
wire            n15386;
wire            n15387;
wire            n15388;
wire            n15389;
wire            n1539;
wire            n15390;
wire            n15391;
wire            n15392;
wire            n15393;
wire            n15394;
wire            n15395;
wire            n15396;
wire            n15397;
wire            n15398;
wire            n15399;
wire            n154;
wire            n1540;
wire            n15400;
wire            n15401;
wire            n15402;
wire            n15403;
wire            n15404;
wire            n15405;
wire            n15406;
wire            n15407;
wire            n15408;
wire            n15409;
wire            n1541;
wire            n15410;
wire            n15411;
wire            n15412;
wire            n15413;
wire            n15414;
wire            n15415;
wire            n15416;
wire            n15417;
wire            n15418;
wire            n15419;
wire            n1542;
wire            n15420;
wire            n15421;
wire            n15422;
wire            n15423;
wire            n15424;
wire            n15425;
wire            n15426;
wire            n15427;
wire            n15428;
wire            n15429;
wire            n1543;
wire            n15430;
wire            n15431;
wire            n15432;
wire            n15433;
wire            n15434;
wire            n15435;
wire            n15436;
wire            n15437;
wire            n15438;
wire            n15439;
wire            n1544;
wire            n15440;
wire            n15441;
wire            n15442;
wire            n15443;
wire            n15444;
wire            n15445;
wire            n15446;
wire            n15447;
wire            n15448;
wire            n15449;
wire            n1545;
wire            n15450;
wire            n15451;
wire            n15452;
wire            n15453;
wire            n15454;
wire            n15455;
wire            n15456;
wire            n15457;
wire            n15458;
wire            n15459;
wire            n1546;
wire            n15460;
wire            n15461;
wire            n15462;
wire            n15463;
wire            n15464;
wire            n15465;
wire            n15466;
wire            n15467;
wire            n15468;
wire            n15469;
wire            n1547;
wire            n15470;
wire            n15471;
wire            n15472;
wire            n15473;
wire            n15474;
wire            n15475;
wire            n15476;
wire            n15477;
wire            n15478;
wire            n15479;
wire            n1548;
wire            n15480;
wire            n15481;
wire            n15482;
wire            n15483;
wire            n15484;
wire            n15485;
wire            n15486;
wire            n15487;
wire            n15488;
wire            n15489;
wire            n1549;
wire            n15490;
wire            n15491;
wire            n15492;
wire            n15493;
wire            n15494;
wire            n15495;
wire            n15496;
wire            n15497;
wire            n15498;
wire            n15499;
wire            n155;
wire            n1550;
wire            n15500;
wire            n15501;
wire            n15502;
wire            n15503;
wire            n15504;
wire            n15505;
wire            n15506;
wire            n15507;
wire            n15508;
wire            n15509;
wire            n1551;
wire            n15510;
wire            n15511;
wire            n15512;
wire            n15513;
wire            n15514;
wire            n15515;
wire            n15516;
wire            n15517;
wire            n15518;
wire            n15519;
wire            n1552;
wire            n15520;
wire            n15521;
wire            n15522;
wire            n15523;
wire            n15524;
wire            n15525;
wire            n15526;
wire            n15527;
wire            n15528;
wire            n15529;
wire            n1553;
wire            n15530;
wire            n15531;
wire            n15532;
wire            n15533;
wire            n15534;
wire            n15535;
wire            n15536;
wire            n15537;
wire            n15538;
wire            n15539;
wire            n1554;
wire            n15540;
wire            n15541;
wire            n15542;
wire            n15543;
wire            n15544;
wire            n15545;
wire            n15546;
wire            n15547;
wire            n15548;
wire            n15549;
wire            n1555;
wire            n15550;
wire            n15551;
wire            n15552;
wire            n15553;
wire            n15554;
wire            n15555;
wire            n15556;
wire            n15557;
wire            n15558;
wire            n15559;
wire            n1556;
wire            n15560;
wire            n15561;
wire            n15562;
wire            n15563;
wire            n15564;
wire            n15565;
wire            n15566;
wire            n15567;
wire            n15568;
wire            n15569;
wire            n1557;
wire            n15570;
wire            n15571;
wire            n15572;
wire            n15573;
wire            n15574;
wire            n15575;
wire            n15576;
wire            n15577;
wire      [1:0] n15578;
wire            n15579;
wire            n1558;
wire            n15580;
wire            n15581;
wire            n15582;
wire            n15583;
wire            n15584;
wire            n15585;
wire            n15586;
wire            n15587;
wire            n15588;
wire            n15589;
wire            n1559;
wire      [2:0] n15590;
wire            n15591;
wire            n15592;
wire            n15593;
wire            n15594;
wire            n15595;
wire            n15596;
wire            n15597;
wire            n15598;
wire            n15599;
wire            n156;
wire            n1560;
wire            n15600;
wire            n15601;
wire            n15602;
wire            n15603;
wire            n15604;
wire            n15605;
wire            n15606;
wire            n15607;
wire            n15608;
wire            n15609;
wire            n1561;
wire            n15610;
wire            n15611;
wire            n15612;
wire            n15613;
wire            n15614;
wire            n15615;
wire            n15616;
wire            n15617;
wire            n15618;
wire            n15619;
wire            n1562;
wire            n15620;
wire            n15621;
wire            n15622;
wire            n15623;
wire            n15624;
wire            n15625;
wire            n15626;
wire            n15627;
wire            n15628;
wire            n15629;
wire            n1563;
wire            n15630;
wire            n15631;
wire            n15632;
wire            n15633;
wire            n15634;
wire            n15635;
wire            n15636;
wire            n15637;
wire            n15638;
wire            n15639;
wire            n1564;
wire            n15640;
wire            n15641;
wire            n15642;
wire            n15643;
wire            n15644;
wire            n15645;
wire            n15646;
wire            n15647;
wire            n15648;
wire            n15649;
wire            n1565;
wire            n15650;
wire            n15651;
wire            n15652;
wire            n15653;
wire            n15654;
wire            n15655;
wire            n15656;
wire            n15657;
wire            n15658;
wire            n15659;
wire            n1566;
wire            n15660;
wire            n15661;
wire            n15662;
wire            n15663;
wire            n15664;
wire            n15665;
wire            n15666;
wire            n15667;
wire            n15668;
wire            n15669;
wire            n1567;
wire            n15670;
wire            n15671;
wire            n15672;
wire            n15673;
wire            n15674;
wire            n15675;
wire            n15676;
wire            n15677;
wire            n15678;
wire            n15679;
wire            n1568;
wire            n15680;
wire            n15681;
wire            n15682;
wire            n15683;
wire            n15684;
wire            n15685;
wire            n15686;
wire            n15687;
wire            n15688;
wire            n15689;
wire            n1569;
wire            n15690;
wire            n15691;
wire            n15692;
wire            n15693;
wire            n15694;
wire            n15695;
wire            n15696;
wire            n15697;
wire            n15698;
wire            n15699;
wire            n157;
wire            n1570;
wire            n15700;
wire            n15701;
wire            n15702;
wire            n15703;
wire            n15704;
wire            n15705;
wire            n15706;
wire            n15707;
wire            n15708;
wire            n15709;
wire            n1571;
wire            n15710;
wire            n15711;
wire            n15712;
wire            n15713;
wire            n15714;
wire            n15715;
wire            n15716;
wire            n15717;
wire            n15718;
wire            n15719;
wire            n1572;
wire            n15720;
wire            n15721;
wire            n15722;
wire            n15723;
wire            n15724;
wire            n15725;
wire            n15726;
wire            n15727;
wire            n15728;
wire            n15729;
wire            n1573;
wire            n15730;
wire            n15731;
wire            n15732;
wire            n15733;
wire            n15734;
wire            n15735;
wire            n15736;
wire            n15737;
wire            n15738;
wire            n15739;
wire            n1574;
wire            n15740;
wire            n15741;
wire            n15742;
wire            n15743;
wire            n15744;
wire            n15745;
wire            n15746;
wire            n15747;
wire            n15748;
wire            n15749;
wire            n1575;
wire            n15750;
wire            n15751;
wire            n15752;
wire            n15753;
wire            n15754;
wire            n15755;
wire            n15756;
wire            n15757;
wire            n15758;
wire            n15759;
wire            n1576;
wire            n15760;
wire            n15761;
wire            n15762;
wire            n15763;
wire            n15764;
wire            n15765;
wire            n15766;
wire            n15767;
wire            n15768;
wire            n15769;
wire            n1577;
wire            n15770;
wire            n15771;
wire            n15772;
wire            n15773;
wire            n15774;
wire            n15775;
wire            n15776;
wire            n15777;
wire            n15778;
wire            n15779;
wire            n1578;
wire            n15780;
wire            n15781;
wire            n15782;
wire            n15783;
wire            n15784;
wire            n15785;
wire            n15786;
wire            n15787;
wire            n15788;
wire            n15789;
wire            n1579;
wire            n15790;
wire            n15791;
wire            n15792;
wire            n15793;
wire            n15794;
wire            n15795;
wire            n15796;
wire            n15797;
wire            n15798;
wire            n15799;
wire            n158;
wire            n1580;
wire            n15800;
wire            n15801;
wire            n15802;
wire            n15803;
wire            n15804;
wire            n15805;
wire            n15806;
wire            n15807;
wire            n15808;
wire            n15809;
wire            n1581;
wire            n15810;
wire            n15811;
wire      [3:0] n15812;
wire            n15813;
wire            n15814;
wire            n15815;
wire            n15816;
wire            n15817;
wire            n15818;
wire            n15819;
wire            n1582;
wire            n15820;
wire            n15821;
wire            n15822;
wire            n15823;
wire            n15824;
wire            n15825;
wire            n15826;
wire            n15827;
wire            n15828;
wire            n15829;
wire            n1583;
wire      [4:0] n15830;
wire            n15831;
wire            n15832;
wire            n15833;
wire            n15834;
wire            n15835;
wire            n15836;
wire            n15837;
wire            n15838;
wire            n15839;
wire            n1584;
wire            n15840;
wire            n15841;
wire            n15842;
wire            n15843;
wire            n15844;
wire            n15845;
wire            n15846;
wire            n15847;
wire            n15848;
wire            n15849;
wire            n1585;
wire            n15850;
wire            n15851;
wire            n15852;
wire            n15853;
wire            n15854;
wire            n15855;
wire            n15856;
wire            n15857;
wire            n15858;
wire            n15859;
wire            n1586;
wire            n15860;
wire            n15861;
wire            n15862;
wire            n15863;
wire            n15864;
wire            n15865;
wire            n15866;
wire            n15867;
wire            n15868;
wire            n15869;
wire            n1587;
wire            n15870;
wire            n15871;
wire            n15872;
wire            n15873;
wire            n15874;
wire            n15875;
wire            n15876;
wire            n15877;
wire            n15878;
wire            n15879;
wire            n1588;
wire            n15880;
wire            n15881;
wire            n15882;
wire            n15883;
wire            n15884;
wire            n15885;
wire            n15886;
wire            n15887;
wire            n15888;
wire            n15889;
wire            n1589;
wire            n15890;
wire            n15891;
wire            n15892;
wire            n15893;
wire            n15894;
wire            n15895;
wire            n15896;
wire            n15897;
wire            n15898;
wire            n15899;
wire            n159;
wire            n1590;
wire            n15900;
wire            n15901;
wire            n15902;
wire            n15903;
wire            n15904;
wire            n15905;
wire            n15906;
wire            n15907;
wire            n15908;
wire            n15909;
wire            n1591;
wire            n15910;
wire            n15911;
wire            n15912;
wire            n15913;
wire            n15914;
wire            n15915;
wire            n15916;
wire            n15917;
wire            n15918;
wire            n15919;
wire            n1592;
wire            n15920;
wire            n15921;
wire            n15922;
wire            n15923;
wire            n15924;
wire            n15925;
wire            n15926;
wire            n15927;
wire            n15928;
wire            n15929;
wire            n1593;
wire            n15930;
wire            n15931;
wire            n15932;
wire            n15933;
wire            n15934;
wire            n15935;
wire            n15936;
wire            n15937;
wire            n15938;
wire            n15939;
wire            n1594;
wire            n15940;
wire            n15941;
wire            n15942;
wire            n15943;
wire            n15944;
wire            n15945;
wire            n15946;
wire            n15947;
wire            n15948;
wire            n15949;
wire            n1595;
wire            n15950;
wire            n15951;
wire            n15952;
wire            n15953;
wire            n15954;
wire            n15955;
wire            n15956;
wire            n15957;
wire            n15958;
wire            n15959;
wire            n1596;
wire            n15960;
wire            n15961;
wire            n15962;
wire            n15963;
wire            n15964;
wire            n15965;
wire            n15966;
wire            n15967;
wire            n15968;
wire            n15969;
wire            n1597;
wire            n15970;
wire            n15971;
wire            n15972;
wire            n15973;
wire            n15974;
wire            n15975;
wire            n15976;
wire            n15977;
wire            n15978;
wire            n15979;
wire            n1598;
wire            n15980;
wire            n15981;
wire            n15982;
wire            n15983;
wire            n15984;
wire            n15985;
wire            n15986;
wire            n15987;
wire            n15988;
wire            n15989;
wire            n1599;
wire            n15990;
wire            n15991;
wire            n15992;
wire            n15993;
wire            n15994;
wire            n15995;
wire            n15996;
wire            n15997;
wire            n15998;
wire            n15999;
wire            n16;
wire            n160;
wire            n1600;
wire            n16000;
wire            n16001;
wire            n16002;
wire            n16003;
wire            n16004;
wire            n16005;
wire            n16006;
wire            n16007;
wire            n16008;
wire            n16009;
wire            n1601;
wire            n16010;
wire            n16011;
wire            n16012;
wire            n16013;
wire            n16014;
wire            n16015;
wire            n16016;
wire            n16017;
wire            n16018;
wire            n16019;
wire            n1602;
wire            n16020;
wire            n16021;
wire            n16022;
wire            n16023;
wire            n16024;
wire            n16025;
wire            n16026;
wire            n16027;
wire            n16028;
wire            n16029;
wire            n1603;
wire            n16030;
wire            n16031;
wire            n16032;
wire            n16033;
wire            n16034;
wire            n16035;
wire            n16036;
wire            n16037;
wire            n16038;
wire            n16039;
wire            n1604;
wire            n16040;
wire            n16041;
wire            n16042;
wire            n16043;
wire            n16044;
wire            n16045;
wire            n16046;
wire            n16047;
wire            n16048;
wire            n16049;
wire            n1605;
wire            n16050;
wire            n16051;
wire            n16052;
wire      [5:0] n16053;
wire            n16054;
wire            n16055;
wire            n16056;
wire            n16057;
wire            n16058;
wire            n16059;
wire            n1606;
wire            n16060;
wire            n16061;
wire            n16062;
wire            n16063;
wire            n16064;
wire            n16065;
wire            n16066;
wire            n16067;
wire            n16068;
wire            n16069;
wire            n1607;
wire            n16070;
wire            n16071;
wire            n16072;
wire            n16073;
wire            n16074;
wire            n16075;
wire            n16076;
wire      [6:0] n16077;
wire            n16078;
wire            n16079;
wire            n1608;
wire            n16080;
wire            n16081;
wire            n16082;
wire            n16083;
wire            n16084;
wire            n16085;
wire            n16086;
wire            n16087;
wire            n16088;
wire            n16089;
wire            n1609;
wire            n16090;
wire            n16091;
wire            n16092;
wire            n16093;
wire            n16094;
wire            n16095;
wire            n16096;
wire            n16097;
wire            n16098;
wire            n16099;
wire            n161;
wire            n1610;
wire            n16100;
wire            n16101;
wire            n16102;
wire            n16103;
wire            n16104;
wire            n16105;
wire            n16106;
wire            n16107;
wire            n16108;
wire            n16109;
wire            n1611;
wire            n16110;
wire            n16111;
wire            n16112;
wire            n16113;
wire            n16114;
wire            n16115;
wire            n16116;
wire            n16117;
wire            n16118;
wire            n16119;
wire            n1612;
wire            n16120;
wire            n16121;
wire            n16122;
wire            n16123;
wire            n16124;
wire            n16125;
wire            n16126;
wire            n16127;
wire            n16128;
wire            n16129;
wire            n1613;
wire            n16130;
wire            n16131;
wire            n16132;
wire            n16133;
wire            n16134;
wire            n16135;
wire            n16136;
wire            n16137;
wire            n16138;
wire            n16139;
wire            n1614;
wire            n16140;
wire            n16141;
wire            n16142;
wire            n16143;
wire            n16144;
wire            n16145;
wire            n16146;
wire            n16147;
wire            n16148;
wire            n16149;
wire            n1615;
wire            n16150;
wire            n16151;
wire            n16152;
wire            n16153;
wire            n16154;
wire            n16155;
wire            n16156;
wire            n16157;
wire            n16158;
wire            n16159;
wire            n1616;
wire            n16160;
wire            n16161;
wire            n16162;
wire            n16163;
wire            n16164;
wire            n16165;
wire            n16166;
wire            n16167;
wire            n16168;
wire            n16169;
wire            n1617;
wire            n16170;
wire            n16171;
wire            n16172;
wire            n16173;
wire            n16174;
wire            n16175;
wire            n16176;
wire            n16177;
wire            n16178;
wire            n16179;
wire            n1618;
wire            n16180;
wire            n16181;
wire            n16182;
wire            n16183;
wire            n16184;
wire            n16185;
wire            n16186;
wire            n16187;
wire            n16188;
wire            n16189;
wire            n1619;
wire            n16190;
wire            n16191;
wire            n16192;
wire            n16193;
wire            n16194;
wire            n16195;
wire            n16196;
wire            n16197;
wire            n16198;
wire            n16199;
wire            n162;
wire            n1620;
wire            n16200;
wire            n16201;
wire            n16202;
wire            n16203;
wire      [7:0] n16204;
wire            n16205;
wire            n16206;
wire            n16207;
wire            n16208;
wire            n16209;
wire            n1621;
wire            n16210;
wire            n16211;
wire            n16212;
wire            n16213;
wire            n16214;
wire            n16215;
wire            n16216;
wire            n16217;
wire            n16218;
wire            n16219;
wire            n1622;
wire            n16220;
wire            n16221;
wire            n16222;
wire            n16223;
wire            n16224;
wire            n16225;
wire            n16226;
wire            n16227;
wire            n16228;
wire            n16229;
wire            n1623;
wire            n16230;
wire            n16231;
wire            n16232;
wire            n16233;
wire      [8:0] n16234;
wire            n16235;
wire            n16236;
wire            n16237;
wire            n16238;
wire            n16239;
wire            n1624;
wire            n16240;
wire            n16241;
wire            n16242;
wire            n16243;
wire            n16244;
wire            n16245;
wire            n16246;
wire            n16247;
wire            n16248;
wire            n16249;
wire            n1625;
wire            n16250;
wire            n16251;
wire            n16252;
wire            n16253;
wire            n16254;
wire            n16255;
wire            n16256;
wire            n16257;
wire            n16258;
wire            n16259;
wire            n1626;
wire            n16260;
wire            n16261;
wire            n16262;
wire            n16263;
wire            n16264;
wire            n16265;
wire            n16266;
wire            n16267;
wire            n16268;
wire            n16269;
wire            n1627;
wire            n16270;
wire            n16271;
wire            n16272;
wire            n16273;
wire            n16274;
wire            n16275;
wire            n16276;
wire            n16277;
wire            n16278;
wire            n16279;
wire            n1628;
wire            n16280;
wire            n16281;
wire            n16282;
wire            n16283;
wire            n16284;
wire            n16285;
wire            n16286;
wire            n16287;
wire            n16288;
wire            n16289;
wire            n1629;
wire            n16290;
wire            n16291;
wire            n16292;
wire            n16293;
wire            n16294;
wire            n16295;
wire            n16296;
wire            n16297;
wire            n16298;
wire            n16299;
wire            n163;
wire            n1630;
wire            n16300;
wire            n16301;
wire            n16302;
wire            n16303;
wire            n16304;
wire            n16305;
wire            n16306;
wire            n16307;
wire            n16308;
wire            n16309;
wire            n1631;
wire            n16310;
wire            n16311;
wire            n16312;
wire            n16313;
wire            n16314;
wire            n16315;
wire            n16316;
wire            n16317;
wire            n16318;
wire            n16319;
wire            n1632;
wire            n16320;
wire            n16321;
wire            n16322;
wire            n16323;
wire            n16324;
wire            n16325;
wire            n16326;
wire            n16327;
wire            n16328;
wire            n16329;
wire            n1633;
wire            n16330;
wire            n16331;
wire            n16332;
wire            n16333;
wire            n16334;
wire            n16335;
wire            n16336;
wire            n16337;
wire            n16338;
wire            n16339;
wire            n1634;
wire            n16340;
wire            n16341;
wire            n16342;
wire            n16343;
wire            n16344;
wire            n16345;
wire            n16346;
wire            n16347;
wire            n16348;
wire            n16349;
wire            n1635;
wire            n16350;
wire            n16351;
wire            n16352;
wire            n16353;
wire            n16354;
wire            n16355;
wire            n16356;
wire            n16357;
wire            n16358;
wire            n16359;
wire            n1636;
wire            n16360;
wire            n16361;
wire            n16362;
wire            n16363;
wire            n16364;
wire            n16365;
wire            n16366;
wire            n16367;
wire            n16368;
wire            n16369;
wire            n1637;
wire            n16370;
wire            n16371;
wire            n16372;
wire            n16373;
wire            n16374;
wire            n16375;
wire            n16376;
wire            n16377;
wire            n16378;
wire            n16379;
wire            n1638;
wire            n16380;
wire      [9:0] n16381;
wire            n16382;
wire            n16383;
wire            n16384;
wire            n16385;
wire            n16386;
wire            n16387;
wire            n16388;
wire            n16389;
wire            n1639;
wire            n16390;
wire            n16391;
wire            n16392;
wire            n16393;
wire            n16394;
wire            n16395;
wire            n16396;
wire            n16397;
wire            n16398;
wire            n16399;
wire            n164;
wire            n1640;
wire            n16400;
wire            n16401;
wire            n16402;
wire            n16403;
wire            n16404;
wire            n16405;
wire            n16406;
wire            n16407;
wire            n16408;
wire            n16409;
wire            n1641;
wire            n16410;
wire            n16411;
wire            n16412;
wire            n16413;
wire            n16414;
wire            n16415;
wire            n16416;
wire     [10:0] n16417;
wire            n16418;
wire            n16419;
wire            n1642;
wire            n16420;
wire            n16421;
wire            n16422;
wire            n16423;
wire            n16424;
wire            n16425;
wire            n16426;
wire            n16427;
wire            n16428;
wire            n16429;
wire            n1643;
wire            n16430;
wire            n16431;
wire            n16432;
wire            n16433;
wire            n16434;
wire            n16435;
wire            n16436;
wire            n16437;
wire            n16438;
wire            n16439;
wire            n1644;
wire            n16440;
wire            n16441;
wire            n16442;
wire            n16443;
wire            n16444;
wire            n16445;
wire            n16446;
wire            n16447;
wire            n16448;
wire            n16449;
wire            n1645;
wire            n16450;
wire            n16451;
wire            n16452;
wire            n16453;
wire            n16454;
wire            n16455;
wire            n16456;
wire            n16457;
wire            n16458;
wire            n16459;
wire            n1646;
wire            n16460;
wire            n16461;
wire            n16462;
wire            n16463;
wire            n16464;
wire            n16465;
wire            n16466;
wire            n16467;
wire            n16468;
wire            n16469;
wire            n1647;
wire            n16470;
wire            n16471;
wire            n16472;
wire            n16473;
wire            n16474;
wire            n16475;
wire            n16476;
wire            n16477;
wire            n16478;
wire            n16479;
wire            n1648;
wire            n16480;
wire            n16481;
wire            n16482;
wire            n16483;
wire            n16484;
wire            n16485;
wire            n16486;
wire            n16487;
wire            n16488;
wire            n16489;
wire            n1649;
wire            n16490;
wire            n16491;
wire            n16492;
wire            n16493;
wire            n16494;
wire            n16495;
wire            n16496;
wire            n16497;
wire            n16498;
wire            n16499;
wire            n165;
wire            n1650;
wire            n16500;
wire            n16501;
wire            n16502;
wire            n16503;
wire            n16504;
wire            n16505;
wire            n16506;
wire            n16507;
wire            n16508;
wire            n16509;
wire            n1651;
wire            n16510;
wire            n16511;
wire            n16512;
wire            n16513;
wire            n16514;
wire            n16515;
wire            n16516;
wire            n16517;
wire            n16518;
wire            n16519;
wire            n1652;
wire            n16520;
wire            n16521;
wire            n16522;
wire            n16523;
wire            n16524;
wire            n16525;
wire            n16526;
wire            n16527;
wire            n16528;
wire            n16529;
wire            n1653;
wire            n16530;
wire            n16531;
wire            n16532;
wire            n16533;
wire            n16534;
wire            n16535;
wire            n16536;
wire            n16537;
wire            n16538;
wire            n16539;
wire            n1654;
wire            n16540;
wire            n16541;
wire            n16542;
wire            n16543;
wire            n16544;
wire            n16545;
wire            n16546;
wire            n16547;
wire            n16548;
wire            n16549;
wire            n1655;
wire            n16550;
wire            n16551;
wire            n16552;
wire            n16553;
wire            n16554;
wire            n16555;
wire            n16556;
wire            n16557;
wire            n16558;
wire            n16559;
wire            n1656;
wire            n16560;
wire            n16561;
wire            n16562;
wire            n16563;
wire            n16564;
wire            n16565;
wire            n16566;
wire            n16567;
wire            n16568;
wire            n16569;
wire            n1657;
wire            n16570;
wire            n16571;
wire            n16572;
wire     [11:0] n16573;
wire            n16574;
wire            n16575;
wire            n16576;
wire            n16577;
wire            n16578;
wire            n16579;
wire            n1658;
wire            n16580;
wire            n16581;
wire            n16582;
wire            n16583;
wire            n16584;
wire            n16585;
wire            n16586;
wire            n16587;
wire            n16588;
wire            n16589;
wire            n1659;
wire            n16590;
wire            n16591;
wire            n16592;
wire            n16593;
wire            n16594;
wire            n16595;
wire            n16596;
wire            n16597;
wire            n16598;
wire            n16599;
wire            n166;
wire            n1660;
wire            n16600;
wire            n16601;
wire            n16602;
wire            n16603;
wire            n16604;
wire            n16605;
wire            n16606;
wire            n16607;
wire            n16608;
wire            n16609;
wire            n1661;
wire            n16610;
wire            n16611;
wire            n16612;
wire            n16613;
wire            n16614;
wire            n16615;
wire            n16616;
wire            n16617;
wire            n16618;
wire            n16619;
wire            n1662;
wire     [12:0] n16620;
wire            n16621;
wire            n16622;
wire            n16623;
wire            n16624;
wire            n16625;
wire            n16626;
wire            n16627;
wire            n16628;
wire            n16629;
wire            n1663;
wire            n16630;
wire            n16631;
wire            n16632;
wire            n16633;
wire            n16634;
wire            n16635;
wire            n16636;
wire            n16637;
wire            n16638;
wire            n16639;
wire            n1664;
wire            n16640;
wire            n16641;
wire            n16642;
wire            n16643;
wire            n16644;
wire            n16645;
wire            n16646;
wire            n16647;
wire            n16648;
wire            n16649;
wire            n1665;
wire            n16650;
wire            n16651;
wire            n16652;
wire            n16653;
wire            n16654;
wire            n16655;
wire            n16656;
wire            n16657;
wire            n16658;
wire            n16659;
wire            n1666;
wire            n16660;
wire            n16661;
wire            n16662;
wire            n16663;
wire            n16664;
wire            n16665;
wire            n16666;
wire            n16667;
wire            n16668;
wire            n16669;
wire            n1667;
wire            n16670;
wire            n16671;
wire            n16672;
wire            n16673;
wire            n16674;
wire            n16675;
wire            n16676;
wire            n16677;
wire            n16678;
wire            n16679;
wire            n1668;
wire            n16680;
wire            n16681;
wire            n16682;
wire            n16683;
wire            n16684;
wire            n16685;
wire            n16686;
wire            n16687;
wire            n16688;
wire            n16689;
wire            n1669;
wire            n16690;
wire            n16691;
wire            n16692;
wire            n16693;
wire            n16694;
wire            n16695;
wire            n16696;
wire            n16697;
wire            n16698;
wire            n16699;
wire            n167;
wire            n1670;
wire            n16700;
wire            n16701;
wire            n16702;
wire            n16703;
wire            n16704;
wire            n16705;
wire            n16706;
wire            n16707;
wire            n16708;
wire            n16709;
wire            n1671;
wire            n16710;
wire            n16711;
wire            n16712;
wire            n16713;
wire            n16714;
wire            n16715;
wire            n16716;
wire            n16717;
wire            n16718;
wire            n16719;
wire            n1672;
wire            n16720;
wire            n16721;
wire            n16722;
wire            n16723;
wire            n16724;
wire            n16725;
wire            n16726;
wire            n16727;
wire            n16728;
wire            n16729;
wire            n1673;
wire            n16730;
wire            n16731;
wire            n16732;
wire            n16733;
wire            n16734;
wire            n16735;
wire            n16736;
wire            n16737;
wire            n16738;
wire            n16739;
wire            n1674;
wire            n16740;
wire            n16741;
wire            n16742;
wire            n16743;
wire            n16744;
wire            n16745;
wire            n16746;
wire            n16747;
wire            n16748;
wire            n16749;
wire            n1675;
wire            n16750;
wire            n16751;
wire            n16752;
wire            n16753;
wire            n16754;
wire            n16755;
wire            n16756;
wire            n16757;
wire            n16758;
wire            n16759;
wire            n1676;
wire            n16760;
wire            n16761;
wire            n16762;
wire            n16763;
wire            n16764;
wire            n16765;
wire            n16766;
wire            n16767;
wire            n16768;
wire            n16769;
wire            n1677;
wire            n16770;
wire            n16771;
wire            n16772;
wire            n16773;
wire            n16774;
wire            n16775;
wire            n16776;
wire            n16777;
wire            n16778;
wire            n16779;
wire            n1678;
wire            n16780;
wire            n16781;
wire            n16782;
wire            n16783;
wire            n16784;
wire            n16785;
wire            n16786;
wire            n16787;
wire            n16788;
wire     [13:0] n16789;
wire            n1679;
wire            n16790;
wire            n16791;
wire            n16792;
wire            n16793;
wire            n16794;
wire            n16795;
wire            n16796;
wire            n16797;
wire            n16798;
wire            n16799;
wire            n168;
wire            n1680;
wire            n16800;
wire            n16801;
wire            n16802;
wire            n16803;
wire            n16804;
wire            n16805;
wire            n16806;
wire            n16807;
wire            n16808;
wire            n16809;
wire            n1681;
wire            n16810;
wire            n16811;
wire            n16812;
wire            n16813;
wire            n16814;
wire            n16815;
wire            n16816;
wire            n16817;
wire            n16818;
wire            n16819;
wire            n1682;
wire            n16820;
wire            n16821;
wire            n16822;
wire            n16823;
wire            n16824;
wire            n16825;
wire            n16826;
wire            n16827;
wire            n16828;
wire            n16829;
wire            n1683;
wire            n16830;
wire            n16831;
wire            n16832;
wire            n16833;
wire            n16834;
wire            n16835;
wire            n16836;
wire            n16837;
wire            n16838;
wire            n16839;
wire            n1684;
wire            n16840;
wire            n16841;
wire            n16842;
wire            n16843;
wire            n16844;
wire            n16845;
wire            n16846;
wire            n16847;
wire            n16848;
wire            n16849;
wire            n1685;
wire            n16850;
wire            n16851;
wire            n16852;
wire            n16853;
wire            n16854;
wire            n16855;
wire     [14:0] n16856;
wire            n16857;
wire            n16858;
wire            n16859;
wire            n1686;
wire            n16860;
wire            n16861;
wire            n16862;
wire            n16863;
wire            n16864;
wire            n16865;
wire            n16866;
wire            n16867;
wire            n16868;
wire            n16869;
wire            n1687;
wire            n16870;
wire            n16871;
wire            n16872;
wire            n16873;
wire            n16874;
wire            n16875;
wire            n16876;
wire            n16877;
wire            n16878;
wire            n16879;
wire            n1688;
wire            n16880;
wire            n16881;
wire            n16882;
wire            n16883;
wire            n16884;
wire            n16885;
wire            n16886;
wire            n16887;
wire            n16888;
wire            n16889;
wire            n1689;
wire            n16890;
wire            n16891;
wire            n16892;
wire            n16893;
wire            n16894;
wire            n16895;
wire            n16896;
wire            n16897;
wire            n16898;
wire            n16899;
wire            n169;
wire            n1690;
wire            n16900;
wire            n16901;
wire            n16902;
wire            n16903;
wire            n16904;
wire            n16905;
wire            n16906;
wire            n16907;
wire            n16908;
wire            n16909;
wire            n1691;
wire            n16910;
wire            n16911;
wire            n16912;
wire            n16913;
wire            n16914;
wire            n16915;
wire            n16916;
wire            n16917;
wire            n16918;
wire            n16919;
wire            n1692;
wire            n16920;
wire            n16921;
wire            n16922;
wire            n16923;
wire            n16924;
wire            n16925;
wire            n16926;
wire            n16927;
wire            n16928;
wire            n16929;
wire            n1693;
wire            n16930;
wire            n16931;
wire            n16932;
wire            n16933;
wire     [15:0] n16934;
wire            n16935;
wire            n16936;
wire            n16937;
wire            n16938;
wire            n16939;
wire            n1694;
wire            n16940;
wire            n16941;
wire            n16942;
wire            n16943;
wire            n16944;
wire            n16945;
wire            n16946;
wire            n16947;
wire            n16948;
wire            n16949;
wire            n1695;
wire            n16950;
wire            n16951;
wire            n16952;
wire            n16953;
wire            n16954;
wire            n16955;
wire            n16956;
wire            n16957;
wire            n16958;
wire            n16959;
wire            n1696;
wire            n16960;
wire            n16961;
wire            n16962;
wire            n16963;
wire            n16964;
wire            n16965;
wire            n16966;
wire            n16967;
wire            n16968;
wire            n16969;
wire            n1697;
wire            n16970;
wire            n16971;
wire            n16972;
wire            n16973;
wire            n16974;
wire            n16975;
wire            n16976;
wire            n16977;
wire            n16978;
wire            n16979;
wire            n1698;
wire            n16980;
wire            n16981;
wire            n16982;
wire            n16983;
wire            n16984;
wire            n16985;
wire            n16986;
wire            n16987;
wire            n16988;
wire            n16989;
wire            n1699;
wire            n16990;
wire            n16991;
wire            n16992;
wire            n16993;
wire            n16994;
wire            n16995;
wire            n16996;
wire            n16997;
wire            n16998;
wire            n16999;
wire            n17;
wire            n170;
wire            n1700;
wire            n17000;
wire            n17001;
wire     [16:0] n17002;
wire            n17003;
wire            n17004;
wire            n17005;
wire            n17006;
wire            n17007;
wire            n17008;
wire            n17009;
wire            n1701;
wire            n17010;
wire            n17011;
wire            n17012;
wire            n17013;
wire            n17014;
wire            n17015;
wire            n17016;
wire            n17017;
wire            n17018;
wire            n17019;
wire            n1702;
wire            n17020;
wire            n17021;
wire            n17022;
wire            n17023;
wire            n17024;
wire            n17025;
wire            n17026;
wire            n17027;
wire            n17028;
wire            n17029;
wire            n1703;
wire            n17030;
wire            n17031;
wire            n17032;
wire            n17033;
wire            n17034;
wire            n17035;
wire            n17036;
wire            n17037;
wire            n17038;
wire            n17039;
wire            n1704;
wire            n17040;
wire            n17041;
wire            n17042;
wire            n17043;
wire            n17044;
wire            n17045;
wire            n17046;
wire            n17047;
wire            n17048;
wire            n17049;
wire            n1705;
wire            n17050;
wire            n17051;
wire            n17052;
wire            n17053;
wire            n17054;
wire            n17055;
wire            n17056;
wire            n17057;
wire            n17058;
wire            n17059;
wire            n1706;
wire            n17060;
wire            n17061;
wire            n17062;
wire            n17063;
wire            n17064;
wire            n17065;
wire            n17066;
wire            n17067;
wire            n17068;
wire            n17069;
wire            n1707;
wire            n17070;
wire            n17071;
wire            n17072;
wire            n17073;
wire     [17:0] n17074;
wire            n17075;
wire            n17076;
wire            n17077;
wire            n17078;
wire            n17079;
wire            n1708;
wire            n17080;
wire            n17081;
wire            n17082;
wire            n17083;
wire            n17084;
wire            n17085;
wire            n17086;
wire            n17087;
wire            n17088;
wire            n17089;
wire            n1709;
wire            n17090;
wire            n17091;
wire            n17092;
wire            n17093;
wire            n17094;
wire            n17095;
wire            n17096;
wire            n17097;
wire            n17098;
wire            n17099;
wire            n171;
wire            n1710;
wire            n17100;
wire            n17101;
wire            n17102;
wire            n17103;
wire            n17104;
wire            n17105;
wire            n17106;
wire            n17107;
wire            n17108;
wire            n17109;
wire            n1711;
wire            n17110;
wire            n17111;
wire            n17112;
wire            n17113;
wire            n17114;
wire            n17115;
wire            n17116;
wire            n17117;
wire            n17118;
wire            n17119;
wire            n1712;
wire            n17120;
wire            n17121;
wire            n17122;
wire            n17123;
wire            n17124;
wire            n17125;
wire            n17126;
wire            n17127;
wire            n17128;
wire            n17129;
wire            n1713;
wire            n17130;
wire            n17131;
wire     [18:0] n17132;
wire            n17133;
wire            n17134;
wire            n17135;
wire            n17136;
wire            n17137;
wire            n17138;
wire            n17139;
wire            n1714;
wire            n17140;
wire            n17141;
wire            n17142;
wire            n17143;
wire            n17144;
wire            n17145;
wire            n17146;
wire            n17147;
wire            n17148;
wire            n17149;
wire            n1715;
wire            n17150;
wire            n17151;
wire            n17152;
wire            n17153;
wire            n17154;
wire            n17155;
wire            n17156;
wire            n17157;
wire            n17158;
wire            n17159;
wire            n1716;
wire            n17160;
wire            n17161;
wire            n17162;
wire            n17163;
wire            n17164;
wire            n17165;
wire            n17166;
wire            n17167;
wire            n17168;
wire            n17169;
wire            n1717;
wire            n17170;
wire            n17171;
wire            n17172;
wire            n17173;
wire            n17174;
wire            n17175;
wire            n17176;
wire            n17177;
wire            n17178;
wire            n17179;
wire            n1718;
wire            n17180;
wire            n17181;
wire            n17182;
wire            n17183;
wire            n17184;
wire            n17185;
wire            n17186;
wire            n17187;
wire            n17188;
wire            n17189;
wire            n1719;
wire            n17190;
wire            n17191;
wire            n17192;
wire            n17193;
wire            n17194;
wire     [19:0] n17195;
wire            n17196;
wire            n17197;
wire            n17198;
wire            n17199;
wire            n172;
wire            n1720;
wire            n17200;
wire            n17201;
wire            n17202;
wire            n17203;
wire            n17204;
wire            n17205;
wire            n17206;
wire            n17207;
wire            n17208;
wire            n17209;
wire            n1721;
wire            n17210;
wire            n17211;
wire            n17212;
wire            n17213;
wire            n17214;
wire            n17215;
wire            n17216;
wire            n17217;
wire            n17218;
wire            n17219;
wire            n1722;
wire            n17220;
wire            n17221;
wire            n17222;
wire            n17223;
wire            n17224;
wire            n17225;
wire            n17226;
wire            n17227;
wire            n17228;
wire            n17229;
wire            n1723;
wire            n17230;
wire            n17231;
wire            n17232;
wire            n17233;
wire            n17234;
wire            n17235;
wire            n17236;
wire            n17237;
wire            n17238;
wire            n17239;
wire            n1724;
wire            n17240;
wire            n17241;
wire            n17242;
wire            n17243;
wire            n17244;
wire            n17245;
wire            n17246;
wire            n17247;
wire            n17248;
wire            n17249;
wire            n1725;
wire            n17250;
wire     [20:0] n17251;
wire            n17252;
wire            n17253;
wire            n17254;
wire            n17255;
wire            n17256;
wire            n17257;
wire            n17258;
wire            n17259;
wire            n1726;
wire            n17260;
wire            n17261;
wire            n17262;
wire            n17263;
wire            n17264;
wire            n17265;
wire            n17266;
wire            n17267;
wire            n17268;
wire            n17269;
wire            n1727;
wire            n17270;
wire            n17271;
wire            n17272;
wire            n17273;
wire            n17274;
wire            n17275;
wire            n17276;
wire            n17277;
wire            n17278;
wire            n17279;
wire            n1728;
wire            n17280;
wire            n17281;
wire            n17282;
wire            n17283;
wire            n17284;
wire            n17285;
wire            n17286;
wire            n17287;
wire            n17288;
wire            n17289;
wire            n1729;
wire            n17290;
wire            n17291;
wire            n17292;
wire            n17293;
wire            n17294;
wire            n17295;
wire            n17296;
wire            n17297;
wire            n17298;
wire            n17299;
wire            n173;
wire            n1730;
wire            n17300;
wire            n17301;
wire            n17302;
wire            n17303;
wire            n17304;
wire            n17305;
wire            n17306;
wire     [21:0] n17307;
wire            n17308;
wire            n17309;
wire            n1731;
wire            n17310;
wire            n17311;
wire            n17312;
wire            n17313;
wire            n17314;
wire            n17315;
wire            n17316;
wire            n17317;
wire            n17318;
wire            n17319;
wire            n1732;
wire            n17320;
wire            n17321;
wire            n17322;
wire            n17323;
wire            n17324;
wire            n17325;
wire            n17326;
wire            n17327;
wire            n17328;
wire            n17329;
wire            n1733;
wire            n17330;
wire            n17331;
wire            n17332;
wire            n17333;
wire            n17334;
wire            n17335;
wire            n17336;
wire            n17337;
wire            n17338;
wire            n17339;
wire            n1734;
wire            n17340;
wire            n17341;
wire            n17342;
wire            n17343;
wire            n17344;
wire            n17345;
wire            n17346;
wire            n17347;
wire            n17348;
wire     [22:0] n17349;
wire            n1735;
wire            n17350;
wire            n17351;
wire            n17352;
wire            n17353;
wire            n17354;
wire            n17355;
wire            n17356;
wire            n17357;
wire            n17358;
wire            n17359;
wire            n1736;
wire            n17360;
wire            n17361;
wire            n17362;
wire            n17363;
wire            n17364;
wire            n17365;
wire            n17366;
wire            n17367;
wire            n17368;
wire            n17369;
wire            n1737;
wire            n17370;
wire            n17371;
wire            n17372;
wire            n17373;
wire            n17374;
wire            n17375;
wire            n17376;
wire            n17377;
wire            n17378;
wire            n17379;
wire            n1738;
wire            n17380;
wire            n17381;
wire            n17382;
wire            n17383;
wire            n17384;
wire            n17385;
wire            n17386;
wire            n17387;
wire            n17388;
wire     [23:0] n17389;
wire            n1739;
wire            n17390;
wire            n17391;
wire            n17392;
wire            n17393;
wire            n17394;
wire            n17395;
wire            n17396;
wire            n17397;
wire            n17398;
wire            n17399;
wire            n174;
wire            n1740;
wire            n17400;
wire            n17401;
wire            n17402;
wire            n17403;
wire            n17404;
wire            n17405;
wire            n17406;
wire            n17407;
wire            n17408;
wire            n17409;
wire            n1741;
wire            n17410;
wire            n17411;
wire            n17412;
wire            n17413;
wire            n17414;
wire            n17415;
wire            n17416;
wire            n17417;
wire            n17418;
wire            n17419;
wire            n1742;
wire            n17420;
wire            n17421;
wire            n17422;
wire            n17423;
wire     [24:0] n17424;
wire            n17425;
wire            n17426;
wire            n17427;
wire            n17428;
wire            n17429;
wire            n1743;
wire            n17430;
wire            n17431;
wire            n17432;
wire            n17433;
wire            n17434;
wire            n17435;
wire            n17436;
wire            n17437;
wire            n17438;
wire            n17439;
wire            n1744;
wire            n17440;
wire            n17441;
wire            n17442;
wire            n17443;
wire            n17444;
wire            n17445;
wire            n17446;
wire            n17447;
wire            n17448;
wire            n17449;
wire            n1745;
wire            n17450;
wire            n17451;
wire            n17452;
wire            n17453;
wire            n17454;
wire            n17455;
wire            n17456;
wire            n17457;
wire     [25:0] n17458;
wire            n17459;
wire            n1746;
wire            n17460;
wire            n17461;
wire            n17462;
wire            n17463;
wire            n17464;
wire            n17465;
wire            n17466;
wire            n17467;
wire            n17468;
wire            n17469;
wire            n1747;
wire            n17470;
wire            n17471;
wire            n17472;
wire            n17473;
wire            n17474;
wire            n17475;
wire            n17476;
wire     [26:0] n17477;
wire            n17478;
wire            n17479;
wire            n1748;
wire            n17480;
wire            n17481;
wire            n17482;
wire            n17483;
wire            n17484;
wire            n17485;
wire            n17486;
wire            n17487;
wire            n17488;
wire            n17489;
wire            n1749;
wire            n17490;
wire            n17491;
wire            n17492;
wire            n17493;
wire            n17494;
wire            n17495;
wire            n17496;
wire            n17497;
wire            n17498;
wire            n17499;
wire            n175;
wire            n1750;
wire            n17500;
wire            n17501;
wire            n17502;
wire            n17503;
wire            n17504;
wire            n17505;
wire            n17506;
wire            n17507;
wire            n17508;
wire            n17509;
wire            n1751;
wire            n17510;
wire     [27:0] n17511;
wire            n17512;
wire            n17513;
wire            n17514;
wire            n17515;
wire            n17516;
wire            n17517;
wire            n17518;
wire            n17519;
wire            n1752;
wire            n17520;
wire            n17521;
wire            n17522;
wire            n17523;
wire            n17524;
wire     [28:0] n17525;
wire            n17526;
wire            n17527;
wire            n17528;
wire            n17529;
wire            n1753;
wire            n17530;
wire            n17531;
wire            n17532;
wire            n17533;
wire            n17534;
wire            n17535;
wire            n17536;
wire            n17537;
wire            n17538;
wire            n17539;
wire            n1754;
wire            n17540;
wire            n17541;
wire            n17542;
wire            n17543;
wire            n17544;
wire            n17545;
wire            n17546;
wire            n17547;
wire            n17548;
wire            n17549;
wire            n1755;
wire            n17550;
wire            n17551;
wire            n17552;
wire            n17553;
wire     [29:0] n17554;
wire            n17555;
wire            n17556;
wire            n17557;
wire            n17558;
wire            n17559;
wire            n1756;
wire            n17560;
wire            n17561;
wire            n17562;
wire            n17563;
wire            n17564;
wire            n17565;
wire            n17566;
wire     [30:0] n17567;
wire            n17568;
wire            n17569;
wire            n1757;
wire            n17570;
wire            n17571;
wire            n17572;
wire     [31:0] n17573;
wire            n1758;
wire            n1759;
wire            n176;
wire            n1760;
wire            n1761;
wire            n1762;
wire            n1763;
wire            n1764;
wire            n1765;
wire            n1766;
wire            n1767;
wire            n1768;
wire            n1769;
wire            n177;
wire            n1770;
wire            n1771;
wire            n1772;
wire            n1773;
wire            n1774;
wire            n1775;
wire            n1776;
wire            n1777;
wire            n1778;
wire            n1779;
wire            n178;
wire            n1780;
wire            n1781;
wire            n1782;
wire            n1783;
wire            n1784;
wire            n1785;
wire            n1786;
wire            n1787;
wire            n1788;
wire            n1789;
wire            n179;
wire            n1790;
wire            n1791;
wire            n1792;
wire            n1793;
wire            n1794;
wire            n1795;
wire            n1796;
wire            n1797;
wire            n1798;
wire            n1799;
wire            n18;
wire            n180;
wire            n1800;
wire            n1801;
wire            n1802;
wire            n1803;
wire            n1804;
wire            n1805;
wire            n1806;
wire            n1807;
wire            n1808;
wire            n1809;
wire            n181;
wire            n1810;
wire            n1811;
wire            n1812;
wire            n1813;
wire            n1814;
wire            n1815;
wire            n1816;
wire            n1817;
wire            n1818;
wire            n1819;
wire            n182;
wire            n1820;
wire            n1821;
wire            n1822;
wire            n1823;
wire            n1824;
wire            n1825;
wire            n1826;
wire            n1827;
wire            n1828;
wire            n1829;
wire            n183;
wire            n1830;
wire            n1831;
wire            n1832;
wire            n1833;
wire            n1834;
wire            n1835;
wire            n1836;
wire            n1837;
wire            n1838;
wire            n1839;
wire            n184;
wire            n1840;
wire            n1841;
wire            n1842;
wire            n1843;
wire            n1844;
wire            n1845;
wire            n1846;
wire            n1847;
wire            n1848;
wire            n1849;
wire            n185;
wire            n1850;
wire            n1851;
wire            n1852;
wire            n1853;
wire            n1854;
wire            n1855;
wire            n1856;
wire            n1857;
wire            n1858;
wire            n1859;
wire            n186;
wire            n1860;
wire            n1861;
wire            n1862;
wire            n1863;
wire            n1864;
wire            n1865;
wire            n1866;
wire            n1867;
wire            n1868;
wire            n1869;
wire            n187;
wire            n1870;
wire            n1871;
wire            n1872;
wire            n1873;
wire            n1874;
wire            n1875;
wire            n1876;
wire            n1877;
wire            n1878;
wire            n1879;
wire            n188;
wire            n1880;
wire            n1881;
wire            n1882;
wire            n1883;
wire            n1884;
wire            n1885;
wire            n1886;
wire            n1887;
wire            n1888;
wire            n1889;
wire            n189;
wire            n1890;
wire            n1891;
wire            n1892;
wire            n1893;
wire            n1894;
wire            n1895;
wire            n1896;
wire            n1897;
wire            n1898;
wire            n1899;
wire            n19;
wire            n190;
wire            n1900;
wire            n1901;
wire            n1902;
wire            n1903;
wire            n1904;
wire            n1905;
wire            n1906;
wire            n1907;
wire            n1908;
wire            n1909;
wire            n191;
wire            n1910;
wire            n1911;
wire            n1912;
wire            n1913;
wire            n1914;
wire            n1915;
wire            n1916;
wire            n1917;
wire            n1918;
wire            n1919;
wire            n192;
wire            n1920;
wire            n1921;
wire            n1922;
wire            n1923;
wire            n1924;
wire            n1925;
wire            n1926;
wire            n1927;
wire            n1928;
wire            n1929;
wire            n193;
wire            n1930;
wire            n1931;
wire            n1932;
wire            n1933;
wire            n1934;
wire            n1935;
wire            n1936;
wire            n1937;
wire            n1938;
wire            n1939;
wire            n194;
wire            n1940;
wire            n1941;
wire            n1942;
wire            n1943;
wire            n1944;
wire            n1945;
wire            n1946;
wire            n1947;
wire            n1948;
wire            n1949;
wire            n195;
wire            n1950;
wire            n1951;
wire            n1952;
wire            n1953;
wire            n1954;
wire            n1955;
wire            n1956;
wire            n1957;
wire            n1958;
wire            n1959;
wire            n196;
wire            n1960;
wire            n1961;
wire            n1962;
wire            n1963;
wire            n1964;
wire            n1965;
wire            n1966;
wire            n1967;
wire            n1968;
wire            n1969;
wire            n197;
wire            n1970;
wire            n1971;
wire            n1972;
wire            n1973;
wire            n1974;
wire            n1975;
wire            n1976;
wire            n1977;
wire            n1978;
wire            n1979;
wire            n198;
wire            n1980;
wire            n1981;
wire            n1982;
wire            n1983;
wire            n1984;
wire            n1985;
wire            n1986;
wire            n1987;
wire            n1988;
wire            n1989;
wire            n199;
wire            n1990;
wire            n1991;
wire            n1992;
wire            n1993;
wire            n1994;
wire            n1995;
wire            n1996;
wire            n1997;
wire            n1998;
wire            n1999;
wire            n20;
wire            n200;
wire            n2000;
wire            n2001;
wire            n2002;
wire            n2003;
wire            n2004;
wire            n2005;
wire            n2006;
wire            n2007;
wire            n2008;
wire            n2009;
wire            n201;
wire            n2010;
wire            n2011;
wire            n2012;
wire            n2013;
wire            n2014;
wire            n2015;
wire            n2016;
wire            n2017;
wire            n2018;
wire            n2019;
wire            n202;
wire            n2020;
wire            n2021;
wire            n2022;
wire            n2023;
wire            n2024;
wire            n2025;
wire            n2026;
wire            n2027;
wire            n2028;
wire            n2029;
wire            n203;
wire            n2030;
wire            n2031;
wire            n2032;
wire            n2033;
wire            n2034;
wire            n2035;
wire            n2036;
wire            n2037;
wire            n2038;
wire            n2039;
wire            n204;
wire            n2040;
wire            n2041;
wire            n2042;
wire            n2043;
wire            n2044;
wire            n2045;
wire            n2046;
wire            n2047;
wire            n2048;
wire            n2049;
wire            n205;
wire            n2050;
wire            n2051;
wire            n2052;
wire            n2053;
wire            n2054;
wire            n2055;
wire            n2056;
wire            n2057;
wire            n2058;
wire            n2059;
wire            n206;
wire            n2060;
wire            n2061;
wire            n2062;
wire            n2063;
wire            n2064;
wire            n2065;
wire            n2066;
wire            n2067;
wire            n2068;
wire            n2069;
wire            n207;
wire            n2070;
wire            n2071;
wire            n2072;
wire            n2073;
wire            n2074;
wire            n2075;
wire            n2076;
wire            n2077;
wire            n2078;
wire            n2079;
wire            n208;
wire            n2080;
wire            n2081;
wire            n2082;
wire            n2083;
wire            n2084;
wire            n2085;
wire            n2086;
wire            n2087;
wire            n2088;
wire            n2089;
wire            n209;
wire            n2090;
wire            n2091;
wire            n2092;
wire            n2093;
wire            n2094;
wire            n2095;
wire            n2096;
wire            n2097;
wire            n2098;
wire            n2099;
wire            n21;
wire            n210;
wire            n2100;
wire            n2101;
wire            n2102;
wire            n2103;
wire            n2104;
wire            n2105;
wire            n2106;
wire            n2107;
wire            n2108;
wire            n2109;
wire            n211;
wire            n2110;
wire            n2111;
wire            n2112;
wire            n2113;
wire            n2114;
wire            n2115;
wire            n2116;
wire            n2117;
wire            n2118;
wire            n2119;
wire            n212;
wire            n2120;
wire            n2121;
wire            n2122;
wire            n2123;
wire            n2124;
wire            n2125;
wire            n2126;
wire            n2127;
wire            n2128;
wire            n2129;
wire            n213;
wire            n2130;
wire            n2131;
wire            n2132;
wire            n2133;
wire            n2134;
wire            n2135;
wire            n2136;
wire            n2137;
wire            n2138;
wire            n2139;
wire            n214;
wire            n2140;
wire            n2141;
wire            n2142;
wire            n2143;
wire            n2144;
wire            n2145;
wire            n2146;
wire            n2147;
wire            n2148;
wire            n2149;
wire            n215;
wire            n2150;
wire            n2151;
wire            n2152;
wire            n2153;
wire            n2154;
wire            n2155;
wire            n2156;
wire            n2157;
wire            n2158;
wire            n2159;
wire            n216;
wire            n2160;
wire            n2161;
wire            n2162;
wire            n2163;
wire            n2164;
wire            n2165;
wire            n2166;
wire            n2167;
wire            n2168;
wire            n2169;
wire            n217;
wire            n2170;
wire            n2171;
wire            n2172;
wire            n2173;
wire            n2174;
wire            n2175;
wire            n2176;
wire            n2177;
wire            n2178;
wire            n2179;
wire            n218;
wire            n2180;
wire            n2181;
wire            n2182;
wire            n2183;
wire            n2184;
wire            n2185;
wire            n2186;
wire            n2187;
wire            n2188;
wire            n2189;
wire            n219;
wire            n2190;
wire            n2191;
wire            n2192;
wire            n2193;
wire            n2194;
wire            n2195;
wire            n2196;
wire            n2197;
wire            n2198;
wire            n2199;
wire            n22;
wire            n220;
wire            n2200;
wire            n2201;
wire            n2202;
wire            n2203;
wire            n2204;
wire            n2205;
wire            n2206;
wire            n2207;
wire            n2208;
wire            n2209;
wire            n221;
wire            n2210;
wire            n2211;
wire            n2212;
wire            n2213;
wire            n2214;
wire            n2215;
wire            n2216;
wire            n2217;
wire            n2218;
wire            n2219;
wire            n222;
wire            n2220;
wire            n2221;
wire            n2222;
wire            n2223;
wire            n2224;
wire            n2225;
wire            n2226;
wire            n2227;
wire            n2228;
wire            n2229;
wire            n223;
wire            n2230;
wire            n2231;
wire            n2232;
wire            n2233;
wire            n2234;
wire            n2235;
wire            n2236;
wire            n2237;
wire            n2238;
wire            n2239;
wire            n224;
wire            n2240;
wire            n2241;
wire            n2242;
wire            n2243;
wire            n2244;
wire            n2245;
wire            n2246;
wire            n2247;
wire            n2248;
wire            n2249;
wire            n225;
wire            n2250;
wire            n2251;
wire            n2252;
wire            n2253;
wire            n2254;
wire            n2255;
wire            n2256;
wire            n2257;
wire            n2258;
wire            n2259;
wire            n226;
wire            n2260;
wire            n2261;
wire            n2262;
wire            n2263;
wire            n2264;
wire            n2265;
wire            n2266;
wire            n2267;
wire            n2268;
wire            n2269;
wire            n227;
wire            n2270;
wire            n2271;
wire            n2272;
wire            n2273;
wire            n2274;
wire            n2275;
wire            n2276;
wire            n2277;
wire            n2278;
wire            n2279;
wire            n228;
wire            n2280;
wire            n2281;
wire            n2282;
wire            n2283;
wire            n2284;
wire            n2285;
wire            n2286;
wire            n2287;
wire            n2288;
wire            n2289;
wire            n229;
wire            n2290;
wire            n2291;
wire            n2292;
wire            n2293;
wire            n2294;
wire            n2295;
wire            n2296;
wire            n2297;
wire            n2298;
wire            n2299;
wire            n23;
wire            n230;
wire            n2300;
wire            n2301;
wire            n2302;
wire            n2303;
wire            n2304;
wire            n2305;
wire            n2306;
wire            n2307;
wire            n2308;
wire            n2309;
wire            n231;
wire            n2310;
wire            n2311;
wire            n2312;
wire            n2313;
wire            n2314;
wire            n2315;
wire            n2316;
wire            n2317;
wire            n2318;
wire            n2319;
wire            n232;
wire            n2320;
wire            n2321;
wire            n2322;
wire            n2323;
wire            n2324;
wire            n2325;
wire            n2326;
wire            n2327;
wire            n2328;
wire            n2329;
wire            n233;
wire            n2330;
wire            n2331;
wire            n2332;
wire            n2333;
wire            n2334;
wire            n2335;
wire            n2336;
wire            n2337;
wire            n2338;
wire            n2339;
wire            n234;
wire            n2340;
wire            n2341;
wire            n2342;
wire            n2343;
wire            n2344;
wire            n2345;
wire            n2346;
wire            n2347;
wire            n2348;
wire            n2349;
wire            n235;
wire            n2350;
wire            n2351;
wire            n2352;
wire            n2353;
wire            n2354;
wire            n2355;
wire            n2356;
wire            n2357;
wire            n2358;
wire            n2359;
wire            n236;
wire            n2360;
wire            n2361;
wire            n2362;
wire            n2363;
wire            n2364;
wire            n2365;
wire            n2366;
wire            n2367;
wire            n2368;
wire            n2369;
wire            n237;
wire            n2370;
wire            n2371;
wire            n2372;
wire            n2373;
wire            n2374;
wire            n2375;
wire            n2376;
wire            n2377;
wire            n2378;
wire            n2379;
wire            n238;
wire            n2380;
wire            n2381;
wire            n2382;
wire            n2383;
wire            n2384;
wire            n2385;
wire            n2386;
wire            n2387;
wire            n2388;
wire            n2389;
wire            n239;
wire            n2390;
wire            n2391;
wire            n2392;
wire            n2393;
wire            n2394;
wire            n2395;
wire            n2396;
wire            n2397;
wire            n2398;
wire            n2399;
wire            n24;
wire            n240;
wire            n2400;
wire            n2401;
wire            n2402;
wire            n2403;
wire            n2404;
wire            n2405;
wire            n2406;
wire            n2407;
wire            n2408;
wire            n2409;
wire            n241;
wire            n2410;
wire            n2411;
wire            n2412;
wire            n2413;
wire            n2414;
wire            n2415;
wire            n2416;
wire            n2417;
wire            n2418;
wire            n2419;
wire            n242;
wire            n2420;
wire            n2421;
wire            n2422;
wire            n2423;
wire            n2424;
wire            n2425;
wire            n2426;
wire            n2427;
wire            n2428;
wire            n2429;
wire            n243;
wire            n2430;
wire            n2431;
wire            n2432;
wire            n2433;
wire            n2434;
wire            n2435;
wire            n2436;
wire            n2437;
wire            n2438;
wire            n2439;
wire            n244;
wire            n2440;
wire            n2441;
wire            n2442;
wire            n2443;
wire            n2444;
wire            n2445;
wire            n2446;
wire            n2447;
wire            n2448;
wire            n2449;
wire            n245;
wire            n2450;
wire            n2451;
wire            n2452;
wire            n2453;
wire            n2454;
wire            n2455;
wire            n2456;
wire            n2457;
wire            n2458;
wire            n2459;
wire            n246;
wire            n2460;
wire            n2461;
wire            n2462;
wire            n2463;
wire            n2464;
wire            n2465;
wire            n2466;
wire            n2467;
wire            n2468;
wire            n2469;
wire            n247;
wire            n2470;
wire            n2471;
wire            n2472;
wire            n2473;
wire            n2474;
wire            n2475;
wire            n2476;
wire            n2477;
wire            n2478;
wire            n2479;
wire            n248;
wire            n2480;
wire            n2481;
wire            n2482;
wire            n2483;
wire            n2484;
wire            n2485;
wire            n2486;
wire            n2487;
wire            n2488;
wire            n2489;
wire            n249;
wire            n2490;
wire            n2491;
wire            n2492;
wire            n2493;
wire            n2494;
wire            n2495;
wire            n2496;
wire            n2497;
wire            n2498;
wire            n2499;
wire            n25;
wire            n250;
wire            n2500;
wire            n2501;
wire            n2502;
wire            n2503;
wire            n2504;
wire            n2505;
wire            n2506;
wire            n2507;
wire            n2508;
wire            n2509;
wire            n251;
wire            n2510;
wire            n2511;
wire            n2512;
wire            n2513;
wire            n2514;
wire            n2515;
wire            n2516;
wire            n2517;
wire            n2518;
wire            n2519;
wire            n252;
wire            n2520;
wire            n2521;
wire            n2522;
wire            n2523;
wire            n2524;
wire            n2525;
wire            n2526;
wire            n2527;
wire            n2528;
wire            n2529;
wire            n253;
wire            n2530;
wire            n2531;
wire            n2532;
wire            n2533;
wire            n2534;
wire            n2535;
wire            n2536;
wire            n2537;
wire            n2538;
wire            n2539;
wire            n254;
wire            n2540;
wire            n2541;
wire            n2542;
wire            n2543;
wire            n2544;
wire            n2545;
wire            n2546;
wire            n2547;
wire            n2548;
wire            n2549;
wire            n255;
wire            n2550;
wire            n2551;
wire            n2552;
wire            n2553;
wire            n2554;
wire            n2555;
wire            n2556;
wire            n2557;
wire            n2558;
wire            n2559;
wire            n256;
wire            n2560;
wire            n2561;
wire            n2562;
wire            n2563;
wire            n2564;
wire            n2565;
wire            n2566;
wire            n2567;
wire            n2568;
wire            n2569;
wire            n257;
wire            n2570;
wire            n2571;
wire            n2572;
wire            n2573;
wire            n2574;
wire            n2575;
wire            n2576;
wire            n2577;
wire            n2578;
wire            n2579;
wire            n258;
wire            n2580;
wire            n2581;
wire            n2582;
wire            n2583;
wire            n2584;
wire            n2585;
wire            n2586;
wire            n2587;
wire            n2588;
wire            n2589;
wire            n259;
wire            n2590;
wire            n2591;
wire            n2592;
wire            n2593;
wire            n2594;
wire            n2595;
wire            n2596;
wire            n2597;
wire            n2598;
wire            n2599;
wire            n26;
wire            n260;
wire            n2600;
wire            n2601;
wire            n2602;
wire            n2603;
wire            n2604;
wire            n2605;
wire            n2606;
wire            n2607;
wire            n2608;
wire            n2609;
wire            n261;
wire            n2610;
wire            n2611;
wire            n2612;
wire            n2613;
wire            n2614;
wire            n2615;
wire            n2616;
wire            n2617;
wire            n2618;
wire            n2619;
wire            n262;
wire            n2620;
wire            n2621;
wire            n2622;
wire            n2623;
wire            n2624;
wire            n2625;
wire            n2626;
wire            n2627;
wire            n2628;
wire            n2629;
wire            n263;
wire            n2630;
wire            n2631;
wire            n2632;
wire            n2633;
wire            n2634;
wire            n2635;
wire            n2636;
wire            n2637;
wire            n2638;
wire            n2639;
wire            n264;
wire            n2640;
wire            n2641;
wire            n2642;
wire            n2643;
wire            n2644;
wire            n2645;
wire            n2646;
wire            n2647;
wire            n2648;
wire            n2649;
wire            n265;
wire            n2650;
wire            n2651;
wire            n2652;
wire            n2653;
wire            n2654;
wire            n2655;
wire            n2656;
wire            n2657;
wire            n2658;
wire            n2659;
wire            n266;
wire            n2660;
wire            n2661;
wire            n2662;
wire            n2663;
wire            n2664;
wire            n2665;
wire            n2666;
wire            n2667;
wire            n2668;
wire            n2669;
wire            n267;
wire            n2670;
wire            n2671;
wire            n2672;
wire            n2673;
wire            n2674;
wire            n2675;
wire            n2676;
wire            n2677;
wire            n2678;
wire            n2679;
wire            n268;
wire            n2680;
wire            n2681;
wire            n2682;
wire            n2683;
wire            n2684;
wire            n2685;
wire            n2686;
wire            n2687;
wire            n2688;
wire            n2689;
wire            n269;
wire            n2690;
wire            n2691;
wire            n2692;
wire            n2693;
wire            n2694;
wire            n2695;
wire            n2696;
wire            n2697;
wire            n2698;
wire            n2699;
wire            n27;
wire            n270;
wire            n2700;
wire            n2701;
wire            n2702;
wire            n2703;
wire            n2704;
wire            n2705;
wire            n2706;
wire            n2707;
wire            n2708;
wire            n2709;
wire            n271;
wire            n2710;
wire            n2711;
wire            n2712;
wire            n2713;
wire            n2714;
wire            n2715;
wire            n2716;
wire            n2717;
wire            n2718;
wire            n2719;
wire            n272;
wire            n2720;
wire            n2721;
wire            n2722;
wire            n2723;
wire            n2724;
wire            n2725;
wire            n2726;
wire            n2727;
wire            n2728;
wire            n2729;
wire            n273;
wire            n2730;
wire            n2731;
wire            n2732;
wire            n2733;
wire            n2734;
wire            n2735;
wire            n2736;
wire            n2737;
wire            n2738;
wire            n2739;
wire            n274;
wire            n2740;
wire            n2741;
wire            n2742;
wire            n2743;
wire            n2744;
wire            n2745;
wire            n2746;
wire            n2747;
wire            n2748;
wire            n2749;
wire            n275;
wire            n2750;
wire            n2751;
wire            n2752;
wire            n2753;
wire            n2754;
wire            n2755;
wire            n2756;
wire            n2757;
wire            n2758;
wire            n2759;
wire            n276;
wire            n2760;
wire            n2761;
wire            n2762;
wire            n2763;
wire            n2764;
wire            n2765;
wire            n2766;
wire            n2767;
wire            n2768;
wire            n2769;
wire            n277;
wire            n2770;
wire            n2771;
wire            n2772;
wire            n2773;
wire            n2774;
wire            n2775;
wire            n2776;
wire            n2777;
wire            n2778;
wire            n2779;
wire            n278;
wire            n2780;
wire            n2781;
wire            n2782;
wire            n2783;
wire            n2784;
wire            n2785;
wire            n2786;
wire            n2787;
wire            n2788;
wire            n2789;
wire            n279;
wire            n2790;
wire            n2791;
wire            n2792;
wire            n2793;
wire            n2794;
wire            n2795;
wire            n2796;
wire            n2797;
wire            n2798;
wire            n2799;
wire            n28;
wire            n280;
wire            n2800;
wire            n2801;
wire            n2802;
wire            n2803;
wire            n2804;
wire            n2805;
wire            n2806;
wire            n2807;
wire            n2808;
wire            n2809;
wire            n281;
wire            n2810;
wire            n2811;
wire            n2812;
wire            n2813;
wire            n2814;
wire            n2815;
wire            n2816;
wire            n2817;
wire            n2818;
wire            n2819;
wire            n282;
wire            n2820;
wire            n2821;
wire            n2822;
wire            n2823;
wire            n2824;
wire            n2825;
wire            n2826;
wire            n2827;
wire            n2828;
wire            n2829;
wire            n283;
wire            n2830;
wire            n2831;
wire            n2832;
wire            n2833;
wire            n2834;
wire            n2835;
wire            n2836;
wire            n2837;
wire            n2838;
wire            n2839;
wire            n284;
wire            n2840;
wire            n2841;
wire            n2842;
wire            n2843;
wire            n2844;
wire            n2845;
wire            n2846;
wire            n2847;
wire            n2848;
wire            n2849;
wire            n285;
wire            n2850;
wire            n2851;
wire            n2852;
wire            n2853;
wire            n2854;
wire            n2855;
wire            n2856;
wire            n2857;
wire            n2858;
wire            n2859;
wire            n286;
wire            n2860;
wire            n2861;
wire            n2862;
wire            n2863;
wire            n2864;
wire            n2865;
wire            n2866;
wire            n2867;
wire            n2868;
wire            n2869;
wire            n287;
wire            n2870;
wire            n2871;
wire            n2872;
wire            n2873;
wire            n2874;
wire            n2875;
wire            n2876;
wire            n2877;
wire            n2878;
wire            n2879;
wire            n288;
wire            n2880;
wire            n2881;
wire            n2882;
wire            n2883;
wire            n2884;
wire            n2885;
wire            n2886;
wire            n2887;
wire            n2888;
wire            n2889;
wire            n289;
wire            n2890;
wire            n2891;
wire            n2892;
wire            n2893;
wire            n2894;
wire            n2895;
wire            n2896;
wire            n2897;
wire            n2898;
wire            n2899;
wire            n29;
wire            n290;
wire            n2900;
wire            n2901;
wire            n2902;
wire            n2903;
wire            n2904;
wire            n2905;
wire            n2906;
wire            n2907;
wire            n2908;
wire            n2909;
wire            n291;
wire            n2910;
wire            n2911;
wire            n2912;
wire            n2913;
wire            n2914;
wire            n2915;
wire            n2916;
wire            n2917;
wire            n2918;
wire            n2919;
wire            n292;
wire            n2920;
wire            n2921;
wire            n2922;
wire            n2923;
wire            n2924;
wire            n2925;
wire            n2926;
wire            n2927;
wire            n2928;
wire            n2929;
wire            n293;
wire            n2930;
wire            n2931;
wire            n2932;
wire            n2933;
wire            n2934;
wire            n2935;
wire            n2936;
wire            n2937;
wire            n2938;
wire            n2939;
wire            n294;
wire            n2940;
wire            n2941;
wire            n2942;
wire            n2943;
wire            n2944;
wire            n2945;
wire            n2946;
wire            n2947;
wire            n2948;
wire            n2949;
wire            n295;
wire            n2950;
wire            n2951;
wire            n2952;
wire            n2953;
wire            n2954;
wire            n2955;
wire            n2956;
wire            n2957;
wire            n2958;
wire            n2959;
wire            n296;
wire            n2960;
wire            n2961;
wire            n2962;
wire            n2963;
wire            n2964;
wire            n2965;
wire            n2966;
wire            n2967;
wire            n2968;
wire            n2969;
wire            n297;
wire            n2970;
wire            n2971;
wire            n2972;
wire            n2973;
wire            n2974;
wire            n2975;
wire            n2976;
wire            n2977;
wire            n2978;
wire            n2979;
wire            n298;
wire            n2980;
wire            n2981;
wire            n2982;
wire            n2983;
wire            n2984;
wire            n2985;
wire            n2986;
wire            n2987;
wire            n2988;
wire            n2989;
wire            n299;
wire            n2990;
wire            n2991;
wire            n2992;
wire            n2993;
wire            n2994;
wire            n2995;
wire            n2996;
wire            n2997;
wire            n2998;
wire            n2999;
wire            n3;
wire            n30;
wire            n300;
wire            n3000;
wire            n3001;
wire            n3002;
wire            n3003;
wire            n3004;
wire            n3005;
wire            n3006;
wire            n3007;
wire            n3008;
wire            n3009;
wire            n301;
wire            n3010;
wire            n3011;
wire            n3012;
wire            n3013;
wire            n3014;
wire            n3015;
wire            n3016;
wire            n3017;
wire            n3018;
wire            n3019;
wire            n302;
wire            n3020;
wire            n3021;
wire            n3022;
wire            n3023;
wire            n3024;
wire            n3025;
wire            n3026;
wire            n3027;
wire            n3028;
wire            n3029;
wire            n303;
wire            n3030;
wire            n3031;
wire            n3032;
wire            n3033;
wire            n3034;
wire            n3035;
wire            n3036;
wire            n3037;
wire            n3038;
wire            n3039;
wire            n304;
wire            n3040;
wire            n3041;
wire            n3042;
wire            n3043;
wire            n3044;
wire            n3045;
wire            n3046;
wire            n3047;
wire            n3048;
wire            n3049;
wire            n305;
wire            n3050;
wire            n3051;
wire            n3052;
wire            n3053;
wire            n3054;
wire            n3055;
wire            n3056;
wire            n3057;
wire            n3058;
wire            n3059;
wire            n306;
wire            n3060;
wire            n3061;
wire            n3062;
wire            n3063;
wire            n3064;
wire            n3065;
wire            n3066;
wire            n3067;
wire            n3068;
wire            n3069;
wire            n307;
wire            n3070;
wire            n3071;
wire            n3072;
wire            n3073;
wire            n3074;
wire            n3075;
wire            n3076;
wire            n3077;
wire            n3078;
wire            n3079;
wire            n308;
wire            n3080;
wire            n3081;
wire            n3082;
wire            n3083;
wire            n3084;
wire            n3085;
wire            n3086;
wire            n3087;
wire            n3088;
wire            n3089;
wire            n309;
wire            n3090;
wire            n3091;
wire            n3092;
wire            n3093;
wire            n3094;
wire            n3095;
wire            n3096;
wire            n3097;
wire            n3098;
wire            n3099;
wire            n31;
wire            n310;
wire            n3100;
wire            n3101;
wire            n3102;
wire            n3103;
wire            n3104;
wire            n3105;
wire            n3106;
wire            n3107;
wire            n3108;
wire            n3109;
wire            n311;
wire            n3110;
wire            n3111;
wire            n3112;
wire            n3113;
wire            n3114;
wire            n3115;
wire            n3116;
wire            n3117;
wire            n3118;
wire            n3119;
wire            n312;
wire            n3120;
wire            n3121;
wire            n3122;
wire            n3123;
wire            n3124;
wire            n3125;
wire            n3126;
wire            n3127;
wire            n3128;
wire            n3129;
wire            n313;
wire            n3130;
wire            n3131;
wire            n3132;
wire            n3133;
wire            n3134;
wire            n3135;
wire            n3136;
wire            n3137;
wire            n3138;
wire            n3139;
wire            n314;
wire            n3140;
wire            n3141;
wire            n3142;
wire            n3143;
wire            n3144;
wire            n3145;
wire            n3146;
wire            n3147;
wire            n3148;
wire            n3149;
wire            n315;
wire            n3150;
wire            n3151;
wire            n3152;
wire            n3153;
wire            n3154;
wire            n3155;
wire            n3156;
wire            n3157;
wire            n3158;
wire            n3159;
wire            n316;
wire            n3160;
wire            n3161;
wire            n3162;
wire            n3163;
wire            n3164;
wire            n3165;
wire            n3166;
wire            n3167;
wire            n3168;
wire            n3169;
wire            n317;
wire            n3170;
wire            n3171;
wire            n3172;
wire            n3173;
wire            n3174;
wire            n3175;
wire            n3176;
wire            n3177;
wire            n3178;
wire            n3179;
wire            n318;
wire            n3180;
wire            n3181;
wire            n3182;
wire            n3183;
wire            n3184;
wire            n3185;
wire            n3186;
wire            n3187;
wire            n3188;
wire            n3189;
wire            n319;
wire            n3190;
wire            n3191;
wire            n3192;
wire            n3193;
wire            n3194;
wire            n3195;
wire            n3196;
wire            n3197;
wire            n3198;
wire            n3199;
wire            n32;
wire            n320;
wire            n3200;
wire            n3201;
wire            n3202;
wire            n3203;
wire            n3204;
wire            n3205;
wire            n3206;
wire            n3207;
wire            n3208;
wire            n3209;
wire            n321;
wire            n3210;
wire            n3211;
wire            n3212;
wire            n3213;
wire            n3214;
wire            n3215;
wire            n3216;
wire            n3217;
wire            n3218;
wire            n3219;
wire            n322;
wire            n3220;
wire            n3221;
wire            n3222;
wire            n3223;
wire            n3224;
wire            n3225;
wire            n3226;
wire            n3227;
wire            n3228;
wire            n3229;
wire            n323;
wire            n3230;
wire            n3231;
wire            n3232;
wire            n3233;
wire            n3234;
wire            n3235;
wire            n3236;
wire            n3237;
wire            n3238;
wire            n3239;
wire            n324;
wire            n3240;
wire            n3241;
wire            n3242;
wire            n3243;
wire            n3244;
wire            n3245;
wire            n3246;
wire            n3247;
wire            n3248;
wire            n3249;
wire            n325;
wire            n3250;
wire            n3251;
wire            n3252;
wire            n3253;
wire            n3254;
wire            n3255;
wire            n3256;
wire            n3257;
wire            n3258;
wire            n3259;
wire            n326;
wire            n3260;
wire            n3261;
wire            n3262;
wire            n3263;
wire            n3264;
wire            n3265;
wire            n3266;
wire            n3267;
wire            n3268;
wire            n3269;
wire            n327;
wire            n3270;
wire            n3271;
wire            n3272;
wire            n3273;
wire            n3274;
wire            n3275;
wire            n3276;
wire            n3277;
wire            n3278;
wire            n3279;
wire            n328;
wire            n3280;
wire            n3281;
wire            n3282;
wire            n3283;
wire            n3284;
wire            n3285;
wire            n3286;
wire            n3287;
wire            n3288;
wire            n3289;
wire            n329;
wire            n3290;
wire            n3291;
wire            n3292;
wire            n3293;
wire            n3294;
wire            n3295;
wire            n3296;
wire            n3297;
wire            n3298;
wire            n3299;
wire            n33;
wire            n330;
wire            n3300;
wire            n3301;
wire            n3302;
wire            n3303;
wire            n3304;
wire            n3305;
wire            n3306;
wire            n3307;
wire            n3308;
wire            n3309;
wire            n331;
wire            n3310;
wire            n3311;
wire            n3312;
wire            n3313;
wire            n3314;
wire            n3315;
wire            n3316;
wire            n3317;
wire            n3318;
wire            n3319;
wire            n332;
wire            n3320;
wire            n3321;
wire            n3322;
wire            n3323;
wire            n3324;
wire            n3325;
wire            n3326;
wire            n3327;
wire            n3328;
wire            n3329;
wire            n333;
wire            n3330;
wire            n3331;
wire            n3332;
wire            n3333;
wire            n3334;
wire            n3335;
wire            n3336;
wire            n3337;
wire            n3338;
wire            n3339;
wire            n334;
wire            n3340;
wire            n3341;
wire            n3342;
wire            n3343;
wire            n3344;
wire            n3345;
wire            n3346;
wire            n3347;
wire            n3348;
wire            n3349;
wire            n335;
wire            n3350;
wire            n3351;
wire            n3352;
wire            n3353;
wire            n3354;
wire            n3355;
wire            n3356;
wire            n3357;
wire            n3358;
wire            n3359;
wire            n336;
wire            n3360;
wire            n3361;
wire            n3362;
wire            n3363;
wire            n3364;
wire            n3365;
wire            n3366;
wire            n3367;
wire            n3368;
wire            n3369;
wire            n337;
wire            n3370;
wire            n3371;
wire            n3372;
wire            n3373;
wire            n3374;
wire            n3375;
wire            n3376;
wire            n3377;
wire            n3378;
wire            n3379;
wire            n338;
wire            n3380;
wire            n3381;
wire            n3382;
wire            n3383;
wire            n3384;
wire            n3385;
wire            n3386;
wire            n3387;
wire            n3388;
wire            n3389;
wire            n339;
wire            n3390;
wire            n3391;
wire            n3392;
wire            n3393;
wire            n3394;
wire            n3395;
wire            n3396;
wire            n3397;
wire            n3398;
wire            n3399;
wire            n34;
wire            n340;
wire            n3400;
wire            n3401;
wire            n3402;
wire            n3403;
wire            n3404;
wire            n3405;
wire            n3406;
wire            n3407;
wire            n3408;
wire            n3409;
wire            n341;
wire            n3410;
wire            n3411;
wire            n3412;
wire            n3413;
wire            n3414;
wire            n3415;
wire            n3416;
wire            n3417;
wire            n3418;
wire            n3419;
wire            n342;
wire            n3420;
wire            n3421;
wire            n3422;
wire            n3423;
wire            n3424;
wire            n3425;
wire            n3426;
wire            n3427;
wire            n3428;
wire            n3429;
wire            n343;
wire            n3430;
wire            n3431;
wire            n3432;
wire            n3433;
wire            n3434;
wire            n3435;
wire            n3436;
wire            n3437;
wire            n3438;
wire            n3439;
wire            n344;
wire            n3440;
wire            n3441;
wire            n3442;
wire            n3443;
wire            n3444;
wire            n3445;
wire            n3446;
wire            n3447;
wire            n3448;
wire            n3449;
wire            n345;
wire            n3450;
wire            n3451;
wire            n3452;
wire            n3453;
wire            n3454;
wire            n3455;
wire            n3456;
wire            n3457;
wire            n3458;
wire            n3459;
wire            n346;
wire            n3460;
wire            n3461;
wire            n3462;
wire            n3463;
wire            n3464;
wire            n3465;
wire            n3466;
wire            n3467;
wire            n3468;
wire            n3469;
wire            n347;
wire            n3470;
wire            n3471;
wire            n3472;
wire            n3473;
wire            n3474;
wire            n3475;
wire            n3476;
wire            n3477;
wire            n3478;
wire            n3479;
wire            n348;
wire            n3480;
wire            n3481;
wire            n3482;
wire            n3483;
wire            n3484;
wire            n3485;
wire            n3486;
wire            n3487;
wire            n3488;
wire            n3489;
wire            n349;
wire            n3490;
wire            n3491;
wire            n3492;
wire            n3493;
wire            n3494;
wire            n3495;
wire            n3496;
wire            n3497;
wire            n3498;
wire            n3499;
wire            n35;
wire            n350;
wire            n3500;
wire            n3501;
wire            n3502;
wire            n3503;
wire            n3504;
wire            n3505;
wire            n3506;
wire            n3507;
wire            n3508;
wire            n3509;
wire            n351;
wire            n3510;
wire            n3511;
wire            n3512;
wire            n3513;
wire            n3514;
wire            n3515;
wire            n3516;
wire            n3517;
wire            n3518;
wire            n3519;
wire            n352;
wire            n3520;
wire            n3521;
wire            n3522;
wire            n3523;
wire            n3524;
wire            n3525;
wire            n3526;
wire            n3527;
wire            n3528;
wire            n3529;
wire            n353;
wire            n3530;
wire            n3531;
wire            n3532;
wire            n3533;
wire            n3534;
wire            n3535;
wire            n3536;
wire            n3537;
wire            n3538;
wire            n3539;
wire            n354;
wire            n3540;
wire            n3541;
wire            n3542;
wire            n3543;
wire            n3544;
wire            n3545;
wire            n3546;
wire            n3547;
wire            n3548;
wire            n3549;
wire            n355;
wire            n3550;
wire            n3551;
wire            n3552;
wire            n3553;
wire            n3554;
wire            n3555;
wire            n3556;
wire            n3557;
wire            n3558;
wire            n3559;
wire            n356;
wire            n3560;
wire            n3561;
wire            n3562;
wire            n3563;
wire            n3564;
wire            n3565;
wire            n3566;
wire            n3567;
wire            n3568;
wire            n3569;
wire            n357;
wire            n3570;
wire            n3571;
wire            n3572;
wire            n3573;
wire            n3574;
wire            n3575;
wire            n3576;
wire            n3577;
wire            n3578;
wire            n3579;
wire            n358;
wire            n3580;
wire            n3581;
wire            n3582;
wire            n3583;
wire            n3584;
wire            n3585;
wire            n3586;
wire            n3587;
wire            n3588;
wire            n3589;
wire            n359;
wire            n3590;
wire            n3591;
wire            n3592;
wire            n3593;
wire            n3594;
wire            n3595;
wire            n3596;
wire            n3597;
wire            n3598;
wire            n3599;
wire            n36;
wire            n360;
wire            n3600;
wire            n3601;
wire            n3602;
wire            n3603;
wire            n3604;
wire            n3605;
wire            n3606;
wire            n3607;
wire            n3608;
wire            n3609;
wire            n361;
wire            n3610;
wire            n3611;
wire            n3612;
wire            n3613;
wire            n3614;
wire            n3615;
wire            n3616;
wire            n3617;
wire            n3618;
wire            n3619;
wire            n362;
wire            n3620;
wire            n3621;
wire            n3622;
wire            n3623;
wire            n3624;
wire            n3625;
wire            n3626;
wire            n3627;
wire            n3628;
wire            n3629;
wire            n363;
wire            n3630;
wire            n3631;
wire            n3632;
wire            n3633;
wire            n3634;
wire            n3635;
wire            n3636;
wire            n3637;
wire            n3638;
wire            n3639;
wire            n364;
wire            n3640;
wire            n3641;
wire            n3642;
wire            n3643;
wire            n3644;
wire            n3645;
wire            n3646;
wire            n3647;
wire            n3648;
wire            n3649;
wire            n365;
wire            n3650;
wire            n3651;
wire            n3652;
wire            n3653;
wire            n3654;
wire            n3655;
wire            n3656;
wire            n3657;
wire            n3658;
wire            n3659;
wire            n366;
wire            n3660;
wire            n3661;
wire            n3662;
wire            n3663;
wire            n3664;
wire            n3665;
wire            n3666;
wire            n3667;
wire            n3668;
wire            n3669;
wire            n367;
wire            n3670;
wire            n3671;
wire            n3672;
wire            n3673;
wire            n3674;
wire            n3675;
wire            n3676;
wire            n3677;
wire            n3678;
wire            n3679;
wire            n368;
wire            n3680;
wire            n3681;
wire            n3682;
wire            n3683;
wire            n3684;
wire            n3685;
wire            n3686;
wire            n3687;
wire            n3688;
wire            n3689;
wire            n369;
wire            n3690;
wire            n3691;
wire            n3692;
wire            n3693;
wire            n3694;
wire            n3695;
wire            n3696;
wire            n3697;
wire            n3698;
wire            n3699;
wire            n37;
wire            n370;
wire            n3700;
wire            n3701;
wire            n3702;
wire            n3703;
wire            n3704;
wire            n3705;
wire            n3706;
wire            n3707;
wire            n3708;
wire            n3709;
wire            n371;
wire            n3710;
wire            n3711;
wire            n3712;
wire            n3713;
wire            n3714;
wire            n3715;
wire            n3716;
wire            n3717;
wire            n3718;
wire            n3719;
wire            n372;
wire            n3720;
wire            n3721;
wire            n3722;
wire            n3723;
wire            n3724;
wire            n3725;
wire            n3726;
wire            n3727;
wire            n3728;
wire            n3729;
wire            n373;
wire            n3730;
wire            n3731;
wire            n3732;
wire            n3733;
wire            n3734;
wire            n3735;
wire            n3736;
wire            n3737;
wire            n3738;
wire            n3739;
wire            n374;
wire            n3740;
wire            n3741;
wire            n3742;
wire            n3743;
wire            n3744;
wire            n3745;
wire            n3746;
wire            n3747;
wire            n3748;
wire            n3749;
wire            n375;
wire            n3750;
wire            n3751;
wire            n3752;
wire            n3753;
wire            n3754;
wire            n3755;
wire            n3756;
wire            n3757;
wire            n3758;
wire            n3759;
wire            n376;
wire            n3760;
wire            n3761;
wire            n3762;
wire            n3763;
wire            n3764;
wire            n3765;
wire            n3766;
wire            n3767;
wire            n3768;
wire            n3769;
wire            n377;
wire            n3770;
wire            n3771;
wire            n3772;
wire            n3773;
wire            n3774;
wire            n3775;
wire            n3776;
wire            n3777;
wire            n3778;
wire            n3779;
wire            n378;
wire            n3780;
wire            n3781;
wire            n3782;
wire            n3783;
wire            n3784;
wire            n3785;
wire            n3786;
wire            n3787;
wire            n3788;
wire            n3789;
wire            n379;
wire            n3790;
wire            n3791;
wire            n3792;
wire            n3793;
wire            n3794;
wire            n3795;
wire            n3796;
wire            n3797;
wire            n3798;
wire            n3799;
wire            n38;
wire            n380;
wire            n3800;
wire            n3801;
wire            n3802;
wire            n3803;
wire            n3804;
wire            n3805;
wire            n3806;
wire            n3807;
wire            n3808;
wire            n3809;
wire            n381;
wire            n3810;
wire            n3811;
wire            n3812;
wire            n3813;
wire            n3814;
wire            n3815;
wire            n3816;
wire            n3817;
wire            n3818;
wire            n3819;
wire            n382;
wire            n3820;
wire            n3821;
wire            n3822;
wire            n3823;
wire            n3824;
wire            n3825;
wire            n3826;
wire            n3827;
wire            n3828;
wire            n3829;
wire            n383;
wire            n3830;
wire            n3831;
wire            n3832;
wire            n3833;
wire            n3834;
wire            n3835;
wire            n3836;
wire            n3837;
wire            n3838;
wire            n3839;
wire            n384;
wire            n3840;
wire            n3841;
wire            n3842;
wire            n3843;
wire            n3844;
wire            n3845;
wire            n3846;
wire            n3847;
wire            n3848;
wire            n3849;
wire            n385;
wire            n3850;
wire            n3851;
wire            n3852;
wire            n3853;
wire            n3854;
wire            n3855;
wire            n3856;
wire            n3857;
wire            n3858;
wire            n3859;
wire            n386;
wire            n3860;
wire            n3861;
wire            n3862;
wire            n3863;
wire            n3864;
wire            n3865;
wire            n3866;
wire            n3867;
wire            n3868;
wire            n3869;
wire            n387;
wire            n3870;
wire            n3871;
wire            n3872;
wire            n3873;
wire            n3874;
wire            n3875;
wire            n3876;
wire            n3877;
wire            n3878;
wire            n3879;
wire            n388;
wire            n3880;
wire            n3881;
wire            n3882;
wire            n3883;
wire            n3884;
wire            n3885;
wire            n3886;
wire            n3887;
wire            n3888;
wire            n3889;
wire            n389;
wire            n3890;
wire            n3891;
wire            n3892;
wire            n3893;
wire            n3894;
wire            n3895;
wire            n3896;
wire            n3897;
wire            n3898;
wire            n3899;
wire            n39;
wire            n390;
wire            n3900;
wire            n3901;
wire            n3902;
wire            n3903;
wire            n3904;
wire            n3905;
wire            n3906;
wire            n3907;
wire            n3908;
wire            n3909;
wire            n391;
wire            n3910;
wire            n3911;
wire            n3912;
wire            n3913;
wire            n3914;
wire            n3915;
wire            n3916;
wire            n3917;
wire            n3918;
wire            n3919;
wire            n392;
wire            n3920;
wire            n3921;
wire            n3922;
wire            n3923;
wire            n3924;
wire            n3925;
wire            n3926;
wire            n3927;
wire            n3928;
wire            n3929;
wire            n393;
wire            n3930;
wire            n3931;
wire            n3932;
wire            n3933;
wire            n3934;
wire            n3935;
wire            n3936;
wire            n3937;
wire            n3938;
wire            n3939;
wire            n394;
wire            n3940;
wire            n3941;
wire            n3942;
wire            n3943;
wire            n3944;
wire            n3945;
wire            n3946;
wire            n3947;
wire            n3948;
wire            n3949;
wire            n395;
wire            n3950;
wire            n3951;
wire            n3952;
wire            n3953;
wire            n3954;
wire            n3955;
wire            n3956;
wire            n3957;
wire            n3958;
wire            n3959;
wire            n396;
wire            n3960;
wire            n3961;
wire            n3962;
wire            n3963;
wire            n3964;
wire            n3965;
wire            n3966;
wire            n3967;
wire            n3968;
wire            n3969;
wire            n397;
wire            n3970;
wire            n3971;
wire            n3972;
wire            n3973;
wire            n3974;
wire            n3975;
wire            n3976;
wire            n3977;
wire            n3978;
wire            n3979;
wire            n398;
wire            n3980;
wire            n3981;
wire            n3982;
wire            n3983;
wire            n3984;
wire            n3985;
wire            n3986;
wire            n3987;
wire            n3988;
wire            n3989;
wire            n399;
wire            n3990;
wire            n3991;
wire            n3992;
wire            n3993;
wire            n3994;
wire            n3995;
wire            n3996;
wire            n3997;
wire            n3998;
wire            n3999;
wire            n4;
wire            n40;
wire            n400;
wire            n4000;
wire            n4001;
wire            n4002;
wire            n4003;
wire            n4004;
wire            n4005;
wire            n4006;
wire            n4007;
wire            n4008;
wire            n4009;
wire            n401;
wire            n4010;
wire            n4011;
wire            n4012;
wire            n4013;
wire            n4014;
wire            n4015;
wire            n4016;
wire            n4017;
wire            n4018;
wire            n4019;
wire            n402;
wire            n4020;
wire            n4021;
wire            n4022;
wire            n4023;
wire            n4024;
wire            n4025;
wire            n4026;
wire            n4027;
wire            n4028;
wire            n4029;
wire            n403;
wire            n4030;
wire            n4031;
wire            n4032;
wire            n4033;
wire            n4034;
wire            n4035;
wire            n4036;
wire            n4037;
wire            n4038;
wire            n4039;
wire            n404;
wire            n4040;
wire            n4041;
wire            n4042;
wire            n4043;
wire            n4044;
wire            n4045;
wire            n4046;
wire            n4047;
wire            n4048;
wire            n4049;
wire            n405;
wire            n4050;
wire            n4051;
wire            n4052;
wire            n4053;
wire            n4054;
wire            n4055;
wire            n4056;
wire            n4057;
wire            n4058;
wire            n4059;
wire            n406;
wire            n4060;
wire            n4061;
wire            n4062;
wire            n4063;
wire            n4064;
wire            n4065;
wire            n4066;
wire            n4067;
wire            n4068;
wire            n4069;
wire            n407;
wire            n4070;
wire            n4071;
wire            n4072;
wire            n4073;
wire            n4074;
wire            n4075;
wire            n4076;
wire            n4077;
wire            n4078;
wire            n4079;
wire            n408;
wire            n4080;
wire            n4081;
wire            n4082;
wire            n4083;
wire            n4084;
wire            n4085;
wire            n4086;
wire            n4087;
wire            n4088;
wire            n4089;
wire            n409;
wire            n4090;
wire            n4091;
wire            n4092;
wire            n4093;
wire            n4094;
wire            n4095;
wire            n4096;
wire            n4097;
wire            n4098;
wire            n4099;
wire            n41;
wire            n410;
wire            n4100;
wire            n4101;
wire            n4102;
wire            n4103;
wire            n4104;
wire            n4105;
wire            n4106;
wire            n4107;
wire            n4108;
wire            n4109;
wire            n411;
wire            n4110;
wire            n4111;
wire            n4112;
wire            n4113;
wire            n4114;
wire            n4115;
wire            n4116;
wire            n4117;
wire            n4118;
wire            n4119;
wire            n412;
wire            n4120;
wire            n4121;
wire            n4122;
wire            n4123;
wire            n4124;
wire            n4125;
wire            n4126;
wire            n4127;
wire            n4128;
wire            n4129;
wire            n413;
wire            n4130;
wire            n4131;
wire            n4132;
wire            n4133;
wire            n4134;
wire            n4135;
wire            n4136;
wire            n4137;
wire            n4138;
wire            n4139;
wire            n414;
wire            n4140;
wire            n4141;
wire            n4142;
wire            n4143;
wire            n4144;
wire            n4145;
wire            n4146;
wire            n4147;
wire            n4148;
wire            n4149;
wire            n415;
wire            n4150;
wire            n4151;
wire            n4152;
wire            n4153;
wire            n4154;
wire            n4155;
wire            n4156;
wire            n4157;
wire            n4158;
wire            n4159;
wire            n416;
wire            n4160;
wire            n4161;
wire            n4162;
wire            n4163;
wire            n4164;
wire            n4165;
wire            n4166;
wire            n4167;
wire            n4168;
wire            n4169;
wire            n417;
wire            n4170;
wire            n4171;
wire            n4172;
wire            n4173;
wire            n4174;
wire            n4175;
wire            n4176;
wire            n4177;
wire            n4178;
wire            n4179;
wire            n418;
wire            n4180;
wire            n4181;
wire            n4182;
wire            n4183;
wire            n4184;
wire            n4185;
wire            n4186;
wire            n4187;
wire            n4188;
wire            n4189;
wire            n419;
wire            n4190;
wire            n4191;
wire            n4192;
wire            n4193;
wire            n4194;
wire            n4195;
wire            n4196;
wire            n4197;
wire            n4198;
wire            n4199;
wire            n42;
wire            n420;
wire            n4200;
wire            n4201;
wire            n4202;
wire            n4203;
wire            n4204;
wire            n4205;
wire            n4206;
wire            n4207;
wire            n4208;
wire            n4209;
wire            n421;
wire            n4210;
wire            n4211;
wire            n4212;
wire            n4213;
wire            n4214;
wire            n4215;
wire            n4216;
wire            n4217;
wire            n4218;
wire            n4219;
wire            n422;
wire            n4220;
wire            n4221;
wire            n4222;
wire            n4223;
wire            n4224;
wire            n4225;
wire            n4226;
wire            n4227;
wire            n4228;
wire            n4229;
wire            n423;
wire            n4230;
wire            n4231;
wire            n4232;
wire            n4233;
wire            n4234;
wire            n4235;
wire            n4236;
wire            n4237;
wire            n4238;
wire            n4239;
wire            n424;
wire            n4240;
wire            n4241;
wire            n4242;
wire            n4243;
wire            n4244;
wire            n4245;
wire            n4246;
wire            n4247;
wire            n4248;
wire            n4249;
wire            n425;
wire            n4250;
wire            n4251;
wire            n4252;
wire            n4253;
wire            n4254;
wire            n4255;
wire            n4256;
wire            n4257;
wire            n4258;
wire            n4259;
wire            n426;
wire            n4260;
wire            n4261;
wire            n4262;
wire            n4263;
wire            n4264;
wire            n4265;
wire            n4266;
wire            n4267;
wire            n4268;
wire            n4269;
wire            n427;
wire            n4270;
wire            n4271;
wire            n4272;
wire            n4273;
wire            n4274;
wire            n4275;
wire            n4276;
wire            n4277;
wire            n4278;
wire            n4279;
wire            n428;
wire            n4280;
wire            n4281;
wire            n4282;
wire            n4283;
wire            n4284;
wire            n4285;
wire            n4286;
wire            n4287;
wire            n4288;
wire            n4289;
wire            n429;
wire            n4290;
wire            n4291;
wire            n4292;
wire            n4293;
wire            n4294;
wire            n4295;
wire            n4296;
wire            n4297;
wire            n4298;
wire            n4299;
wire            n43;
wire            n430;
wire            n4300;
wire            n4301;
wire            n4302;
wire            n4303;
wire            n4304;
wire            n4305;
wire            n4306;
wire            n4307;
wire            n4308;
wire            n4309;
wire            n431;
wire            n4310;
wire            n4311;
wire            n4312;
wire            n4313;
wire            n4314;
wire            n4315;
wire            n4316;
wire            n4317;
wire            n4318;
wire            n4319;
wire            n432;
wire            n4320;
wire            n4321;
wire            n4322;
wire            n4323;
wire            n4324;
wire            n4325;
wire            n4326;
wire            n4327;
wire            n4328;
wire            n4329;
wire            n433;
wire            n4330;
wire            n4331;
wire            n4332;
wire            n4333;
wire            n4334;
wire            n4335;
wire            n4336;
wire            n4337;
wire            n4338;
wire            n4339;
wire            n434;
wire            n4340;
wire            n4341;
wire            n4342;
wire            n4343;
wire            n4344;
wire            n4345;
wire            n4346;
wire            n4347;
wire            n4348;
wire            n4349;
wire            n435;
wire            n4350;
wire            n4351;
wire            n4352;
wire            n4353;
wire            n4354;
wire            n4355;
wire            n4356;
wire            n4357;
wire            n4358;
wire            n4359;
wire            n436;
wire            n4360;
wire            n4361;
wire            n4362;
wire            n4363;
wire            n4364;
wire            n4365;
wire            n4366;
wire            n4367;
wire            n4368;
wire            n4369;
wire            n437;
wire            n4370;
wire            n4371;
wire            n4372;
wire            n4373;
wire            n4374;
wire            n4375;
wire            n4376;
wire            n4377;
wire            n4378;
wire            n4379;
wire            n438;
wire            n4380;
wire            n4381;
wire            n4382;
wire            n4383;
wire            n4384;
wire            n4385;
wire            n4386;
wire            n4387;
wire            n4388;
wire            n4389;
wire            n439;
wire            n4390;
wire            n4391;
wire            n4392;
wire            n4393;
wire            n4394;
wire            n4395;
wire            n4396;
wire            n4397;
wire            n4398;
wire            n4399;
wire            n44;
wire            n440;
wire            n4400;
wire            n4401;
wire            n4402;
wire            n4403;
wire            n4404;
wire            n4405;
wire            n4406;
wire            n4407;
wire            n4408;
wire            n4409;
wire            n441;
wire            n4410;
wire            n4411;
wire            n4412;
wire            n4413;
wire            n4414;
wire            n4415;
wire            n4416;
wire            n4417;
wire            n4418;
wire            n4419;
wire            n442;
wire            n4420;
wire            n4421;
wire            n4422;
wire            n4423;
wire            n4424;
wire            n4425;
wire            n4426;
wire            n4427;
wire            n4428;
wire            n4429;
wire            n443;
wire            n4430;
wire            n4431;
wire            n4432;
wire            n4433;
wire            n4434;
wire            n4435;
wire            n4436;
wire            n4437;
wire            n4438;
wire            n4439;
wire            n444;
wire            n4440;
wire            n4441;
wire            n4442;
wire            n4443;
wire            n4444;
wire            n4445;
wire            n4446;
wire            n4447;
wire            n4448;
wire            n4449;
wire            n445;
wire            n4450;
wire            n4451;
wire            n4452;
wire            n4453;
wire            n4454;
wire            n4455;
wire            n4456;
wire            n4457;
wire            n4458;
wire            n4459;
wire            n446;
wire            n4460;
wire            n4461;
wire            n4462;
wire            n4463;
wire            n4464;
wire            n4465;
wire            n4466;
wire            n4467;
wire            n4468;
wire            n4469;
wire            n447;
wire            n4470;
wire            n4471;
wire            n4472;
wire            n4473;
wire            n4474;
wire            n4475;
wire            n4476;
wire            n4477;
wire            n4478;
wire            n4479;
wire            n448;
wire            n4480;
wire            n4481;
wire            n4482;
wire            n4483;
wire            n4484;
wire            n4485;
wire            n4486;
wire            n4487;
wire            n4488;
wire            n4489;
wire            n449;
wire            n4490;
wire            n4491;
wire            n4492;
wire            n4493;
wire            n4494;
wire            n4495;
wire            n4496;
wire            n4497;
wire            n4498;
wire            n4499;
wire            n45;
wire            n450;
wire            n4500;
wire            n4501;
wire            n4502;
wire            n4503;
wire            n4504;
wire            n4505;
wire            n4506;
wire            n4507;
wire            n4508;
wire            n4509;
wire            n451;
wire            n4510;
wire            n4511;
wire            n4512;
wire            n4513;
wire            n4514;
wire            n4515;
wire            n4516;
wire            n4517;
wire            n4518;
wire            n4519;
wire            n452;
wire            n4520;
wire            n4521;
wire            n4522;
wire            n4523;
wire            n4524;
wire            n4525;
wire            n4526;
wire            n4527;
wire            n4528;
wire            n4529;
wire            n453;
wire            n4530;
wire            n4531;
wire            n4532;
wire            n4533;
wire            n4534;
wire            n4535;
wire            n4536;
wire            n4537;
wire            n4538;
wire            n4539;
wire            n454;
wire            n4540;
wire            n4541;
wire            n4542;
wire            n4543;
wire            n4544;
wire            n4545;
wire            n4546;
wire            n4547;
wire            n4548;
wire            n4549;
wire            n455;
wire            n4550;
wire            n4551;
wire            n4552;
wire            n4553;
wire            n4554;
wire            n4555;
wire            n4556;
wire            n4557;
wire            n4558;
wire            n4559;
wire            n456;
wire            n4560;
wire            n4561;
wire            n4562;
wire            n4563;
wire            n4564;
wire            n4565;
wire            n4566;
wire            n4567;
wire            n4568;
wire            n4569;
wire            n457;
wire            n4570;
wire            n4571;
wire            n4572;
wire            n4573;
wire            n4574;
wire            n4575;
wire            n4576;
wire            n4577;
wire            n4578;
wire            n4579;
wire            n458;
wire            n4580;
wire            n4581;
wire            n4582;
wire            n4583;
wire            n4584;
wire            n4585;
wire            n4586;
wire            n4587;
wire            n4588;
wire            n4589;
wire            n459;
wire            n4590;
wire            n4591;
wire            n4592;
wire            n4593;
wire            n4594;
wire            n4595;
wire            n4596;
wire            n4597;
wire            n4598;
wire            n4599;
wire            n46;
wire            n460;
wire            n4600;
wire            n4601;
wire            n4602;
wire            n4603;
wire            n4604;
wire            n4605;
wire            n4606;
wire            n4607;
wire            n4608;
wire            n4609;
wire            n461;
wire            n4610;
wire            n4611;
wire            n4612;
wire            n4613;
wire            n4614;
wire            n4615;
wire            n4616;
wire            n4617;
wire            n4618;
wire            n4619;
wire            n462;
wire            n4620;
wire            n4621;
wire            n4622;
wire            n4623;
wire            n4624;
wire            n4625;
wire            n4626;
wire            n4627;
wire            n4628;
wire            n4629;
wire            n463;
wire            n4630;
wire            n4631;
wire            n4632;
wire            n4633;
wire            n4634;
wire            n4635;
wire            n4636;
wire            n4637;
wire            n4638;
wire            n4639;
wire            n464;
wire            n4640;
wire            n4641;
wire            n4642;
wire            n4643;
wire            n4644;
wire            n4645;
wire            n4646;
wire            n4647;
wire            n4648;
wire            n4649;
wire            n465;
wire            n4650;
wire            n4651;
wire            n4652;
wire            n4653;
wire            n4654;
wire            n4655;
wire            n4656;
wire            n4657;
wire            n4658;
wire            n4659;
wire            n466;
wire            n4660;
wire            n4661;
wire            n4662;
wire            n4663;
wire            n4664;
wire            n4665;
wire            n4666;
wire            n4667;
wire            n4668;
wire            n4669;
wire            n467;
wire            n4670;
wire            n4671;
wire            n4672;
wire            n4673;
wire            n4674;
wire            n4675;
wire            n4676;
wire            n4677;
wire            n4678;
wire            n4679;
wire            n468;
wire            n4680;
wire            n4681;
wire            n4682;
wire            n4683;
wire            n4684;
wire            n4685;
wire            n4686;
wire            n4687;
wire            n4688;
wire            n4689;
wire            n469;
wire            n4690;
wire            n4691;
wire            n4692;
wire            n4693;
wire            n4694;
wire            n4695;
wire            n4696;
wire            n4697;
wire            n4698;
wire            n4699;
wire            n47;
wire            n470;
wire            n4700;
wire            n4701;
wire            n4702;
wire            n4703;
wire            n4704;
wire            n4705;
wire            n4706;
wire            n4707;
wire            n4708;
wire            n4709;
wire            n471;
wire            n4710;
wire            n4711;
wire            n4712;
wire            n4713;
wire            n4714;
wire            n4715;
wire            n4716;
wire            n4717;
wire            n4718;
wire            n4719;
wire            n472;
wire            n4720;
wire            n4721;
wire            n4722;
wire            n4723;
wire            n4724;
wire            n4725;
wire            n4726;
wire            n4727;
wire            n4728;
wire            n4729;
wire            n473;
wire            n4730;
wire            n4731;
wire            n4732;
wire            n4733;
wire            n4734;
wire            n4735;
wire            n4736;
wire            n4737;
wire            n4738;
wire            n4739;
wire            n474;
wire            n4740;
wire            n4741;
wire            n4742;
wire            n4743;
wire            n4744;
wire            n4745;
wire            n4746;
wire            n4747;
wire            n4748;
wire            n4749;
wire            n475;
wire            n4750;
wire            n4751;
wire            n4752;
wire            n4753;
wire            n4754;
wire            n4755;
wire            n4756;
wire            n4757;
wire            n4758;
wire            n4759;
wire            n476;
wire            n4760;
wire            n4761;
wire            n4762;
wire            n4763;
wire            n4764;
wire            n4765;
wire            n4766;
wire            n4767;
wire            n4768;
wire            n4769;
wire            n477;
wire            n4770;
wire            n4771;
wire            n4772;
wire            n4773;
wire            n4774;
wire            n4775;
wire            n4776;
wire            n4777;
wire            n4778;
wire            n4779;
wire            n478;
wire            n4780;
wire            n4781;
wire            n4782;
wire            n4783;
wire            n4784;
wire            n4785;
wire            n4786;
wire            n4787;
wire            n4788;
wire            n4789;
wire            n479;
wire            n4790;
wire            n4791;
wire            n4792;
wire            n4793;
wire            n4794;
wire            n4795;
wire            n4796;
wire            n4797;
wire            n4798;
wire            n4799;
wire            n48;
wire            n480;
wire            n4800;
wire            n4801;
wire            n4802;
wire            n4803;
wire            n4804;
wire            n4805;
wire            n4806;
wire            n4807;
wire            n4808;
wire            n4809;
wire            n481;
wire            n4810;
wire            n4811;
wire            n4812;
wire            n4813;
wire            n4814;
wire            n4815;
wire            n4816;
wire            n4817;
wire            n4818;
wire            n4819;
wire            n482;
wire            n4820;
wire            n4821;
wire            n4822;
wire            n4823;
wire            n4824;
wire            n4825;
wire            n4826;
wire            n4827;
wire            n4828;
wire            n4829;
wire            n483;
wire            n4830;
wire            n4831;
wire            n4832;
wire            n4833;
wire            n4834;
wire            n4835;
wire            n4836;
wire            n4837;
wire            n4838;
wire            n4839;
wire            n484;
wire            n4840;
wire            n4841;
wire            n4842;
wire            n4843;
wire            n4844;
wire            n4845;
wire            n4846;
wire            n4847;
wire            n4848;
wire            n4849;
wire            n485;
wire            n4850;
wire            n4851;
wire            n4852;
wire            n4853;
wire            n4854;
wire            n4855;
wire            n4856;
wire            n4857;
wire            n4858;
wire            n4859;
wire            n486;
wire            n4860;
wire            n4861;
wire            n4862;
wire            n4863;
wire            n4864;
wire            n4865;
wire            n4866;
wire            n4867;
wire            n4868;
wire            n4869;
wire            n487;
wire            n4870;
wire            n4871;
wire            n4872;
wire            n4873;
wire            n4874;
wire            n4875;
wire            n4876;
wire            n4877;
wire            n4878;
wire            n4879;
wire            n488;
wire            n4880;
wire            n4881;
wire            n4882;
wire            n4883;
wire            n4884;
wire            n4885;
wire            n4886;
wire            n4887;
wire            n4888;
wire            n4889;
wire            n489;
wire            n4890;
wire            n4891;
wire            n4892;
wire            n4893;
wire            n4894;
wire            n4895;
wire            n4896;
wire            n4897;
wire            n4898;
wire            n4899;
wire            n49;
wire            n490;
wire            n4900;
wire            n4901;
wire            n4902;
wire            n4903;
wire            n4904;
wire            n4905;
wire            n4906;
wire            n4907;
wire            n4908;
wire            n4909;
wire            n491;
wire            n4910;
wire            n4911;
wire            n4912;
wire            n4913;
wire            n4914;
wire            n4915;
wire            n4916;
wire            n4917;
wire            n4918;
wire            n4919;
wire            n492;
wire            n4920;
wire            n4921;
wire            n4922;
wire            n4923;
wire            n4924;
wire            n4925;
wire            n4926;
wire            n4927;
wire            n4928;
wire            n4929;
wire            n493;
wire            n4930;
wire            n4931;
wire            n4932;
wire            n4933;
wire            n4934;
wire            n4935;
wire            n4936;
wire            n4937;
wire            n4938;
wire            n4939;
wire            n494;
wire            n4940;
wire            n4941;
wire            n4942;
wire            n4943;
wire            n4944;
wire            n4945;
wire            n4946;
wire            n4947;
wire            n4948;
wire            n4949;
wire            n495;
wire            n4950;
wire            n4951;
wire            n4952;
wire            n4953;
wire            n4954;
wire            n4955;
wire            n4956;
wire            n4957;
wire            n4958;
wire            n4959;
wire            n496;
wire            n4960;
wire            n4961;
wire            n4962;
wire            n4963;
wire            n4964;
wire            n4965;
wire            n4966;
wire            n4967;
wire            n4968;
wire            n4969;
wire            n497;
wire            n4970;
wire            n4971;
wire            n4972;
wire            n4973;
wire            n4974;
wire            n4975;
wire            n4976;
wire            n4977;
wire            n4978;
wire            n4979;
wire            n498;
wire            n4980;
wire            n4981;
wire            n4982;
wire            n4983;
wire            n4984;
wire            n4985;
wire            n4986;
wire            n4987;
wire            n4988;
wire            n4989;
wire            n499;
wire            n4990;
wire            n4991;
wire            n4992;
wire            n4993;
wire            n4994;
wire            n4995;
wire            n4996;
wire            n4997;
wire            n4998;
wire            n4999;
wire            n50;
wire            n500;
wire            n5000;
wire            n5001;
wire            n5002;
wire            n5003;
wire            n5004;
wire            n5005;
wire            n5006;
wire            n5007;
wire            n5008;
wire            n5009;
wire            n501;
wire            n5010;
wire            n5011;
wire            n5012;
wire            n5013;
wire            n5014;
wire            n5015;
wire            n5016;
wire            n5017;
wire            n5018;
wire            n5019;
wire            n502;
wire            n5020;
wire            n5021;
wire            n5022;
wire            n5023;
wire            n5024;
wire            n5025;
wire            n5026;
wire            n5027;
wire            n5028;
wire            n5029;
wire            n503;
wire            n5030;
wire            n5031;
wire            n5032;
wire            n5033;
wire            n5034;
wire            n5035;
wire            n5036;
wire            n5037;
wire            n5038;
wire            n5039;
wire            n504;
wire            n5040;
wire            n5041;
wire            n5042;
wire            n5043;
wire            n5044;
wire            n5045;
wire            n5046;
wire            n5047;
wire            n5048;
wire            n5049;
wire            n505;
wire            n5050;
wire            n5051;
wire            n5052;
wire            n5053;
wire            n5054;
wire            n5055;
wire            n5056;
wire            n5057;
wire            n5058;
wire            n5059;
wire            n506;
wire            n5060;
wire            n5061;
wire            n5062;
wire            n5063;
wire            n5064;
wire            n5065;
wire            n5066;
wire            n5067;
wire            n5068;
wire            n5069;
wire            n507;
wire            n5070;
wire            n5071;
wire            n5072;
wire            n5073;
wire            n5074;
wire            n5075;
wire            n5076;
wire            n5077;
wire            n5078;
wire            n5079;
wire            n508;
wire            n5080;
wire            n5081;
wire            n5082;
wire            n5083;
wire            n5084;
wire            n5085;
wire            n5086;
wire            n5087;
wire            n5088;
wire            n5089;
wire            n509;
wire            n5090;
wire            n5091;
wire            n5092;
wire            n5093;
wire            n5094;
wire            n5095;
wire            n5096;
wire            n5097;
wire            n5098;
wire            n5099;
wire            n51;
wire            n510;
wire            n5100;
wire            n5101;
wire            n5102;
wire            n5103;
wire            n5104;
wire            n5105;
wire            n5106;
wire            n5107;
wire            n5108;
wire            n5109;
wire            n511;
wire            n5110;
wire            n5111;
wire            n5112;
wire            n5113;
wire            n5114;
wire            n5115;
wire            n5116;
wire            n5117;
wire            n5118;
wire            n5119;
wire            n512;
wire            n5120;
wire            n5121;
wire            n5122;
wire            n5123;
wire            n5124;
wire            n5125;
wire            n5126;
wire            n5127;
wire            n5128;
wire            n5129;
wire            n513;
wire            n5130;
wire            n5131;
wire            n5132;
wire            n5133;
wire            n5134;
wire            n5135;
wire            n5136;
wire            n5137;
wire            n5138;
wire            n5139;
wire            n514;
wire            n5140;
wire            n5141;
wire            n5142;
wire            n5143;
wire            n5144;
wire            n5145;
wire            n5146;
wire            n5147;
wire            n5148;
wire            n5149;
wire            n515;
wire            n5150;
wire            n5151;
wire            n5152;
wire            n5153;
wire            n5154;
wire            n5155;
wire            n5156;
wire            n5157;
wire            n5158;
wire            n5159;
wire            n516;
wire            n5160;
wire            n5161;
wire            n5162;
wire            n5163;
wire            n5164;
wire            n5165;
wire            n5166;
wire            n5167;
wire            n5168;
wire            n5169;
wire            n517;
wire            n5170;
wire            n5171;
wire            n5172;
wire            n5173;
wire            n5174;
wire            n5175;
wire            n5176;
wire            n5177;
wire            n5178;
wire            n5179;
wire            n518;
wire            n5180;
wire            n5181;
wire            n5182;
wire            n5183;
wire            n5184;
wire            n5185;
wire            n5186;
wire            n5187;
wire            n5188;
wire            n5189;
wire            n519;
wire            n5190;
wire            n5191;
wire            n5192;
wire            n5193;
wire            n5194;
wire            n5195;
wire            n5196;
wire            n5197;
wire            n5198;
wire            n5199;
wire            n52;
wire            n520;
wire            n5200;
wire            n5201;
wire            n5202;
wire            n5203;
wire            n5204;
wire            n5205;
wire            n5206;
wire            n5207;
wire            n5208;
wire            n5209;
wire            n521;
wire            n5210;
wire            n5211;
wire            n5212;
wire            n5213;
wire            n5214;
wire            n5215;
wire            n5216;
wire            n5217;
wire            n5218;
wire            n5219;
wire            n522;
wire            n5220;
wire            n5221;
wire            n5222;
wire            n5223;
wire            n5224;
wire            n5225;
wire            n5226;
wire            n5227;
wire            n5228;
wire            n5229;
wire            n523;
wire            n5230;
wire            n5231;
wire            n5232;
wire            n5233;
wire            n5234;
wire            n5235;
wire            n5236;
wire            n5237;
wire            n5238;
wire            n5239;
wire            n524;
wire            n5240;
wire            n5241;
wire            n5242;
wire            n5243;
wire            n5244;
wire            n5245;
wire            n5246;
wire            n5247;
wire            n5248;
wire            n5249;
wire            n525;
wire            n5250;
wire            n5251;
wire            n5252;
wire            n5253;
wire            n5254;
wire            n5255;
wire            n5256;
wire            n5257;
wire            n5258;
wire            n5259;
wire            n526;
wire            n5260;
wire            n5261;
wire            n5262;
wire            n5263;
wire            n5264;
wire            n5265;
wire            n5266;
wire            n5267;
wire            n5268;
wire            n5269;
wire            n527;
wire            n5270;
wire            n5271;
wire            n5272;
wire            n5273;
wire            n5274;
wire            n5275;
wire            n5276;
wire            n5277;
wire            n5278;
wire            n5279;
wire            n528;
wire            n5280;
wire            n5281;
wire            n5282;
wire            n5283;
wire            n5284;
wire            n5285;
wire            n5286;
wire            n5287;
wire            n5288;
wire            n5289;
wire            n529;
wire            n5290;
wire            n5291;
wire            n5292;
wire            n5293;
wire            n5294;
wire            n5295;
wire            n5296;
wire            n5297;
wire            n5298;
wire            n5299;
wire            n53;
wire            n530;
wire            n5300;
wire            n5301;
wire            n5302;
wire            n5303;
wire            n5304;
wire            n5305;
wire            n5306;
wire            n5307;
wire            n5308;
wire            n5309;
wire            n531;
wire            n5310;
wire            n5311;
wire            n5312;
wire            n5313;
wire            n5314;
wire            n5315;
wire            n5316;
wire            n5317;
wire            n5318;
wire            n5319;
wire            n532;
wire            n5320;
wire            n5321;
wire            n5322;
wire            n5323;
wire            n5324;
wire            n5325;
wire            n5326;
wire            n5327;
wire            n5328;
wire            n5329;
wire            n533;
wire            n5330;
wire            n5331;
wire            n5332;
wire            n5333;
wire            n5334;
wire            n5335;
wire            n5336;
wire            n5337;
wire            n5338;
wire            n5339;
wire            n534;
wire            n5340;
wire            n5341;
wire            n5342;
wire            n5343;
wire            n5344;
wire            n5345;
wire            n5346;
wire            n5347;
wire            n5348;
wire            n5349;
wire            n535;
wire            n5350;
wire            n5351;
wire            n5352;
wire            n5353;
wire            n5354;
wire            n5355;
wire            n5356;
wire            n5357;
wire            n5358;
wire            n5359;
wire            n536;
wire            n5360;
wire            n5361;
wire            n5362;
wire            n5363;
wire            n5364;
wire            n5365;
wire            n5366;
wire            n5367;
wire            n5368;
wire            n5369;
wire            n537;
wire            n5370;
wire            n5371;
wire            n5372;
wire            n5373;
wire            n5374;
wire            n5375;
wire            n5376;
wire            n5377;
wire            n5378;
wire            n5379;
wire            n538;
wire            n5380;
wire            n5381;
wire            n5382;
wire            n5383;
wire            n5384;
wire            n5385;
wire            n5386;
wire            n5387;
wire            n5388;
wire            n5389;
wire            n539;
wire            n5390;
wire            n5391;
wire            n5392;
wire            n5393;
wire            n5394;
wire            n5395;
wire            n5396;
wire            n5397;
wire            n5398;
wire            n5399;
wire            n54;
wire            n540;
wire            n5400;
wire            n5401;
wire            n5402;
wire            n5403;
wire            n5404;
wire            n5405;
wire            n5406;
wire            n5407;
wire            n5408;
wire            n5409;
wire            n541;
wire            n5410;
wire            n5411;
wire            n5412;
wire            n5413;
wire            n5414;
wire            n5415;
wire            n5416;
wire            n5417;
wire            n5418;
wire            n5419;
wire            n542;
wire            n5420;
wire            n5421;
wire            n5422;
wire            n5423;
wire            n5424;
wire            n5425;
wire            n5426;
wire            n5427;
wire            n5428;
wire            n5429;
wire            n543;
wire            n5430;
wire            n5431;
wire            n5432;
wire            n5433;
wire            n5434;
wire            n5435;
wire            n5436;
wire            n5437;
wire            n5438;
wire            n5439;
wire            n544;
wire            n5440;
wire            n5441;
wire            n5442;
wire            n5443;
wire            n5444;
wire            n5445;
wire            n5446;
wire            n5447;
wire            n5448;
wire            n5449;
wire            n545;
wire            n5450;
wire            n5451;
wire            n5452;
wire            n5453;
wire            n5454;
wire            n5455;
wire            n5456;
wire            n5457;
wire            n5458;
wire            n5459;
wire            n546;
wire            n5460;
wire            n5461;
wire            n5462;
wire            n5463;
wire            n5464;
wire            n5465;
wire            n5466;
wire            n5467;
wire            n5468;
wire            n5469;
wire            n547;
wire            n5470;
wire            n5471;
wire            n5472;
wire            n5473;
wire            n5474;
wire            n5475;
wire            n5476;
wire            n5477;
wire            n5478;
wire            n5479;
wire            n548;
wire            n5480;
wire            n5481;
wire            n5482;
wire            n5483;
wire            n5484;
wire            n5485;
wire            n5486;
wire            n5487;
wire            n5488;
wire            n5489;
wire            n549;
wire            n5490;
wire            n5491;
wire            n5492;
wire            n5493;
wire            n5494;
wire            n5495;
wire            n5496;
wire            n5497;
wire            n5498;
wire            n5499;
wire            n55;
wire            n550;
wire            n5500;
wire            n5501;
wire            n5502;
wire            n5503;
wire            n5504;
wire            n5505;
wire            n5506;
wire            n5507;
wire            n5508;
wire            n5509;
wire            n551;
wire            n5510;
wire            n5511;
wire            n5512;
wire            n5513;
wire            n5514;
wire            n5515;
wire            n5516;
wire            n5517;
wire            n5518;
wire            n5519;
wire            n552;
wire            n5520;
wire            n5521;
wire            n5522;
wire            n5523;
wire            n5524;
wire            n5525;
wire            n5526;
wire            n5527;
wire            n5528;
wire            n5529;
wire            n553;
wire            n5530;
wire            n5531;
wire            n5532;
wire            n5533;
wire            n5534;
wire            n5535;
wire            n5536;
wire            n5537;
wire            n5538;
wire            n5539;
wire            n554;
wire            n5540;
wire            n5541;
wire            n5542;
wire            n5543;
wire            n5544;
wire            n5545;
wire            n5546;
wire            n5547;
wire            n5548;
wire            n5549;
wire            n555;
wire            n5550;
wire            n5551;
wire            n5552;
wire            n5553;
wire            n5554;
wire            n5555;
wire            n5556;
wire            n5557;
wire            n5558;
wire            n5559;
wire            n556;
wire            n5560;
wire            n5561;
wire            n5562;
wire            n5563;
wire            n5564;
wire            n5565;
wire            n5566;
wire            n5567;
wire            n5568;
wire            n5569;
wire            n557;
wire            n5570;
wire            n5571;
wire            n5572;
wire            n5573;
wire            n5574;
wire            n5575;
wire            n5576;
wire            n5577;
wire            n5578;
wire            n5579;
wire            n558;
wire            n5580;
wire            n5581;
wire            n5582;
wire            n5583;
wire            n5584;
wire            n5585;
wire            n5586;
wire            n5587;
wire            n5588;
wire            n5589;
wire            n559;
wire            n5590;
wire            n5591;
wire            n5592;
wire            n5593;
wire            n5594;
wire            n5595;
wire            n5596;
wire            n5597;
wire            n5598;
wire            n5599;
wire            n56;
wire            n560;
wire            n5600;
wire            n5601;
wire            n5602;
wire            n5603;
wire            n5604;
wire            n5605;
wire            n5606;
wire            n5607;
wire            n5608;
wire            n5609;
wire            n561;
wire            n5610;
wire            n5611;
wire            n5612;
wire            n5613;
wire            n5614;
wire            n5615;
wire            n5616;
wire            n5617;
wire            n5618;
wire            n5619;
wire            n562;
wire            n5620;
wire            n5621;
wire            n5622;
wire            n5623;
wire            n5624;
wire            n5625;
wire            n5626;
wire            n5627;
wire            n5628;
wire            n5629;
wire            n563;
wire            n5630;
wire            n5631;
wire            n5632;
wire            n5633;
wire            n5634;
wire            n5635;
wire            n5636;
wire            n5637;
wire            n5638;
wire            n5639;
wire            n564;
wire            n5640;
wire            n5641;
wire            n5642;
wire            n5643;
wire            n5644;
wire            n5645;
wire            n5646;
wire            n5647;
wire            n5648;
wire            n5649;
wire            n565;
wire            n5650;
wire            n5651;
wire            n5652;
wire            n5653;
wire            n5654;
wire            n5655;
wire            n5656;
wire            n5657;
wire            n5658;
wire            n5659;
wire            n566;
wire            n5660;
wire            n5661;
wire            n5662;
wire            n5663;
wire            n5664;
wire            n5665;
wire            n5666;
wire            n5667;
wire            n5668;
wire            n5669;
wire            n567;
wire            n5670;
wire            n5671;
wire            n5672;
wire            n5673;
wire            n5674;
wire            n5675;
wire            n5676;
wire            n5677;
wire            n5678;
wire            n5679;
wire            n568;
wire            n5680;
wire            n5681;
wire            n5682;
wire            n5683;
wire            n5684;
wire            n5685;
wire            n5686;
wire            n5687;
wire            n5688;
wire            n5689;
wire            n569;
wire            n5690;
wire            n5691;
wire            n5692;
wire            n5693;
wire            n5694;
wire            n5695;
wire            n5696;
wire            n5697;
wire            n5698;
wire            n5699;
wire            n57;
wire            n570;
wire            n5700;
wire            n5701;
wire            n5702;
wire            n5703;
wire            n5704;
wire            n5705;
wire            n5706;
wire            n5707;
wire            n5708;
wire            n5709;
wire            n571;
wire            n5710;
wire            n5711;
wire            n5712;
wire            n5713;
wire            n5714;
wire            n5715;
wire            n5716;
wire            n5717;
wire            n5718;
wire            n5719;
wire            n572;
wire            n5720;
wire            n5721;
wire            n5722;
wire            n5723;
wire            n5724;
wire            n5725;
wire            n5726;
wire            n5727;
wire            n5728;
wire            n5729;
wire            n573;
wire            n5730;
wire            n5731;
wire            n5732;
wire            n5733;
wire            n5734;
wire            n5735;
wire            n5736;
wire            n5737;
wire            n5738;
wire            n5739;
wire            n574;
wire            n5740;
wire            n5741;
wire            n5742;
wire            n5743;
wire            n5744;
wire            n5745;
wire            n5746;
wire            n5747;
wire            n5748;
wire            n5749;
wire            n575;
wire            n5750;
wire            n5751;
wire            n5752;
wire            n5753;
wire            n5754;
wire            n5755;
wire            n5756;
wire            n5757;
wire            n5758;
wire            n5759;
wire            n576;
wire            n5760;
wire            n5761;
wire            n5762;
wire            n5763;
wire            n5764;
wire            n5765;
wire            n5766;
wire            n5767;
wire            n5768;
wire            n5769;
wire            n577;
wire            n5770;
wire            n5771;
wire            n5772;
wire            n5773;
wire            n5774;
wire            n5775;
wire            n5776;
wire            n5777;
wire            n5778;
wire            n5779;
wire            n578;
wire            n5780;
wire            n5781;
wire            n5782;
wire            n5783;
wire            n5784;
wire            n5785;
wire            n5786;
wire            n5787;
wire            n5788;
wire            n5789;
wire            n579;
wire            n5790;
wire            n5791;
wire            n5792;
wire            n5793;
wire            n5794;
wire            n5795;
wire            n5796;
wire            n5797;
wire            n5798;
wire            n5799;
wire            n58;
wire            n580;
wire            n5800;
wire            n5801;
wire            n5802;
wire            n5803;
wire            n5804;
wire            n5805;
wire            n5806;
wire            n5807;
wire            n5808;
wire            n5809;
wire            n581;
wire            n5810;
wire            n5811;
wire            n5812;
wire            n5813;
wire            n5814;
wire            n5815;
wire            n5816;
wire            n5817;
wire            n5818;
wire            n5819;
wire            n582;
wire            n5820;
wire            n5821;
wire            n5822;
wire            n5823;
wire            n5824;
wire            n5825;
wire            n5826;
wire            n5827;
wire            n5828;
wire            n5829;
wire            n583;
wire            n5830;
wire            n5831;
wire            n5832;
wire            n5833;
wire            n5834;
wire            n5835;
wire            n5836;
wire            n5837;
wire            n5838;
wire            n5839;
wire            n584;
wire            n5840;
wire            n5841;
wire            n5842;
wire            n5843;
wire            n5844;
wire            n5845;
wire            n5846;
wire            n5847;
wire            n5848;
wire            n5849;
wire            n585;
wire            n5850;
wire            n5851;
wire            n5852;
wire            n5853;
wire            n5854;
wire            n5855;
wire            n5856;
wire            n5857;
wire            n5858;
wire            n5859;
wire            n586;
wire            n5860;
wire            n5861;
wire            n5862;
wire            n5863;
wire            n5864;
wire            n5865;
wire            n5866;
wire            n5867;
wire            n5868;
wire            n5869;
wire            n587;
wire            n5870;
wire            n5871;
wire            n5872;
wire            n5873;
wire            n5874;
wire            n5875;
wire            n5876;
wire            n5877;
wire            n5878;
wire            n5879;
wire            n588;
wire            n5880;
wire            n5881;
wire            n5882;
wire            n5883;
wire            n5884;
wire            n5885;
wire            n5886;
wire            n5887;
wire            n5888;
wire            n5889;
wire            n589;
wire            n5890;
wire            n5891;
wire            n5892;
wire            n5893;
wire            n5894;
wire            n5895;
wire            n5896;
wire            n5897;
wire            n5898;
wire            n5899;
wire            n59;
wire            n590;
wire            n5900;
wire            n5901;
wire            n5902;
wire            n5903;
wire            n5904;
wire            n5905;
wire            n5906;
wire            n5907;
wire            n5908;
wire            n5909;
wire            n591;
wire            n5910;
wire            n5911;
wire            n5912;
wire            n5913;
wire            n5914;
wire            n5915;
wire            n5916;
wire            n5917;
wire            n5918;
wire            n5919;
wire            n592;
wire            n5920;
wire            n5921;
wire            n5922;
wire            n5923;
wire            n5924;
wire            n5925;
wire            n5926;
wire            n5927;
wire            n5928;
wire            n5929;
wire            n593;
wire            n5930;
wire            n5931;
wire            n5932;
wire            n5933;
wire            n5934;
wire            n5935;
wire            n5936;
wire            n5937;
wire            n5938;
wire            n5939;
wire            n594;
wire            n5940;
wire            n5941;
wire            n5942;
wire            n5943;
wire            n5944;
wire            n5945;
wire            n5946;
wire            n5947;
wire            n5948;
wire            n5949;
wire            n595;
wire            n5950;
wire            n5951;
wire            n5952;
wire            n5953;
wire            n5954;
wire            n5955;
wire            n5956;
wire            n5957;
wire            n5958;
wire            n5959;
wire            n596;
wire            n5960;
wire            n5961;
wire            n5962;
wire            n5963;
wire            n5964;
wire            n5965;
wire            n5966;
wire            n5967;
wire            n5968;
wire            n5969;
wire            n597;
wire            n5970;
wire            n5971;
wire            n5972;
wire            n5973;
wire            n5974;
wire            n5975;
wire            n5976;
wire            n5977;
wire            n5978;
wire            n5979;
wire            n598;
wire            n5980;
wire            n5981;
wire            n5982;
wire            n5983;
wire            n5984;
wire            n5985;
wire            n5986;
wire            n5987;
wire            n5988;
wire            n5989;
wire            n599;
wire            n5990;
wire            n5991;
wire            n5992;
wire            n5993;
wire            n5994;
wire            n5995;
wire            n5996;
wire            n5997;
wire            n5998;
wire            n5999;
wire            n6;
wire            n60;
wire            n600;
wire            n6000;
wire            n6001;
wire            n6002;
wire            n6003;
wire            n6004;
wire            n6005;
wire            n6006;
wire            n6007;
wire            n6008;
wire            n6009;
wire            n601;
wire            n6010;
wire            n6011;
wire            n6012;
wire            n6013;
wire            n6014;
wire            n6015;
wire            n6016;
wire            n6017;
wire            n6018;
wire            n6019;
wire            n602;
wire            n6020;
wire            n6021;
wire            n6022;
wire            n6023;
wire            n6024;
wire            n6025;
wire            n6026;
wire            n6027;
wire            n6028;
wire            n6029;
wire            n603;
wire            n6030;
wire            n6031;
wire            n6032;
wire            n6033;
wire            n6034;
wire            n6035;
wire            n6036;
wire            n6037;
wire            n6038;
wire            n6039;
wire            n604;
wire            n6040;
wire            n6041;
wire            n6042;
wire            n6043;
wire            n6044;
wire            n6045;
wire            n6046;
wire            n6047;
wire            n6048;
wire            n6049;
wire            n605;
wire            n6050;
wire            n6051;
wire            n6052;
wire            n6053;
wire            n6054;
wire            n6055;
wire            n6056;
wire            n6057;
wire            n6058;
wire            n6059;
wire            n606;
wire            n6060;
wire            n6061;
wire            n6062;
wire            n6063;
wire            n6064;
wire            n6065;
wire            n6066;
wire            n6067;
wire            n6068;
wire            n6069;
wire            n607;
wire            n6070;
wire            n6071;
wire            n6072;
wire            n6073;
wire            n6074;
wire            n6075;
wire            n6076;
wire            n6077;
wire            n6078;
wire            n6079;
wire            n608;
wire            n6080;
wire            n6081;
wire            n6082;
wire            n6083;
wire            n6084;
wire            n6085;
wire            n6086;
wire            n6087;
wire            n6088;
wire            n6089;
wire            n609;
wire            n6090;
wire            n6091;
wire            n6092;
wire            n6093;
wire            n6094;
wire            n6095;
wire            n6096;
wire            n6097;
wire            n6098;
wire            n6099;
wire            n61;
wire            n610;
wire            n6100;
wire            n6101;
wire            n6102;
wire            n6103;
wire            n6104;
wire            n6105;
wire            n6106;
wire            n6107;
wire            n6108;
wire            n6109;
wire            n611;
wire            n6110;
wire            n6111;
wire            n6112;
wire            n6113;
wire            n6114;
wire            n6115;
wire            n6116;
wire            n6117;
wire            n6118;
wire            n6119;
wire            n612;
wire            n6120;
wire            n6121;
wire            n6122;
wire            n6123;
wire            n6124;
wire            n6125;
wire            n6126;
wire            n6127;
wire            n6128;
wire            n6129;
wire            n613;
wire            n6130;
wire            n6131;
wire            n6132;
wire            n6133;
wire            n6134;
wire            n6135;
wire            n6136;
wire            n6137;
wire            n6138;
wire            n6139;
wire            n614;
wire            n6140;
wire            n6141;
wire            n6142;
wire            n6143;
wire            n6144;
wire            n6145;
wire            n6146;
wire            n6147;
wire            n6148;
wire            n6149;
wire            n615;
wire            n6150;
wire            n6151;
wire            n6152;
wire            n6153;
wire            n6154;
wire            n6155;
wire            n6156;
wire            n6157;
wire            n6158;
wire            n6159;
wire            n616;
wire            n6160;
wire            n6161;
wire            n6162;
wire            n6163;
wire            n6164;
wire            n6165;
wire            n6166;
wire            n6167;
wire            n6168;
wire            n6169;
wire            n617;
wire            n6170;
wire            n6171;
wire            n6172;
wire            n6173;
wire            n6174;
wire            n6175;
wire            n6176;
wire            n6177;
wire            n6178;
wire            n6179;
wire            n618;
wire            n6180;
wire            n6181;
wire            n6182;
wire            n6183;
wire            n6184;
wire            n6185;
wire            n6186;
wire            n6187;
wire            n6188;
wire            n6189;
wire            n619;
wire            n6190;
wire            n6191;
wire            n6192;
wire            n6193;
wire            n6194;
wire            n6195;
wire            n6196;
wire            n6197;
wire            n6198;
wire            n6199;
wire            n62;
wire            n620;
wire            n6200;
wire            n6201;
wire            n6202;
wire            n6203;
wire            n6204;
wire            n6205;
wire            n6206;
wire            n6207;
wire            n6208;
wire            n6209;
wire            n621;
wire            n6210;
wire            n6211;
wire            n6212;
wire            n6213;
wire            n6214;
wire            n6215;
wire            n6216;
wire            n6217;
wire            n6218;
wire            n6219;
wire            n622;
wire            n6220;
wire            n6221;
wire            n6222;
wire            n6223;
wire            n6224;
wire            n6225;
wire            n6226;
wire            n6227;
wire            n6228;
wire            n6229;
wire            n623;
wire            n6230;
wire            n6231;
wire            n6232;
wire            n6233;
wire            n6234;
wire            n6235;
wire            n6236;
wire            n6237;
wire            n6238;
wire            n6239;
wire            n624;
wire            n6240;
wire            n6241;
wire            n6242;
wire            n6243;
wire            n6244;
wire            n6245;
wire            n6246;
wire            n6247;
wire            n6248;
wire            n6249;
wire            n625;
wire            n6250;
wire            n6251;
wire            n6252;
wire            n6253;
wire            n6254;
wire            n6255;
wire            n6256;
wire            n6257;
wire            n6258;
wire            n6259;
wire            n626;
wire            n6260;
wire            n6261;
wire            n6262;
wire            n6263;
wire            n6264;
wire            n6265;
wire            n6266;
wire            n6267;
wire            n6268;
wire            n6269;
wire            n627;
wire            n6270;
wire            n6271;
wire            n6272;
wire            n6273;
wire            n6274;
wire            n6275;
wire            n6276;
wire            n6277;
wire            n6278;
wire            n6279;
wire            n628;
wire            n6280;
wire            n6281;
wire            n6282;
wire            n6283;
wire            n6284;
wire            n6285;
wire            n6286;
wire            n6287;
wire            n6288;
wire            n6289;
wire            n629;
wire            n6290;
wire            n6291;
wire            n6292;
wire            n6293;
wire            n6294;
wire            n6295;
wire            n6296;
wire            n6297;
wire            n6298;
wire            n6299;
wire            n63;
wire            n630;
wire            n6300;
wire            n6301;
wire            n6302;
wire            n6303;
wire            n6304;
wire            n6305;
wire            n6306;
wire            n6307;
wire            n6308;
wire            n6309;
wire            n631;
wire            n6310;
wire            n6311;
wire            n6312;
wire            n6313;
wire            n6314;
wire            n6315;
wire            n6316;
wire            n6317;
wire            n6318;
wire            n6319;
wire            n632;
wire            n6320;
wire            n6321;
wire            n6322;
wire            n6323;
wire            n6324;
wire            n6325;
wire            n6326;
wire            n6327;
wire            n6328;
wire            n6329;
wire            n633;
wire            n6330;
wire            n6331;
wire            n6332;
wire            n6333;
wire            n6334;
wire            n6335;
wire            n6336;
wire            n6337;
wire            n6338;
wire            n6339;
wire            n634;
wire            n6340;
wire            n6341;
wire            n6342;
wire            n6343;
wire            n6344;
wire            n6345;
wire            n6346;
wire            n6347;
wire            n6348;
wire            n6349;
wire            n635;
wire            n6350;
wire            n6351;
wire            n6352;
wire            n6353;
wire            n6354;
wire            n6355;
wire            n6356;
wire            n6357;
wire            n6358;
wire            n6359;
wire            n636;
wire            n6360;
wire            n6361;
wire            n6362;
wire            n6363;
wire            n6364;
wire            n6365;
wire            n6366;
wire            n6367;
wire            n6368;
wire            n6369;
wire            n637;
wire            n6370;
wire            n6371;
wire            n6372;
wire            n6373;
wire            n6374;
wire            n6375;
wire            n6376;
wire            n6377;
wire            n6378;
wire            n6379;
wire            n638;
wire            n6380;
wire            n6381;
wire            n6382;
wire            n6383;
wire            n6384;
wire            n6385;
wire            n6386;
wire            n6387;
wire            n6388;
wire            n6389;
wire            n639;
wire            n6390;
wire            n6391;
wire            n6392;
wire            n6393;
wire            n6394;
wire            n6395;
wire            n6396;
wire            n6397;
wire            n6398;
wire            n6399;
wire            n64;
wire            n640;
wire            n6400;
wire            n6401;
wire            n6402;
wire            n6403;
wire            n6404;
wire            n6405;
wire            n6406;
wire            n6407;
wire            n6408;
wire            n6409;
wire            n641;
wire            n6410;
wire            n6411;
wire            n6412;
wire            n6413;
wire            n6414;
wire            n6415;
wire            n6416;
wire            n6417;
wire            n6418;
wire            n6419;
wire            n642;
wire            n6420;
wire            n6421;
wire            n6422;
wire            n6423;
wire            n6424;
wire            n6425;
wire            n6426;
wire            n6427;
wire            n6428;
wire            n6429;
wire            n643;
wire            n6430;
wire            n6431;
wire            n6432;
wire            n6433;
wire            n6434;
wire            n6435;
wire            n6436;
wire            n6437;
wire            n6438;
wire            n6439;
wire            n644;
wire            n6440;
wire            n6441;
wire            n6442;
wire            n6443;
wire            n6444;
wire            n6445;
wire            n6446;
wire            n6447;
wire            n6448;
wire            n6449;
wire            n645;
wire            n6450;
wire            n6451;
wire            n6452;
wire            n6453;
wire            n6454;
wire            n6455;
wire            n6456;
wire            n6457;
wire            n6458;
wire            n6459;
wire            n646;
wire            n6460;
wire            n6461;
wire            n6462;
wire            n6463;
wire            n6464;
wire            n6465;
wire            n6466;
wire            n6467;
wire            n6468;
wire            n6469;
wire            n647;
wire            n6470;
wire            n6471;
wire            n6472;
wire            n6473;
wire            n6474;
wire            n6475;
wire            n6476;
wire            n6477;
wire            n6478;
wire            n6479;
wire            n648;
wire            n6480;
wire            n6481;
wire            n6482;
wire            n6483;
wire            n6484;
wire            n6485;
wire            n6486;
wire            n6487;
wire            n6488;
wire            n6489;
wire            n649;
wire            n6490;
wire            n6491;
wire            n6492;
wire            n6493;
wire            n6494;
wire            n6495;
wire            n6496;
wire            n6497;
wire            n6498;
wire            n6499;
wire            n65;
wire            n650;
wire            n6500;
wire            n6501;
wire            n6502;
wire            n6503;
wire            n6504;
wire            n6505;
wire            n6506;
wire            n6507;
wire            n6508;
wire            n6509;
wire            n651;
wire            n6510;
wire            n6511;
wire            n6512;
wire            n6513;
wire            n6514;
wire            n6515;
wire            n6516;
wire            n6517;
wire            n6518;
wire            n6519;
wire            n652;
wire            n6520;
wire            n6521;
wire            n6522;
wire            n6523;
wire            n6524;
wire            n6525;
wire            n6526;
wire            n6527;
wire            n6528;
wire            n6529;
wire            n653;
wire            n6530;
wire            n6531;
wire            n6532;
wire            n6533;
wire            n6534;
wire            n6535;
wire            n6536;
wire            n6537;
wire            n6538;
wire            n6539;
wire            n654;
wire            n6540;
wire            n6541;
wire            n6542;
wire            n6543;
wire            n6544;
wire            n6545;
wire            n6546;
wire            n6547;
wire            n6548;
wire            n6549;
wire            n655;
wire            n6550;
wire            n6551;
wire            n6552;
wire            n6553;
wire            n6554;
wire            n6555;
wire            n6556;
wire            n6557;
wire            n6558;
wire            n6559;
wire            n656;
wire            n6560;
wire            n6561;
wire            n6562;
wire            n6563;
wire            n6564;
wire            n6565;
wire            n6566;
wire            n6567;
wire            n6568;
wire            n6569;
wire            n657;
wire            n6570;
wire            n6571;
wire            n6572;
wire            n6573;
wire            n6574;
wire            n6575;
wire            n6576;
wire            n6577;
wire            n6578;
wire            n6579;
wire            n658;
wire            n6580;
wire            n6581;
wire            n6582;
wire            n6583;
wire            n6584;
wire            n6585;
wire            n6586;
wire            n6587;
wire            n6588;
wire            n6589;
wire            n659;
wire            n6590;
wire            n6591;
wire            n6592;
wire            n6593;
wire            n6594;
wire            n6595;
wire            n6596;
wire            n6597;
wire            n6598;
wire            n6599;
wire            n66;
wire            n660;
wire            n6600;
wire            n6601;
wire            n6602;
wire            n6603;
wire            n6604;
wire            n6605;
wire            n6606;
wire            n6607;
wire            n6608;
wire            n6609;
wire            n661;
wire            n6610;
wire            n6611;
wire            n6612;
wire            n6613;
wire            n6614;
wire            n6615;
wire            n6616;
wire            n6617;
wire            n6618;
wire            n6619;
wire            n662;
wire            n6620;
wire            n6621;
wire            n6622;
wire            n6623;
wire            n6624;
wire            n6625;
wire            n6626;
wire            n6627;
wire            n6628;
wire            n6629;
wire            n663;
wire            n6630;
wire            n6631;
wire            n6632;
wire            n6633;
wire            n6634;
wire            n6635;
wire            n6636;
wire            n6637;
wire            n6638;
wire            n6639;
wire            n664;
wire            n6640;
wire            n6641;
wire            n6642;
wire            n6643;
wire            n6644;
wire            n6645;
wire            n6646;
wire            n6647;
wire            n6648;
wire            n6649;
wire            n665;
wire            n6650;
wire            n6651;
wire            n6652;
wire            n6653;
wire            n6654;
wire            n6655;
wire            n6656;
wire            n6657;
wire            n6658;
wire            n6659;
wire            n666;
wire            n6660;
wire            n6661;
wire            n6662;
wire            n6663;
wire            n6664;
wire            n6665;
wire            n6666;
wire            n6667;
wire            n6668;
wire            n6669;
wire            n667;
wire            n6670;
wire            n6671;
wire            n6672;
wire            n6673;
wire            n6674;
wire            n6675;
wire            n6676;
wire            n6677;
wire            n6678;
wire            n6679;
wire            n668;
wire            n6680;
wire            n6681;
wire            n6682;
wire            n6683;
wire            n6684;
wire            n6685;
wire            n6686;
wire            n6687;
wire            n6688;
wire            n6689;
wire            n669;
wire            n6690;
wire            n6691;
wire            n6692;
wire            n6693;
wire            n6694;
wire            n6695;
wire            n6696;
wire            n6697;
wire            n6698;
wire            n6699;
wire            n67;
wire            n670;
wire            n6700;
wire            n6701;
wire            n6702;
wire            n6703;
wire            n6704;
wire            n6705;
wire            n6706;
wire            n6707;
wire            n6708;
wire            n6709;
wire            n671;
wire            n6710;
wire            n6711;
wire            n6712;
wire            n6713;
wire            n6714;
wire            n6715;
wire            n6716;
wire            n6717;
wire            n6718;
wire            n6719;
wire            n672;
wire            n6720;
wire            n6721;
wire            n6722;
wire            n6723;
wire            n6724;
wire            n6725;
wire            n6726;
wire            n6727;
wire            n6728;
wire            n6729;
wire            n673;
wire            n6730;
wire            n6731;
wire            n6732;
wire            n6733;
wire            n6734;
wire            n6735;
wire            n6736;
wire            n6737;
wire            n6738;
wire            n6739;
wire            n674;
wire            n6740;
wire            n6741;
wire            n6742;
wire            n6743;
wire            n6744;
wire            n6745;
wire            n6746;
wire            n6747;
wire            n6748;
wire            n6749;
wire            n675;
wire            n6750;
wire            n6751;
wire            n6752;
wire            n6753;
wire            n6754;
wire            n6755;
wire            n6756;
wire            n6757;
wire            n6758;
wire            n6759;
wire            n676;
wire            n6760;
wire            n6761;
wire            n6762;
wire            n6763;
wire            n6764;
wire            n6765;
wire            n6766;
wire            n6767;
wire            n6768;
wire            n6769;
wire            n677;
wire            n6770;
wire            n6771;
wire            n6772;
wire            n6773;
wire            n6774;
wire            n6775;
wire            n6776;
wire            n6777;
wire            n6778;
wire            n6779;
wire            n678;
wire            n6780;
wire            n6781;
wire            n6782;
wire            n6783;
wire            n6784;
wire            n6785;
wire            n6786;
wire            n6787;
wire            n6788;
wire            n6789;
wire            n679;
wire            n6790;
wire            n6791;
wire            n6792;
wire            n6793;
wire            n6794;
wire            n6795;
wire            n6796;
wire            n6797;
wire            n6798;
wire            n6799;
wire            n68;
wire            n680;
wire            n6800;
wire            n6801;
wire            n6802;
wire            n6803;
wire            n6804;
wire            n6805;
wire            n6806;
wire            n6807;
wire            n6808;
wire            n6809;
wire            n681;
wire            n6810;
wire            n6811;
wire            n6812;
wire            n6813;
wire            n6814;
wire            n6815;
wire            n6816;
wire            n6817;
wire            n6818;
wire            n6819;
wire            n682;
wire            n6820;
wire            n6821;
wire            n6822;
wire            n6823;
wire            n6824;
wire            n6825;
wire            n6826;
wire            n6827;
wire            n6828;
wire            n6829;
wire            n683;
wire            n6830;
wire            n6831;
wire            n6832;
wire            n6833;
wire            n6834;
wire            n6835;
wire            n6836;
wire            n6837;
wire            n6838;
wire            n6839;
wire            n684;
wire            n6840;
wire            n6841;
wire            n6842;
wire            n6843;
wire            n6844;
wire            n6845;
wire            n6846;
wire            n6847;
wire            n6848;
wire            n6849;
wire            n685;
wire            n6850;
wire            n6851;
wire            n6852;
wire            n6853;
wire            n6854;
wire            n6855;
wire            n6856;
wire            n6857;
wire            n6858;
wire            n6859;
wire            n686;
wire            n6860;
wire            n6861;
wire            n6862;
wire            n6863;
wire            n6864;
wire            n6865;
wire            n6866;
wire            n6867;
wire            n6868;
wire            n6869;
wire            n687;
wire            n6870;
wire            n6871;
wire            n6872;
wire            n6873;
wire            n6874;
wire            n6875;
wire            n6876;
wire            n6877;
wire            n6878;
wire            n6879;
wire            n688;
wire            n6880;
wire            n6881;
wire            n6882;
wire            n6883;
wire            n6884;
wire            n6885;
wire            n6886;
wire            n6887;
wire            n6888;
wire            n6889;
wire            n689;
wire            n6890;
wire            n6891;
wire            n6892;
wire            n6893;
wire            n6894;
wire            n6895;
wire            n6896;
wire            n6897;
wire            n6898;
wire            n6899;
wire            n69;
wire            n690;
wire            n6900;
wire            n6901;
wire            n6902;
wire            n6903;
wire            n6904;
wire            n6905;
wire            n6906;
wire            n6907;
wire            n6908;
wire            n6909;
wire            n691;
wire            n6910;
wire            n6911;
wire            n6912;
wire            n6913;
wire            n6914;
wire            n6915;
wire            n6916;
wire            n6917;
wire            n6918;
wire            n6919;
wire            n692;
wire            n6920;
wire            n6921;
wire            n6922;
wire            n6923;
wire            n6924;
wire            n6925;
wire            n6926;
wire            n6927;
wire            n6928;
wire            n6929;
wire            n693;
wire            n6930;
wire            n6931;
wire            n6932;
wire            n6933;
wire            n6934;
wire            n6935;
wire            n6936;
wire            n6937;
wire            n6938;
wire            n6939;
wire            n694;
wire            n6940;
wire            n6941;
wire            n6942;
wire            n6943;
wire            n6944;
wire            n6945;
wire            n6946;
wire            n6947;
wire            n6948;
wire            n6949;
wire            n695;
wire            n6950;
wire            n6951;
wire            n6952;
wire            n6953;
wire            n6954;
wire            n6955;
wire            n6956;
wire            n6957;
wire            n6958;
wire            n6959;
wire            n696;
wire            n6960;
wire            n6961;
wire            n6962;
wire            n6963;
wire            n6964;
wire            n6965;
wire            n6966;
wire            n6967;
wire            n6968;
wire            n6969;
wire            n697;
wire            n6970;
wire            n6971;
wire            n6972;
wire            n6973;
wire            n6974;
wire            n6975;
wire            n6976;
wire            n6977;
wire            n6978;
wire            n6979;
wire            n698;
wire            n6980;
wire            n6981;
wire            n6982;
wire            n6983;
wire            n6984;
wire            n6985;
wire            n6986;
wire            n6987;
wire            n6988;
wire            n6989;
wire            n699;
wire            n6990;
wire            n6991;
wire            n6992;
wire            n6993;
wire            n6994;
wire            n6995;
wire            n6996;
wire            n6997;
wire            n6998;
wire            n6999;
wire            n7;
wire            n70;
wire            n700;
wire            n7000;
wire            n7001;
wire            n7002;
wire            n7003;
wire            n7004;
wire            n7005;
wire            n7006;
wire            n7007;
wire            n7008;
wire            n7009;
wire            n701;
wire            n7010;
wire            n7011;
wire            n7012;
wire            n7013;
wire            n7014;
wire            n7015;
wire            n7016;
wire            n7017;
wire            n7018;
wire            n7019;
wire            n702;
wire            n7020;
wire            n7021;
wire            n7022;
wire            n7023;
wire            n7024;
wire            n7025;
wire            n7026;
wire            n7027;
wire            n7028;
wire            n7029;
wire            n703;
wire            n7030;
wire            n7031;
wire            n7032;
wire            n7033;
wire            n7034;
wire            n7035;
wire            n7036;
wire            n7037;
wire            n7038;
wire            n7039;
wire            n704;
wire            n7040;
wire            n7041;
wire            n7042;
wire            n7043;
wire            n7044;
wire            n7045;
wire            n7046;
wire            n7047;
wire            n7048;
wire            n7049;
wire            n705;
wire            n7050;
wire            n7051;
wire            n7052;
wire            n7053;
wire            n7054;
wire            n7055;
wire            n7056;
wire            n7057;
wire            n7058;
wire            n7059;
wire            n706;
wire            n7060;
wire            n7061;
wire            n7062;
wire            n7063;
wire            n7064;
wire            n7065;
wire            n7066;
wire            n7067;
wire            n7068;
wire            n7069;
wire            n707;
wire            n7070;
wire            n7071;
wire            n7072;
wire            n7073;
wire            n7074;
wire            n7075;
wire            n7076;
wire            n7077;
wire            n7078;
wire            n7079;
wire            n708;
wire            n7080;
wire            n7081;
wire            n7082;
wire            n7083;
wire            n7084;
wire            n7085;
wire            n7086;
wire            n7087;
wire            n7088;
wire            n7089;
wire            n709;
wire            n7090;
wire            n7091;
wire            n7092;
wire            n7093;
wire            n7094;
wire            n7095;
wire            n7096;
wire            n7097;
wire            n7098;
wire            n7099;
wire            n71;
wire            n710;
wire            n7100;
wire            n7101;
wire            n7102;
wire            n7103;
wire            n7104;
wire            n7105;
wire            n7106;
wire            n7107;
wire            n7108;
wire            n7109;
wire            n711;
wire            n7110;
wire            n7111;
wire            n7112;
wire            n7113;
wire            n7114;
wire            n7115;
wire            n7116;
wire            n7117;
wire            n7118;
wire            n7119;
wire            n712;
wire            n7120;
wire            n7121;
wire            n7122;
wire            n7123;
wire            n7124;
wire            n7125;
wire            n7126;
wire            n7127;
wire            n7128;
wire            n7129;
wire            n713;
wire            n7130;
wire            n7131;
wire            n7132;
wire            n7133;
wire            n7134;
wire            n7135;
wire            n7136;
wire            n7137;
wire            n7138;
wire            n7139;
wire            n714;
wire            n7140;
wire            n7141;
wire            n7142;
wire            n7143;
wire            n7144;
wire            n7145;
wire            n7146;
wire            n7147;
wire            n7148;
wire            n7149;
wire            n715;
wire            n7150;
wire            n7151;
wire            n7152;
wire            n7153;
wire            n7154;
wire            n7155;
wire            n7156;
wire            n7157;
wire            n7158;
wire            n7159;
wire            n716;
wire            n7160;
wire            n7161;
wire            n7162;
wire            n7163;
wire            n7164;
wire            n7165;
wire            n7166;
wire            n7167;
wire            n7168;
wire            n7169;
wire            n717;
wire            n7170;
wire            n7171;
wire            n7172;
wire            n7173;
wire            n7174;
wire            n7175;
wire            n7176;
wire            n7177;
wire            n7178;
wire            n7179;
wire            n718;
wire            n7180;
wire            n7181;
wire            n7182;
wire            n7183;
wire            n7184;
wire            n7185;
wire            n7186;
wire            n7187;
wire            n7188;
wire            n7189;
wire            n719;
wire            n7190;
wire            n7191;
wire            n7192;
wire            n7193;
wire            n7194;
wire            n7195;
wire            n7196;
wire            n7197;
wire            n7198;
wire            n7199;
wire            n72;
wire            n720;
wire            n7200;
wire            n7201;
wire            n7202;
wire            n7203;
wire            n7204;
wire            n7205;
wire            n7206;
wire            n7207;
wire            n7208;
wire            n7209;
wire            n721;
wire            n7210;
wire            n7211;
wire            n7212;
wire            n7213;
wire            n7214;
wire            n7215;
wire            n7216;
wire            n7217;
wire            n7218;
wire            n7219;
wire            n722;
wire            n7220;
wire            n7221;
wire            n7222;
wire            n7223;
wire            n7224;
wire            n7225;
wire            n7226;
wire            n7227;
wire            n7228;
wire            n7229;
wire            n723;
wire            n7230;
wire            n7231;
wire            n7232;
wire            n7233;
wire            n7234;
wire            n7235;
wire            n7236;
wire            n7237;
wire            n7238;
wire            n7239;
wire            n724;
wire            n7240;
wire            n7241;
wire            n7242;
wire            n7243;
wire            n7244;
wire            n7245;
wire            n7246;
wire            n7247;
wire            n7248;
wire            n7249;
wire            n725;
wire            n7250;
wire            n7251;
wire            n7252;
wire            n7253;
wire            n7254;
wire            n7255;
wire            n7256;
wire            n7257;
wire            n7258;
wire            n7259;
wire            n726;
wire            n7260;
wire            n7261;
wire            n7262;
wire            n7263;
wire            n7264;
wire            n7265;
wire            n7266;
wire            n7267;
wire            n7268;
wire            n7269;
wire            n727;
wire            n7270;
wire            n7271;
wire            n7272;
wire            n7273;
wire            n7274;
wire            n7275;
wire            n7276;
wire            n7277;
wire            n7278;
wire            n7279;
wire            n728;
wire            n7280;
wire            n7281;
wire            n7282;
wire            n7283;
wire            n7284;
wire            n7285;
wire            n7286;
wire            n7287;
wire            n7288;
wire            n7289;
wire            n729;
wire            n7290;
wire            n7291;
wire            n7292;
wire            n7293;
wire            n7294;
wire            n7295;
wire            n7296;
wire            n7297;
wire            n7298;
wire            n7299;
wire            n73;
wire            n730;
wire            n7300;
wire            n7301;
wire            n7302;
wire            n7303;
wire            n7304;
wire            n7305;
wire            n7306;
wire            n7307;
wire            n7308;
wire            n7309;
wire            n731;
wire            n7310;
wire            n7311;
wire            n7312;
wire            n7313;
wire            n7314;
wire            n7315;
wire            n7316;
wire            n7317;
wire            n7318;
wire            n7319;
wire            n732;
wire            n7320;
wire            n7321;
wire            n7322;
wire            n7323;
wire            n7324;
wire            n7325;
wire            n7326;
wire            n7327;
wire            n7328;
wire            n7329;
wire            n733;
wire            n7330;
wire            n7331;
wire            n7332;
wire            n7333;
wire            n7334;
wire            n7335;
wire            n7336;
wire            n7337;
wire            n7338;
wire            n7339;
wire            n734;
wire            n7340;
wire            n7341;
wire            n7342;
wire            n7343;
wire            n7344;
wire            n7345;
wire            n7346;
wire            n7347;
wire            n7348;
wire            n7349;
wire            n735;
wire            n7350;
wire            n7351;
wire            n7352;
wire            n7353;
wire            n7354;
wire            n7355;
wire            n7356;
wire            n7357;
wire            n7358;
wire            n7359;
wire            n736;
wire            n7360;
wire            n7361;
wire            n7362;
wire            n7363;
wire            n7364;
wire            n7365;
wire            n7366;
wire            n7367;
wire            n7368;
wire            n7369;
wire            n737;
wire            n7370;
wire            n7371;
wire            n7372;
wire            n7373;
wire            n7374;
wire            n7375;
wire            n7376;
wire            n7377;
wire            n7378;
wire            n7379;
wire            n738;
wire            n7380;
wire            n7381;
wire            n7382;
wire            n7383;
wire            n7384;
wire            n7385;
wire            n7386;
wire            n7387;
wire            n7388;
wire            n7389;
wire            n739;
wire            n7390;
wire            n7391;
wire            n7392;
wire            n7393;
wire            n7394;
wire            n7395;
wire            n7396;
wire            n7397;
wire            n7398;
wire            n7399;
wire            n74;
wire            n740;
wire            n7400;
wire            n7401;
wire            n7402;
wire            n7403;
wire            n7404;
wire            n7405;
wire            n7406;
wire            n7407;
wire            n7408;
wire            n7409;
wire            n741;
wire            n7410;
wire            n7411;
wire            n7412;
wire            n7413;
wire            n7414;
wire            n7415;
wire            n7416;
wire            n7417;
wire            n7418;
wire            n7419;
wire            n742;
wire            n7420;
wire            n7421;
wire            n7422;
wire            n7423;
wire            n7424;
wire            n7425;
wire            n7426;
wire            n7427;
wire            n7428;
wire            n7429;
wire            n743;
wire            n7430;
wire            n7431;
wire            n7432;
wire            n7433;
wire            n7434;
wire            n7435;
wire            n7436;
wire            n7437;
wire            n7438;
wire            n7439;
wire            n744;
wire            n7440;
wire            n7441;
wire            n7442;
wire            n7443;
wire            n7444;
wire            n7445;
wire            n7446;
wire            n7447;
wire            n7448;
wire            n7449;
wire            n745;
wire            n7450;
wire            n7451;
wire            n7452;
wire            n7453;
wire            n7454;
wire            n7455;
wire            n7456;
wire            n7457;
wire            n7458;
wire            n7459;
wire            n746;
wire            n7460;
wire            n7461;
wire            n7462;
wire            n7463;
wire            n7464;
wire            n7465;
wire            n7466;
wire            n7467;
wire            n7468;
wire            n7469;
wire            n747;
wire            n7470;
wire            n7471;
wire            n7472;
wire            n7473;
wire            n7474;
wire            n7475;
wire            n7476;
wire            n7477;
wire            n7478;
wire            n7479;
wire            n748;
wire            n7480;
wire            n7481;
wire            n7482;
wire            n7483;
wire            n7484;
wire            n7485;
wire            n7486;
wire            n7487;
wire            n7488;
wire            n7489;
wire            n749;
wire            n7490;
wire            n7491;
wire            n7492;
wire            n7493;
wire            n7494;
wire            n7495;
wire            n7496;
wire            n7497;
wire            n7498;
wire            n7499;
wire            n75;
wire            n750;
wire            n7500;
wire            n7501;
wire            n7502;
wire            n7503;
wire            n7504;
wire            n7505;
wire            n7506;
wire            n7507;
wire            n7508;
wire            n7509;
wire            n751;
wire            n7510;
wire            n7511;
wire            n7512;
wire            n7513;
wire            n7514;
wire            n7515;
wire            n7516;
wire            n7517;
wire            n7518;
wire            n7519;
wire            n752;
wire            n7520;
wire            n7521;
wire            n7522;
wire            n7523;
wire            n7524;
wire            n7525;
wire            n7526;
wire            n7527;
wire            n7528;
wire            n7529;
wire            n753;
wire            n7530;
wire            n7531;
wire            n7532;
wire            n7533;
wire            n7534;
wire            n7535;
wire            n7536;
wire            n7537;
wire            n7538;
wire            n7539;
wire            n754;
wire            n7540;
wire            n7541;
wire            n7542;
wire            n7543;
wire            n7544;
wire            n7545;
wire            n7546;
wire            n7547;
wire            n7548;
wire            n7549;
wire            n755;
wire            n7550;
wire            n7551;
wire            n7552;
wire            n7553;
wire            n7554;
wire            n7555;
wire            n7556;
wire            n7557;
wire            n7558;
wire            n7559;
wire            n756;
wire            n7560;
wire            n7561;
wire            n7562;
wire            n7563;
wire            n7564;
wire            n7565;
wire            n7566;
wire            n7567;
wire            n7568;
wire            n7569;
wire            n757;
wire            n7570;
wire            n7571;
wire            n7572;
wire            n7573;
wire            n7574;
wire            n7575;
wire            n7576;
wire            n7577;
wire            n7578;
wire            n7579;
wire            n758;
wire            n7580;
wire            n7581;
wire            n7582;
wire            n7583;
wire            n7584;
wire            n7585;
wire            n7586;
wire            n7587;
wire            n7588;
wire            n7589;
wire            n759;
wire            n7590;
wire            n7591;
wire            n7592;
wire            n7593;
wire            n7594;
wire            n7595;
wire            n7596;
wire            n7597;
wire            n7598;
wire            n7599;
wire            n76;
wire            n760;
wire            n7600;
wire            n7601;
wire            n7602;
wire            n7603;
wire            n7604;
wire            n7605;
wire            n7606;
wire            n7607;
wire            n7608;
wire            n7609;
wire            n761;
wire            n7610;
wire            n7611;
wire            n7612;
wire            n7613;
wire            n7614;
wire            n7615;
wire            n7616;
wire            n7617;
wire            n7618;
wire            n7619;
wire            n762;
wire            n7620;
wire            n7621;
wire            n7622;
wire            n7623;
wire            n7624;
wire            n7625;
wire            n7626;
wire            n7627;
wire            n7628;
wire            n7629;
wire            n763;
wire            n7630;
wire            n7631;
wire            n7632;
wire            n7633;
wire            n7634;
wire            n7635;
wire            n7636;
wire            n7637;
wire            n7638;
wire            n7639;
wire            n764;
wire            n7640;
wire            n7641;
wire            n7642;
wire            n7643;
wire            n7644;
wire            n7645;
wire            n7646;
wire            n7647;
wire            n7648;
wire            n7649;
wire            n765;
wire            n7650;
wire            n7651;
wire            n7652;
wire            n7653;
wire            n7654;
wire            n7655;
wire            n7656;
wire            n7657;
wire            n7658;
wire            n7659;
wire            n766;
wire            n7660;
wire            n7661;
wire            n7662;
wire            n7663;
wire            n7664;
wire            n7665;
wire            n7666;
wire            n7667;
wire            n7668;
wire            n7669;
wire            n767;
wire            n7670;
wire            n7671;
wire            n7672;
wire            n7673;
wire            n7674;
wire            n7675;
wire            n7676;
wire            n7677;
wire            n7678;
wire            n7679;
wire            n768;
wire            n7680;
wire            n7681;
wire            n7682;
wire            n7683;
wire            n7684;
wire            n7685;
wire            n7686;
wire            n7687;
wire            n7688;
wire            n7689;
wire            n769;
wire            n7690;
wire            n7691;
wire            n7692;
wire            n7693;
wire            n7694;
wire            n7695;
wire            n7696;
wire            n7697;
wire            n7698;
wire            n7699;
wire            n77;
wire            n770;
wire            n7700;
wire            n7701;
wire            n7702;
wire            n7703;
wire            n7704;
wire            n7705;
wire            n7706;
wire            n7707;
wire            n7708;
wire            n7709;
wire            n771;
wire            n7710;
wire            n7711;
wire            n7712;
wire            n7713;
wire            n7714;
wire            n7715;
wire            n7716;
wire            n7717;
wire            n7718;
wire            n7719;
wire            n772;
wire            n7720;
wire            n7721;
wire            n7722;
wire            n7723;
wire            n7724;
wire            n7725;
wire            n7726;
wire            n7727;
wire            n7728;
wire            n7729;
wire            n773;
wire            n7730;
wire            n7731;
wire            n7732;
wire            n7733;
wire            n7734;
wire            n7735;
wire            n7736;
wire            n7737;
wire            n7738;
wire            n7739;
wire            n774;
wire            n7740;
wire            n7741;
wire            n7742;
wire            n7743;
wire            n7744;
wire            n7745;
wire            n7746;
wire            n7747;
wire            n7748;
wire            n7749;
wire            n775;
wire            n7750;
wire            n7751;
wire            n7752;
wire            n7753;
wire            n7754;
wire            n7755;
wire            n7756;
wire            n7757;
wire            n7758;
wire            n7759;
wire            n776;
wire            n7760;
wire            n7761;
wire            n7762;
wire            n7763;
wire            n7764;
wire            n7765;
wire            n7766;
wire            n7767;
wire            n7768;
wire            n7769;
wire            n777;
wire            n7770;
wire            n7771;
wire            n7772;
wire            n7773;
wire            n7774;
wire            n7775;
wire            n7776;
wire            n7777;
wire            n7778;
wire            n7779;
wire            n778;
wire            n7780;
wire            n7781;
wire            n7782;
wire            n7783;
wire            n7784;
wire            n7785;
wire            n7786;
wire            n7787;
wire            n7788;
wire            n7789;
wire            n779;
wire            n7790;
wire            n7791;
wire            n7792;
wire            n7793;
wire            n7794;
wire            n7795;
wire            n7796;
wire            n7797;
wire            n7798;
wire            n7799;
wire            n78;
wire            n780;
wire            n7800;
wire            n7801;
wire            n7802;
wire            n7803;
wire            n7804;
wire            n7805;
wire            n7806;
wire            n7807;
wire            n7808;
wire            n7809;
wire            n781;
wire            n7810;
wire            n7811;
wire            n7812;
wire            n7813;
wire            n7814;
wire            n7815;
wire            n7816;
wire            n7817;
wire            n7818;
wire            n7819;
wire            n782;
wire            n7820;
wire            n7821;
wire            n7822;
wire            n7823;
wire            n7824;
wire            n7825;
wire            n7826;
wire            n7827;
wire            n7828;
wire            n7829;
wire            n783;
wire            n7830;
wire            n7831;
wire            n7832;
wire            n7833;
wire            n7834;
wire            n7835;
wire            n7836;
wire            n7837;
wire            n7838;
wire            n7839;
wire            n784;
wire            n7840;
wire            n7841;
wire            n7842;
wire            n7843;
wire            n7844;
wire            n7845;
wire            n7846;
wire            n7847;
wire            n7848;
wire            n7849;
wire            n785;
wire            n7850;
wire            n7851;
wire            n7852;
wire            n7853;
wire            n7854;
wire            n7855;
wire            n7856;
wire            n7857;
wire            n7858;
wire            n7859;
wire            n786;
wire            n7860;
wire            n7861;
wire            n7862;
wire            n7863;
wire            n7864;
wire            n7865;
wire            n7866;
wire            n7867;
wire            n7868;
wire            n7869;
wire            n787;
wire            n7870;
wire            n7871;
wire            n7872;
wire            n7873;
wire            n7874;
wire            n7875;
wire            n7876;
wire            n7877;
wire            n7878;
wire            n7879;
wire            n788;
wire            n7880;
wire            n7881;
wire            n7882;
wire            n7883;
wire            n7884;
wire            n7885;
wire            n7886;
wire            n7887;
wire            n7888;
wire            n7889;
wire            n789;
wire            n7890;
wire            n7891;
wire            n7892;
wire            n7893;
wire            n7894;
wire            n7895;
wire            n7896;
wire            n7897;
wire            n7898;
wire            n7899;
wire            n79;
wire            n790;
wire            n7900;
wire            n7901;
wire            n7902;
wire            n7903;
wire            n7904;
wire            n7905;
wire            n7906;
wire            n7907;
wire            n7908;
wire            n7909;
wire            n791;
wire            n7910;
wire            n7911;
wire            n7912;
wire            n7913;
wire            n7914;
wire            n7915;
wire            n7916;
wire            n7917;
wire            n7918;
wire            n7919;
wire            n792;
wire            n7920;
wire            n7921;
wire            n7922;
wire            n7923;
wire            n7924;
wire            n7925;
wire            n7926;
wire            n7927;
wire            n7928;
wire            n7929;
wire            n793;
wire            n7930;
wire            n7931;
wire            n7932;
wire            n7933;
wire            n7934;
wire            n7935;
wire            n7936;
wire            n7937;
wire            n7938;
wire            n7939;
wire            n794;
wire            n7940;
wire            n7941;
wire            n7942;
wire            n7943;
wire            n7944;
wire            n7945;
wire            n7946;
wire            n7947;
wire            n7948;
wire            n7949;
wire            n795;
wire            n7950;
wire            n7951;
wire            n7952;
wire            n7953;
wire            n7954;
wire            n7955;
wire            n7956;
wire            n7957;
wire            n7958;
wire            n7959;
wire            n796;
wire            n7960;
wire            n7961;
wire            n7962;
wire            n7963;
wire            n7964;
wire            n7965;
wire            n7966;
wire            n7967;
wire            n7968;
wire            n7969;
wire            n797;
wire            n7970;
wire            n7971;
wire            n7972;
wire            n7973;
wire            n7974;
wire            n7975;
wire            n7976;
wire            n7977;
wire            n7978;
wire            n7979;
wire            n798;
wire            n7980;
wire            n7981;
wire            n7982;
wire            n7983;
wire            n7984;
wire            n7985;
wire            n7986;
wire            n7987;
wire            n7988;
wire            n7989;
wire            n799;
wire            n7990;
wire            n7991;
wire            n7992;
wire            n7993;
wire            n7994;
wire            n7995;
wire            n7996;
wire            n7997;
wire            n7998;
wire            n7999;
wire            n8;
wire            n80;
wire            n800;
wire            n8000;
wire            n8001;
wire            n8002;
wire            n8003;
wire            n8004;
wire            n8005;
wire            n8006;
wire            n8007;
wire            n8008;
wire            n8009;
wire            n801;
wire            n8010;
wire            n8011;
wire            n8012;
wire            n8013;
wire            n8014;
wire            n8015;
wire            n8016;
wire            n8017;
wire            n8018;
wire            n8019;
wire            n802;
wire            n8020;
wire            n8021;
wire            n8022;
wire            n8023;
wire            n8024;
wire            n8025;
wire            n8026;
wire            n8027;
wire            n8028;
wire            n8029;
wire            n803;
wire            n8030;
wire            n8031;
wire            n8032;
wire            n8033;
wire            n8034;
wire            n8035;
wire            n8036;
wire            n8037;
wire            n8038;
wire            n8039;
wire            n804;
wire            n8040;
wire            n8041;
wire            n8042;
wire            n8043;
wire            n8044;
wire            n8045;
wire            n8046;
wire            n8047;
wire            n8048;
wire            n8049;
wire            n805;
wire            n8050;
wire            n8051;
wire            n8052;
wire            n8053;
wire            n8054;
wire            n8055;
wire            n8056;
wire            n8057;
wire            n8058;
wire            n8059;
wire            n806;
wire            n8060;
wire            n8061;
wire            n8062;
wire            n8063;
wire            n8064;
wire            n8065;
wire            n8066;
wire            n8067;
wire            n8068;
wire            n8069;
wire            n807;
wire            n8070;
wire            n8071;
wire            n8072;
wire            n8073;
wire            n8074;
wire            n8075;
wire            n8076;
wire            n8077;
wire            n8078;
wire            n8079;
wire            n808;
wire            n8080;
wire            n8081;
wire            n8082;
wire            n8083;
wire            n8084;
wire            n8085;
wire            n8086;
wire            n8087;
wire            n8088;
wire            n8089;
wire            n809;
wire            n8090;
wire            n8091;
wire            n8092;
wire            n8093;
wire            n8094;
wire            n8095;
wire            n8096;
wire            n8097;
wire            n8098;
wire            n8099;
wire            n81;
wire            n810;
wire            n8100;
wire            n8101;
wire            n8102;
wire            n8103;
wire            n8104;
wire            n8105;
wire            n8106;
wire            n8107;
wire            n8108;
wire            n8109;
wire            n811;
wire            n8110;
wire            n8111;
wire            n8112;
wire            n8113;
wire            n8114;
wire            n8115;
wire            n8116;
wire            n8117;
wire            n8118;
wire            n8119;
wire            n812;
wire            n8120;
wire            n8121;
wire            n8122;
wire            n8123;
wire            n8124;
wire            n8125;
wire            n8126;
wire            n8127;
wire            n8128;
wire            n8129;
wire            n813;
wire            n8130;
wire            n8131;
wire            n8132;
wire            n8133;
wire            n8134;
wire            n8135;
wire            n8136;
wire            n8137;
wire            n8138;
wire            n8139;
wire            n814;
wire            n8140;
wire            n8141;
wire            n8142;
wire            n8143;
wire            n8144;
wire            n8145;
wire            n8146;
wire            n8147;
wire            n8148;
wire            n8149;
wire            n815;
wire            n8150;
wire            n8151;
wire            n8152;
wire            n8153;
wire            n8154;
wire            n8155;
wire            n8156;
wire            n8157;
wire            n8158;
wire            n8159;
wire            n816;
wire            n8160;
wire            n8161;
wire            n8162;
wire            n8163;
wire            n8164;
wire            n8165;
wire            n8166;
wire            n8167;
wire            n8168;
wire            n8169;
wire            n817;
wire            n8170;
wire            n8171;
wire            n8172;
wire            n8173;
wire            n8174;
wire            n8175;
wire            n8176;
wire            n8177;
wire            n8178;
wire            n8179;
wire            n818;
wire            n8180;
wire            n8181;
wire            n8182;
wire            n8183;
wire            n8184;
wire            n8185;
wire            n8186;
wire            n8187;
wire            n8188;
wire            n8189;
wire            n819;
wire            n8190;
wire            n8191;
wire            n8192;
wire            n8193;
wire            n8194;
wire            n8195;
wire            n8196;
wire            n8197;
wire            n8198;
wire            n8199;
wire            n82;
wire            n820;
wire            n8200;
wire            n8201;
wire            n8202;
wire            n8203;
wire            n8204;
wire            n8205;
wire            n8206;
wire            n8207;
wire            n8208;
wire            n8209;
wire            n821;
wire            n8210;
wire            n8211;
wire            n8212;
wire            n8213;
wire            n8214;
wire            n8215;
wire            n8216;
wire            n8217;
wire            n8218;
wire            n8219;
wire            n822;
wire            n8220;
wire            n8221;
wire            n8222;
wire            n8223;
wire            n8224;
wire            n8225;
wire            n8226;
wire            n8227;
wire            n8228;
wire            n8229;
wire            n823;
wire            n8230;
wire            n8231;
wire            n8232;
wire            n8233;
wire            n8234;
wire            n8235;
wire            n8236;
wire            n8237;
wire            n8238;
wire            n8239;
wire            n824;
wire            n8240;
wire            n8241;
wire            n8242;
wire            n8243;
wire            n8244;
wire            n8245;
wire            n8246;
wire            n8247;
wire            n8248;
wire            n8249;
wire            n825;
wire            n8250;
wire            n8251;
wire            n8252;
wire            n8253;
wire            n8254;
wire            n8255;
wire            n8256;
wire            n8257;
wire            n8258;
wire            n8259;
wire            n826;
wire            n8260;
wire            n8261;
wire            n8262;
wire            n8263;
wire            n8264;
wire            n8265;
wire            n8266;
wire            n8267;
wire            n8268;
wire            n8269;
wire            n827;
wire            n8270;
wire            n8271;
wire            n8272;
wire            n8273;
wire            n8274;
wire            n8275;
wire            n8276;
wire            n8277;
wire            n8278;
wire            n8279;
wire            n828;
wire            n8280;
wire            n8281;
wire            n8282;
wire            n8283;
wire            n8284;
wire            n8285;
wire            n8286;
wire            n8287;
wire            n8288;
wire            n8289;
wire            n829;
wire            n8290;
wire            n8291;
wire            n8292;
wire            n8293;
wire            n8294;
wire            n8295;
wire            n8296;
wire            n8297;
wire            n8298;
wire            n8299;
wire            n83;
wire            n830;
wire            n8300;
wire            n8301;
wire            n8302;
wire            n8303;
wire            n8304;
wire            n8305;
wire            n8306;
wire            n8307;
wire            n8308;
wire            n8309;
wire            n831;
wire            n8310;
wire            n8311;
wire            n8312;
wire            n8313;
wire            n8314;
wire            n8315;
wire            n8316;
wire            n8317;
wire            n8318;
wire            n8319;
wire            n832;
wire            n8320;
wire            n8321;
wire            n8322;
wire            n8323;
wire            n8324;
wire            n8325;
wire            n8326;
wire            n8327;
wire            n8328;
wire            n8329;
wire            n833;
wire            n8330;
wire            n8331;
wire            n8332;
wire            n8333;
wire            n8334;
wire            n8335;
wire            n8336;
wire            n8337;
wire            n8338;
wire            n8339;
wire            n834;
wire            n8340;
wire            n8341;
wire            n8342;
wire            n8343;
wire            n8344;
wire            n8345;
wire            n8346;
wire            n8347;
wire            n8348;
wire            n8349;
wire            n835;
wire            n8350;
wire            n8351;
wire            n8352;
wire            n8353;
wire            n8354;
wire            n8355;
wire            n8356;
wire            n8357;
wire            n8358;
wire            n8359;
wire            n836;
wire            n8360;
wire            n8361;
wire            n8362;
wire            n8363;
wire            n8364;
wire            n8365;
wire            n8366;
wire            n8367;
wire            n8368;
wire            n8369;
wire            n837;
wire            n8370;
wire            n8371;
wire            n8372;
wire            n8373;
wire            n8374;
wire            n8375;
wire            n8376;
wire            n8377;
wire            n8378;
wire            n8379;
wire            n838;
wire            n8380;
wire            n8381;
wire            n8382;
wire            n8383;
wire            n8384;
wire            n8385;
wire            n8386;
wire            n8387;
wire            n8388;
wire            n8389;
wire            n839;
wire            n8390;
wire            n8391;
wire            n8392;
wire            n8393;
wire            n8394;
wire            n8395;
wire            n8396;
wire            n8397;
wire            n8398;
wire            n8399;
wire            n84;
wire            n840;
wire            n8400;
wire            n8401;
wire            n8402;
wire            n8403;
wire            n8404;
wire            n8405;
wire            n8406;
wire            n8407;
wire            n8408;
wire            n8409;
wire            n841;
wire            n8410;
wire            n8411;
wire            n8412;
wire            n8413;
wire            n8414;
wire            n8415;
wire            n8416;
wire            n8417;
wire            n8418;
wire            n8419;
wire            n842;
wire            n8420;
wire            n8421;
wire            n8422;
wire            n8423;
wire            n8424;
wire            n8425;
wire            n8426;
wire            n8427;
wire            n8428;
wire            n8429;
wire            n843;
wire            n8430;
wire            n8431;
wire            n8432;
wire            n8433;
wire            n8434;
wire            n8435;
wire            n8436;
wire            n8437;
wire            n8438;
wire            n8439;
wire            n844;
wire            n8440;
wire            n8441;
wire            n8442;
wire            n8443;
wire            n8444;
wire            n8445;
wire            n8446;
wire            n8447;
wire            n8448;
wire            n8449;
wire            n845;
wire            n8450;
wire            n8451;
wire            n8452;
wire            n8453;
wire            n8454;
wire            n8455;
wire            n8456;
wire            n8457;
wire            n8458;
wire            n8459;
wire            n846;
wire            n8460;
wire            n8461;
wire            n8462;
wire            n8463;
wire            n8464;
wire            n8465;
wire            n8466;
wire            n8467;
wire            n8468;
wire            n8469;
wire            n847;
wire            n8470;
wire            n8471;
wire            n8472;
wire            n8473;
wire            n8474;
wire            n8475;
wire            n8476;
wire            n8477;
wire            n8478;
wire            n8479;
wire            n848;
wire            n8480;
wire            n8481;
wire            n8482;
wire            n8483;
wire            n8484;
wire            n8485;
wire            n8486;
wire            n8487;
wire            n8488;
wire            n8489;
wire            n849;
wire            n8490;
wire            n8491;
wire            n8492;
wire            n8493;
wire            n8494;
wire            n8495;
wire            n8496;
wire            n8497;
wire            n8498;
wire            n8499;
wire            n85;
wire            n850;
wire            n8500;
wire            n8501;
wire            n8502;
wire            n8503;
wire            n8504;
wire            n8505;
wire            n8506;
wire            n8507;
wire            n8508;
wire            n8509;
wire            n851;
wire            n8510;
wire            n8511;
wire            n8512;
wire            n8513;
wire            n8514;
wire            n8515;
wire            n8516;
wire            n8517;
wire            n8518;
wire            n8519;
wire            n852;
wire            n8520;
wire            n8521;
wire            n8522;
wire            n8523;
wire            n8524;
wire            n8525;
wire            n8526;
wire            n8527;
wire            n8528;
wire            n8529;
wire            n853;
wire            n8530;
wire            n8531;
wire            n8532;
wire            n8533;
wire            n8534;
wire            n8535;
wire            n8536;
wire            n8537;
wire            n8538;
wire            n8539;
wire            n854;
wire            n8540;
wire            n8541;
wire            n8542;
wire            n8543;
wire            n8544;
wire            n8545;
wire            n8546;
wire            n8547;
wire            n8548;
wire            n8549;
wire            n855;
wire            n8550;
wire            n8551;
wire            n8552;
wire            n8553;
wire            n8554;
wire            n8555;
wire            n8556;
wire            n8557;
wire            n8558;
wire            n8559;
wire            n856;
wire            n8560;
wire            n8561;
wire            n8562;
wire            n8563;
wire            n8564;
wire            n8565;
wire            n8566;
wire            n8567;
wire            n8568;
wire            n8569;
wire            n857;
wire            n8570;
wire            n8571;
wire            n8572;
wire            n8573;
wire            n8574;
wire            n8575;
wire            n8576;
wire            n8577;
wire            n8578;
wire            n8579;
wire            n858;
wire            n8580;
wire            n8581;
wire            n8582;
wire            n8583;
wire            n8584;
wire            n8585;
wire            n8586;
wire            n8587;
wire            n8588;
wire            n8589;
wire            n859;
wire            n8590;
wire            n8591;
wire            n8592;
wire            n8593;
wire            n8594;
wire            n8595;
wire            n8596;
wire            n8597;
wire            n8598;
wire            n8599;
wire            n86;
wire            n860;
wire            n8600;
wire            n8601;
wire            n8602;
wire            n8603;
wire            n8604;
wire            n8605;
wire            n8606;
wire            n8607;
wire            n8608;
wire            n8609;
wire            n861;
wire            n8610;
wire            n8611;
wire            n8612;
wire            n8613;
wire            n8614;
wire            n8615;
wire            n8616;
wire            n8617;
wire            n8618;
wire            n8619;
wire            n862;
wire            n8620;
wire            n8621;
wire            n8622;
wire            n8623;
wire            n8624;
wire            n8625;
wire            n8626;
wire            n8627;
wire            n8628;
wire            n8629;
wire            n863;
wire            n8630;
wire            n8631;
wire            n8632;
wire            n8633;
wire            n8634;
wire            n8635;
wire            n8636;
wire            n8637;
wire            n8638;
wire            n8639;
wire            n864;
wire            n8640;
wire            n8641;
wire            n8642;
wire            n8643;
wire            n8644;
wire            n8645;
wire            n8646;
wire            n8647;
wire            n8648;
wire            n8649;
wire            n865;
wire            n8650;
wire            n8651;
wire            n8652;
wire            n8653;
wire            n8654;
wire            n8655;
wire            n8656;
wire            n8657;
wire            n8658;
wire            n8659;
wire            n866;
wire            n8660;
wire            n8661;
wire            n8662;
wire            n8663;
wire            n8664;
wire            n8665;
wire            n8666;
wire            n8667;
wire            n8668;
wire            n8669;
wire            n867;
wire            n8670;
wire            n8671;
wire            n8672;
wire            n8673;
wire            n8674;
wire            n8675;
wire            n8676;
wire            n8677;
wire            n8678;
wire            n8679;
wire            n868;
wire            n8680;
wire            n8681;
wire            n8682;
wire            n8683;
wire            n8684;
wire            n8685;
wire            n8686;
wire            n8687;
wire            n8688;
wire            n8689;
wire            n869;
wire            n8690;
wire            n8691;
wire            n8692;
wire            n8693;
wire            n8694;
wire            n8695;
wire            n8696;
wire            n8697;
wire            n8698;
wire            n8699;
wire            n87;
wire            n870;
wire            n8700;
wire            n8701;
wire            n8702;
wire            n8703;
wire            n8704;
wire            n8705;
wire            n8706;
wire            n8707;
wire            n8708;
wire            n8709;
wire            n871;
wire            n8710;
wire            n8711;
wire            n8712;
wire            n8713;
wire            n8714;
wire            n8715;
wire            n8716;
wire            n8717;
wire            n8718;
wire            n8719;
wire            n872;
wire            n8720;
wire            n8721;
wire            n8722;
wire            n8723;
wire            n8724;
wire            n8725;
wire            n8726;
wire            n8727;
wire            n8728;
wire            n8729;
wire            n873;
wire            n8730;
wire            n8731;
wire            n8732;
wire            n8733;
wire            n8734;
wire            n8735;
wire            n8736;
wire            n8737;
wire            n8738;
wire            n8739;
wire            n874;
wire            n8740;
wire            n8741;
wire            n8742;
wire            n8743;
wire            n8744;
wire            n8745;
wire            n8746;
wire            n8747;
wire            n8748;
wire            n8749;
wire            n875;
wire            n8750;
wire            n8751;
wire            n8752;
wire            n8753;
wire            n8754;
wire            n8755;
wire            n8756;
wire            n8757;
wire            n8758;
wire            n8759;
wire            n876;
wire            n8760;
wire            n8761;
wire            n8762;
wire            n8763;
wire            n8764;
wire            n8765;
wire            n8766;
wire            n8767;
wire            n8768;
wire            n8769;
wire            n877;
wire            n8770;
wire            n8771;
wire            n8772;
wire            n8773;
wire            n8774;
wire            n8775;
wire            n8776;
wire            n8777;
wire            n8778;
wire            n8779;
wire            n878;
wire            n8780;
wire            n8781;
wire            n8782;
wire            n8783;
wire            n8784;
wire            n8785;
wire            n8786;
wire            n8787;
wire            n8788;
wire            n8789;
wire            n879;
wire            n8790;
wire            n8791;
wire            n8792;
wire            n8793;
wire            n8794;
wire            n8795;
wire            n8796;
wire            n8797;
wire            n8798;
wire            n8799;
wire            n88;
wire            n880;
wire            n8800;
wire            n8801;
wire            n8802;
wire            n8803;
wire            n8804;
wire            n8805;
wire            n8806;
wire            n8807;
wire            n8808;
wire            n8809;
wire            n881;
wire            n8810;
wire            n8811;
wire            n8812;
wire            n8813;
wire            n8814;
wire            n8815;
wire            n8816;
wire            n8817;
wire            n8818;
wire            n8819;
wire            n882;
wire            n8820;
wire            n8821;
wire            n8822;
wire            n8823;
wire            n8824;
wire            n8825;
wire            n8826;
wire            n8827;
wire            n8828;
wire            n8829;
wire            n883;
wire            n8830;
wire            n8831;
wire            n8832;
wire            n8833;
wire            n8834;
wire            n8835;
wire            n8836;
wire            n8837;
wire            n8838;
wire            n8839;
wire            n884;
wire            n8840;
wire            n8841;
wire            n8842;
wire            n8843;
wire            n8844;
wire            n8845;
wire            n8846;
wire            n8847;
wire            n8848;
wire            n8849;
wire            n885;
wire            n8850;
wire            n8851;
wire            n8852;
wire            n8853;
wire            n8854;
wire            n8855;
wire            n8856;
wire            n8857;
wire            n8858;
wire            n8859;
wire            n886;
wire            n8860;
wire            n8861;
wire            n8862;
wire            n8863;
wire            n8864;
wire            n8865;
wire            n8866;
wire            n8867;
wire            n8868;
wire            n8869;
wire            n887;
wire            n8870;
wire            n8871;
wire            n8872;
wire            n8873;
wire            n8874;
wire            n8875;
wire            n8876;
wire            n8877;
wire            n8878;
wire            n8879;
wire            n888;
wire            n8880;
wire            n8881;
wire            n8882;
wire            n8883;
wire            n8884;
wire            n8885;
wire            n8886;
wire            n8887;
wire            n8888;
wire            n8889;
wire            n889;
wire            n8890;
wire            n8891;
wire            n8892;
wire            n8893;
wire            n8894;
wire            n8895;
wire            n8896;
wire            n8897;
wire            n8898;
wire            n8899;
wire            n89;
wire            n890;
wire            n8900;
wire            n8901;
wire            n8902;
wire            n8903;
wire            n8904;
wire            n8905;
wire            n8906;
wire            n8907;
wire            n8908;
wire            n8909;
wire            n891;
wire            n8910;
wire            n8911;
wire            n8912;
wire            n8913;
wire            n8914;
wire            n8915;
wire            n8916;
wire            n8917;
wire            n8918;
wire            n8919;
wire            n892;
wire            n8920;
wire            n8921;
wire            n8922;
wire            n8923;
wire            n8924;
wire            n8925;
wire            n8926;
wire            n8927;
wire            n8928;
wire            n8929;
wire            n893;
wire            n8930;
wire            n8931;
wire            n8932;
wire            n8933;
wire            n8934;
wire            n8935;
wire            n8936;
wire            n8937;
wire            n8938;
wire            n8939;
wire            n894;
wire            n8940;
wire            n8941;
wire            n8942;
wire            n8943;
wire            n8944;
wire            n8945;
wire            n8946;
wire            n8947;
wire            n8948;
wire            n8949;
wire            n895;
wire            n8950;
wire            n8951;
wire            n8952;
wire            n8953;
wire            n8954;
wire            n8955;
wire            n8956;
wire            n8957;
wire            n8958;
wire            n8959;
wire            n896;
wire            n8960;
wire            n8961;
wire            n8962;
wire            n8963;
wire            n8964;
wire            n8965;
wire            n8966;
wire            n8967;
wire            n8968;
wire            n8969;
wire            n897;
wire            n8970;
wire            n8971;
wire            n8972;
wire            n8973;
wire            n8974;
wire            n8975;
wire            n8976;
wire            n8977;
wire            n8978;
wire            n8979;
wire            n898;
wire            n8980;
wire            n8981;
wire            n8982;
wire            n8983;
wire            n8984;
wire            n8985;
wire            n8986;
wire            n8987;
wire            n8988;
wire            n8989;
wire            n899;
wire            n8990;
wire            n8991;
wire            n8992;
wire            n8993;
wire            n8994;
wire            n8995;
wire            n8996;
wire            n8997;
wire            n8998;
wire            n8999;
wire            n9;
wire            n90;
wire            n900;
wire            n9000;
wire            n9001;
wire            n9002;
wire            n9003;
wire            n9004;
wire            n9005;
wire            n9006;
wire            n9007;
wire            n9008;
wire            n9009;
wire            n901;
wire            n9010;
wire            n9011;
wire            n9012;
wire            n9013;
wire            n9014;
wire            n9015;
wire            n9016;
wire            n9017;
wire            n9018;
wire            n9019;
wire            n902;
wire            n9020;
wire            n9021;
wire            n9022;
wire            n9023;
wire            n9024;
wire            n9025;
wire            n9026;
wire            n9027;
wire            n9028;
wire            n9029;
wire            n903;
wire            n9030;
wire            n9031;
wire            n9032;
wire            n9033;
wire            n9034;
wire            n9035;
wire            n9036;
wire            n9037;
wire            n9038;
wire            n9039;
wire            n904;
wire            n9040;
wire            n9041;
wire            n9042;
wire            n9043;
wire            n9044;
wire            n9045;
wire            n9046;
wire            n9047;
wire            n9048;
wire            n9049;
wire            n905;
wire            n9050;
wire            n9051;
wire            n9052;
wire            n9053;
wire            n9054;
wire            n9055;
wire            n9056;
wire            n9057;
wire            n9058;
wire            n9059;
wire            n906;
wire            n9060;
wire            n9061;
wire            n9062;
wire            n9063;
wire            n9064;
wire            n9065;
wire            n9066;
wire            n9067;
wire            n9068;
wire            n9069;
wire            n907;
wire            n9070;
wire            n9071;
wire            n9072;
wire            n9073;
wire            n9074;
wire            n9075;
wire            n9076;
wire            n9077;
wire            n9078;
wire            n9079;
wire            n908;
wire            n9080;
wire            n9081;
wire            n9082;
wire            n9083;
wire            n9084;
wire            n9085;
wire            n9086;
wire            n9087;
wire            n9088;
wire            n9089;
wire            n909;
wire            n9090;
wire            n9091;
wire            n9092;
wire            n9093;
wire            n9094;
wire            n9095;
wire            n9096;
wire            n9097;
wire            n9098;
wire            n9099;
wire            n91;
wire            n910;
wire            n9100;
wire            n9101;
wire            n9102;
wire            n9103;
wire            n9104;
wire            n9105;
wire            n9106;
wire            n9107;
wire            n9108;
wire            n9109;
wire            n911;
wire            n9110;
wire            n9111;
wire            n9112;
wire            n9113;
wire            n9114;
wire            n9115;
wire            n9116;
wire            n9117;
wire            n9118;
wire            n9119;
wire            n912;
wire            n9120;
wire            n9121;
wire            n9122;
wire            n9123;
wire            n9124;
wire            n9125;
wire            n9126;
wire            n9127;
wire            n9128;
wire            n9129;
wire            n913;
wire            n9130;
wire            n9131;
wire            n9132;
wire            n9133;
wire            n9134;
wire            n9135;
wire            n9136;
wire            n9137;
wire            n9138;
wire            n9139;
wire            n914;
wire            n9140;
wire            n9141;
wire            n9142;
wire            n9143;
wire            n9144;
wire            n9145;
wire            n9146;
wire            n9147;
wire            n9148;
wire            n9149;
wire            n915;
wire            n9150;
wire            n9151;
wire            n9152;
wire            n9153;
wire            n9154;
wire            n9155;
wire            n9156;
wire            n9157;
wire            n9158;
wire            n9159;
wire            n916;
wire            n9160;
wire            n9161;
wire            n9162;
wire            n9163;
wire            n9164;
wire            n9165;
wire            n9166;
wire            n9167;
wire            n9168;
wire            n9169;
wire            n917;
wire            n9170;
wire            n9171;
wire            n9172;
wire            n9173;
wire            n9174;
wire            n9175;
wire            n9176;
wire            n9177;
wire            n9178;
wire            n9179;
wire            n918;
wire            n9180;
wire            n9181;
wire            n9182;
wire            n9183;
wire            n9184;
wire            n9185;
wire            n9186;
wire            n9187;
wire            n9188;
wire            n9189;
wire            n919;
wire            n9190;
wire            n9191;
wire            n9192;
wire            n9193;
wire            n9194;
wire            n9195;
wire            n9196;
wire            n9197;
wire            n9198;
wire            n9199;
wire            n92;
wire            n920;
wire            n9200;
wire            n9201;
wire            n9202;
wire            n9203;
wire            n9204;
wire            n9205;
wire            n9206;
wire            n9207;
wire            n9208;
wire            n9209;
wire            n921;
wire            n9210;
wire            n9211;
wire            n9212;
wire            n9213;
wire            n9214;
wire            n9215;
wire            n9216;
wire            n9217;
wire            n9218;
wire            n9219;
wire            n922;
wire            n9220;
wire            n9221;
wire            n9222;
wire            n9223;
wire            n9224;
wire            n9225;
wire            n9226;
wire            n9227;
wire            n9228;
wire            n9229;
wire            n923;
wire            n9230;
wire            n9231;
wire            n9232;
wire            n9233;
wire            n9234;
wire            n9235;
wire            n9236;
wire            n9237;
wire            n9238;
wire            n9239;
wire            n924;
wire            n9240;
wire            n9241;
wire            n9242;
wire            n9243;
wire            n9244;
wire            n9245;
wire            n9246;
wire            n9247;
wire            n9248;
wire            n9249;
wire            n925;
wire            n9250;
wire            n9251;
wire            n9252;
wire            n9253;
wire            n9254;
wire            n9255;
wire            n9256;
wire            n9257;
wire            n9258;
wire            n9259;
wire            n926;
wire            n9260;
wire            n9261;
wire            n9262;
wire            n9263;
wire            n9264;
wire            n9265;
wire            n9266;
wire            n9267;
wire            n9268;
wire            n9269;
wire            n927;
wire            n9270;
wire            n9271;
wire            n9272;
wire            n9273;
wire            n9274;
wire            n9275;
wire            n9276;
wire            n9277;
wire            n9278;
wire            n9279;
wire            n928;
wire            n9280;
wire            n9281;
wire            n9282;
wire            n9283;
wire            n9284;
wire            n9285;
wire            n9286;
wire            n9287;
wire            n9288;
wire            n9289;
wire            n929;
wire            n9290;
wire            n9291;
wire            n9292;
wire            n9293;
wire            n9294;
wire            n9295;
wire            n9296;
wire            n9297;
wire            n9298;
wire            n9299;
wire            n93;
wire            n930;
wire            n9300;
wire            n9301;
wire            n9302;
wire            n9303;
wire            n9304;
wire            n9305;
wire            n9306;
wire            n9307;
wire            n9308;
wire            n9309;
wire            n931;
wire            n9310;
wire            n9311;
wire            n9312;
wire            n9313;
wire            n9314;
wire            n9315;
wire            n9316;
wire            n9317;
wire            n9318;
wire            n9319;
wire            n932;
wire            n9320;
wire            n9321;
wire            n9322;
wire            n9323;
wire            n9324;
wire            n9325;
wire            n9326;
wire            n9327;
wire            n9328;
wire            n9329;
wire            n933;
wire            n9330;
wire            n9331;
wire            n9332;
wire            n9333;
wire            n9334;
wire            n9335;
wire            n9336;
wire            n9337;
wire            n9338;
wire            n9339;
wire            n934;
wire            n9340;
wire            n9341;
wire            n9342;
wire            n9343;
wire            n9344;
wire            n9345;
wire            n9346;
wire            n9347;
wire            n9348;
wire            n9349;
wire            n935;
wire            n9350;
wire            n9351;
wire            n9352;
wire            n9353;
wire            n9354;
wire            n9355;
wire            n9356;
wire            n9357;
wire            n9358;
wire            n9359;
wire            n936;
wire            n9360;
wire            n9361;
wire            n9362;
wire            n9363;
wire            n9364;
wire            n9365;
wire            n9366;
wire            n9367;
wire            n9368;
wire            n9369;
wire            n937;
wire            n9370;
wire            n9371;
wire            n9372;
wire            n9373;
wire            n9374;
wire            n9375;
wire            n9376;
wire            n9377;
wire            n9378;
wire            n9379;
wire            n938;
wire            n9380;
wire            n9381;
wire            n9382;
wire            n9383;
wire            n9384;
wire            n9385;
wire            n9386;
wire            n9387;
wire            n9388;
wire            n9389;
wire            n939;
wire            n9390;
wire            n9391;
wire            n9392;
wire            n9393;
wire            n9394;
wire            n9395;
wire            n9396;
wire            n9397;
wire            n9398;
wire            n9399;
wire            n94;
wire            n940;
wire            n9400;
wire            n9401;
wire            n9402;
wire            n9403;
wire            n9404;
wire            n9405;
wire            n9406;
wire            n9407;
wire            n9408;
wire            n9409;
wire            n941;
wire            n9410;
wire            n9411;
wire            n9412;
wire            n9413;
wire            n9414;
wire            n9415;
wire            n9416;
wire            n9417;
wire            n9418;
wire            n9419;
wire            n942;
wire            n9420;
wire            n9421;
wire            n9422;
wire            n9423;
wire            n9424;
wire            n9425;
wire            n9426;
wire            n9427;
wire            n9428;
wire            n9429;
wire            n943;
wire            n9430;
wire            n9431;
wire            n9432;
wire            n9433;
wire            n9434;
wire            n9435;
wire            n9436;
wire            n9437;
wire            n9438;
wire            n9439;
wire            n944;
wire            n9440;
wire            n9441;
wire            n9442;
wire            n9443;
wire            n9444;
wire            n9445;
wire            n9446;
wire            n9447;
wire            n9448;
wire            n9449;
wire            n945;
wire            n9450;
wire            n9451;
wire            n9452;
wire            n9453;
wire            n9454;
wire            n9455;
wire            n9456;
wire            n9457;
wire            n9458;
wire            n9459;
wire            n946;
wire            n9460;
wire            n9461;
wire            n9462;
wire            n9463;
wire            n9464;
wire            n9465;
wire            n9466;
wire            n9467;
wire            n9468;
wire            n9469;
wire            n947;
wire            n9470;
wire            n9471;
wire            n9472;
wire            n9473;
wire            n9474;
wire            n9475;
wire            n9476;
wire            n9477;
wire            n9478;
wire            n9479;
wire            n948;
wire            n9480;
wire            n9481;
wire            n9482;
wire            n9483;
wire            n9484;
wire            n9485;
wire            n9486;
wire            n9487;
wire            n9488;
wire            n9489;
wire            n949;
wire            n9490;
wire            n9491;
wire            n9492;
wire            n9493;
wire            n9494;
wire            n9495;
wire            n9496;
wire            n9497;
wire            n9498;
wire            n9499;
wire            n95;
wire            n950;
wire            n9500;
wire            n9501;
wire            n9502;
wire            n9503;
wire            n9504;
wire            n9505;
wire            n9506;
wire            n9507;
wire            n9508;
wire            n9509;
wire            n951;
wire            n9510;
wire            n9511;
wire            n9512;
wire            n9513;
wire            n9514;
wire            n9515;
wire            n9516;
wire            n9517;
wire            n9518;
wire            n9519;
wire            n952;
wire            n9520;
wire            n9521;
wire            n9522;
wire            n9523;
wire            n9524;
wire            n9525;
wire            n9526;
wire            n9527;
wire            n9528;
wire            n9529;
wire            n953;
wire            n9530;
wire            n9531;
wire            n9532;
wire            n9533;
wire            n9534;
wire            n9535;
wire            n9536;
wire            n9537;
wire            n9538;
wire            n9539;
wire            n954;
wire            n9540;
wire            n9541;
wire            n9542;
wire            n9543;
wire            n9544;
wire            n9545;
wire            n9546;
wire            n9547;
wire            n9548;
wire            n9549;
wire            n955;
wire            n9550;
wire            n9551;
wire            n9552;
wire            n9553;
wire            n9554;
wire            n9555;
wire            n9556;
wire            n9557;
wire            n9558;
wire            n9559;
wire            n956;
wire            n9560;
wire            n9561;
wire            n9562;
wire            n9563;
wire            n9564;
wire            n9565;
wire            n9566;
wire            n9567;
wire            n9568;
wire            n9569;
wire            n957;
wire            n9570;
wire            n9571;
wire            n9572;
wire            n9573;
wire            n9574;
wire            n9575;
wire            n9576;
wire            n9577;
wire            n9578;
wire            n9579;
wire            n958;
wire            n9580;
wire            n9581;
wire            n9582;
wire            n9583;
wire            n9584;
wire            n9585;
wire            n9586;
wire            n9587;
wire            n9588;
wire            n9589;
wire            n959;
wire            n9590;
wire            n9591;
wire            n9592;
wire            n9593;
wire            n9594;
wire            n9595;
wire            n9596;
wire            n9597;
wire            n9598;
wire            n9599;
wire            n96;
wire            n960;
wire            n9600;
wire            n9601;
wire            n9602;
wire            n9603;
wire            n9604;
wire            n9605;
wire            n9606;
wire            n9607;
wire            n9608;
wire            n9609;
wire            n961;
wire            n9610;
wire            n9611;
wire            n9612;
wire            n9613;
wire            n9614;
wire            n9615;
wire            n9616;
wire            n9617;
wire            n9618;
wire            n9619;
wire            n962;
wire            n9620;
wire            n9621;
wire            n9622;
wire            n9623;
wire            n9624;
wire            n9625;
wire            n9626;
wire            n9627;
wire            n9628;
wire            n9629;
wire            n963;
wire            n9630;
wire            n9631;
wire            n9632;
wire            n9633;
wire            n9634;
wire            n9635;
wire            n9636;
wire            n9637;
wire            n9638;
wire            n9639;
wire            n964;
wire            n9640;
wire            n9641;
wire            n9642;
wire            n9643;
wire            n9644;
wire            n9645;
wire            n9646;
wire            n9647;
wire            n9648;
wire            n9649;
wire            n965;
wire            n9650;
wire            n9651;
wire            n9652;
wire            n9653;
wire            n9654;
wire            n9655;
wire            n9656;
wire            n9657;
wire            n9658;
wire            n9659;
wire            n966;
wire            n9660;
wire            n9661;
wire            n9662;
wire            n9663;
wire            n9664;
wire            n9665;
wire            n9666;
wire            n9667;
wire            n9668;
wire            n9669;
wire            n967;
wire            n9670;
wire            n9671;
wire            n9672;
wire            n9673;
wire            n9674;
wire            n9675;
wire            n9676;
wire            n9677;
wire            n9678;
wire            n9679;
wire            n968;
wire            n9680;
wire            n9681;
wire            n9682;
wire            n9683;
wire            n9684;
wire            n9685;
wire            n9686;
wire            n9687;
wire            n9688;
wire            n9689;
wire            n969;
wire            n9690;
wire            n9691;
wire            n9692;
wire            n9693;
wire            n9694;
wire            n9695;
wire            n9696;
wire            n9697;
wire            n9698;
wire            n9699;
wire            n97;
wire            n970;
wire            n9700;
wire            n9701;
wire            n9702;
wire            n9703;
wire            n9704;
wire            n9705;
wire            n9706;
wire            n9707;
wire            n9708;
wire            n9709;
wire            n971;
wire            n9710;
wire            n9711;
wire            n9712;
wire            n9713;
wire            n9714;
wire            n9715;
wire            n9716;
wire            n9717;
wire            n9718;
wire            n9719;
wire            n972;
wire            n9720;
wire            n9721;
wire            n9722;
wire            n9723;
wire            n9724;
wire            n9725;
wire            n9726;
wire            n9727;
wire            n9728;
wire            n9729;
wire            n973;
wire            n9730;
wire            n9731;
wire            n9732;
wire            n9733;
wire            n9734;
wire            n9735;
wire            n9736;
wire            n9737;
wire            n9738;
wire            n9739;
wire            n974;
wire            n9740;
wire            n9741;
wire            n9742;
wire            n9743;
wire            n9744;
wire            n9745;
wire            n9746;
wire            n9747;
wire            n9748;
wire            n9749;
wire            n975;
wire            n9750;
wire            n9751;
wire            n9752;
wire            n9753;
wire            n9754;
wire            n9755;
wire            n9756;
wire            n9757;
wire            n9758;
wire            n9759;
wire            n976;
wire            n9760;
wire            n9761;
wire            n9762;
wire            n9763;
wire            n9764;
wire            n9765;
wire            n9766;
wire            n9767;
wire            n9768;
wire            n9769;
wire            n977;
wire            n9770;
wire            n9771;
wire            n9772;
wire            n9773;
wire            n9774;
wire            n9775;
wire            n9776;
wire            n9777;
wire            n9778;
wire            n9779;
wire            n978;
wire            n9780;
wire            n9781;
wire            n9782;
wire            n9783;
wire            n9784;
wire            n9785;
wire            n9786;
wire            n9787;
wire            n9788;
wire            n9789;
wire            n979;
wire            n9790;
wire            n9791;
wire            n9792;
wire            n9793;
wire            n9794;
wire            n9795;
wire            n9796;
wire            n9797;
wire            n9798;
wire            n9799;
wire            n98;
wire            n980;
wire            n9800;
wire            n9801;
wire            n9802;
wire            n9803;
wire            n9804;
wire            n9805;
wire            n9806;
wire            n9807;
wire            n9808;
wire            n9809;
wire            n981;
wire            n9810;
wire            n9811;
wire            n9812;
wire            n9813;
wire            n9814;
wire            n9815;
wire            n9816;
wire            n9817;
wire            n9818;
wire            n9819;
wire            n982;
wire            n9820;
wire            n9821;
wire            n9822;
wire            n9823;
wire            n9824;
wire            n9825;
wire            n9826;
wire            n9827;
wire            n9828;
wire            n9829;
wire            n983;
wire            n9830;
wire            n9831;
wire            n9832;
wire            n9833;
wire            n9834;
wire            n9835;
wire            n9836;
wire            n9837;
wire            n9838;
wire            n9839;
wire            n984;
wire            n9840;
wire            n9841;
wire            n9842;
wire            n9843;
wire            n9844;
wire            n9845;
wire            n9846;
wire            n9847;
wire            n9848;
wire            n9849;
wire            n985;
wire            n9850;
wire            n9851;
wire            n9852;
wire            n9853;
wire            n9854;
wire            n9855;
wire            n9856;
wire            n9857;
wire            n9858;
wire            n9859;
wire            n986;
wire            n9860;
wire            n9861;
wire            n9862;
wire            n9863;
wire            n9864;
wire            n9865;
wire            n9866;
wire            n9867;
wire            n9868;
wire            n9869;
wire            n987;
wire            n9870;
wire            n9871;
wire            n9872;
wire            n9873;
wire            n9874;
wire            n9875;
wire            n9876;
wire            n9877;
wire            n9878;
wire            n9879;
wire            n988;
wire            n9880;
wire            n9881;
wire            n9882;
wire            n9883;
wire            n9884;
wire            n9885;
wire            n9886;
wire            n9887;
wire            n9888;
wire            n9889;
wire            n989;
wire            n9890;
wire            n9891;
wire            n9892;
wire            n9893;
wire            n9894;
wire            n9895;
wire            n9896;
wire            n9897;
wire            n9898;
wire            n9899;
wire            n99;
wire            n990;
wire            n9900;
wire            n9901;
wire            n9902;
wire            n9903;
wire            n9904;
wire            n9905;
wire            n9906;
wire            n9907;
wire            n9908;
wire            n9909;
wire            n991;
wire            n9910;
wire            n9911;
wire            n9912;
wire            n9913;
wire            n9914;
wire            n9915;
wire            n9916;
wire            n9917;
wire            n9918;
wire            n9919;
wire            n992;
wire            n9920;
wire            n9921;
wire            n9922;
wire            n9923;
wire            n9924;
wire            n9925;
wire            n9926;
wire            n9927;
wire            n9928;
wire            n9929;
wire            n993;
wire            n9930;
wire            n9931;
wire            n9932;
wire            n9933;
wire            n9934;
wire            n9935;
wire            n9936;
wire            n9937;
wire            n9938;
wire            n9939;
wire            n994;
wire            n9940;
wire            n9941;
wire            n9942;
wire            n9943;
wire            n9944;
wire            n9945;
wire            n9946;
wire            n9947;
wire            n9948;
wire            n9949;
wire            n995;
wire            n9950;
wire            n9951;
wire            n9952;
wire            n9953;
wire            n9954;
wire            n9955;
wire            n9956;
wire            n9957;
wire            n9958;
wire            n9959;
wire            n996;
wire            n9960;
wire            n9961;
wire            n9962;
wire            n9963;
wire            n9964;
wire            n9965;
wire            n9966;
wire            n9967;
wire            n9968;
wire            n9969;
wire            n997;
wire            n9970;
wire            n9971;
wire            n9972;
wire            n9973;
wire            n9974;
wire            n9975;
wire            n9976;
wire            n9977;
wire            n9978;
wire            n9979;
wire            n998;
wire            n9980;
wire            n9981;
wire            n9982;
wire            n9983;
wire            n9984;
wire            n9985;
wire            n9986;
wire            n9987;
wire            n9988;
wire            n9989;
wire            n999;
wire            n9990;
wire            n9991;
wire            n9992;
wire            n9993;
wire            n9994;
wire            n9995;
wire            n9996;
wire            n9997;
wire            n9998;
wire            n9999;
wire            rst;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign n1 = ki[13:13] ;
assign bv_1_0_n2 = 1'h0 ;
assign n3 =  ( n1 ) == ( bv_1_0_n2 )  ;
assign n4 = ki[12:12] ;
assign bv_1_1_n5 = 1'h1 ;
assign n6 =  ( n4 ) == ( bv_1_1_n5 )  ;
assign n7 =  ( n3 ) | ( n6 )  ;
assign n8 = ki[11:11] ;
assign n9 =  ( n8 ) == ( bv_1_1_n5 )  ;
assign n10 =  ( n7 ) | ( n9 )  ;
assign n11 = ~ ( n10 )  ;
assign n12 = ki[13:13] ;
assign n13 =  ( n12 ) == ( bv_1_1_n5 )  ;
assign n14 = ki[12:12] ;
assign n15 =  ( n14 ) == ( bv_1_0_n2 )  ;
assign n16 =  ( n13 ) | ( n15 )  ;
assign n17 = ki[11:11] ;
assign n18 =  ( n17 ) == ( bv_1_0_n2 )  ;
assign n19 =  ( n16 ) | ( n18 )  ;
assign n20 = ~ ( n19 )  ;
assign n21 =  ( n11 ) | ( n20 )  ;
assign n22 = ki[13:13] ;
assign n23 =  ( n22 ) == ( bv_1_0_n2 )  ;
assign n24 = ki[12:12] ;
assign n25 =  ( n24 ) == ( bv_1_0_n2 )  ;
assign n26 =  ( n23 ) | ( n25 )  ;
assign n27 = ki[11:11] ;
assign n28 =  ( n27 ) == ( bv_1_0_n2 )  ;
assign n29 =  ( n26 ) | ( n28 )  ;
assign n30 = ~ ( n29 )  ;
assign n31 = ki[13:13] ;
assign n32 =  ( n31 ) == ( bv_1_1_n5 )  ;
assign n33 = ki[12:12] ;
assign n34 =  ( n33 ) == ( bv_1_1_n5 )  ;
assign n35 =  ( n32 ) | ( n34 )  ;
assign n36 = ki[11:11] ;
assign n37 =  ( n36 ) == ( bv_1_1_n5 )  ;
assign n38 =  ( n35 ) | ( n37 )  ;
assign n39 = ~ ( n38 )  ;
assign n40 =  ( n30 ) | ( n39 )  ;
assign n41 = ki[13:13] ;
assign n42 =  ( n41 ) == ( bv_1_0_n2 )  ;
assign n43 = ki[12:12] ;
assign n44 =  ( n43 ) == ( bv_1_0_n2 )  ;
assign n45 = ki[11:11] ;
assign n46 =  ( n45 ) == ( bv_1_0_n2 )  ;
assign n47 =  ( n44 ) | ( n46 )  ;
assign n48 = ~ ( n47 )  ;
assign n49 =  ( n42 ) | ( n48 )  ;
assign n50 = i_wb_data[14:14] ;
assign n51 = ~ ( n50 ) ;
assign n52 = sp[14:14] ;
assign n53 =  ( n51 ) ^ ( n52 )  ;
assign n54 = i_wb_data[13:13] ;
assign n55 = sp[13:13] ;
assign n56 = ~ ( n55 ) ;
assign n57 =  ( n54 ) | ( n56 )  ;
assign n58 = ~ ( n57 ) ;
assign n59 = i_wb_data[13:13] ;
assign n60 = ~ ( n59 ) ;
assign n61 = sp[13:13] ;
assign n62 =  ( n60 ) ^ ( n61 )  ;
assign n63 = ~ ( n62 ) ;
assign n64 = i_wb_data[12:12] ;
assign n65 = sp[12:12] ;
assign n66 = ~ ( n65 ) ;
assign n67 =  ( n64 ) | ( n66 )  ;
assign n68 = ~ ( n67 ) ;
assign n69 = i_wb_data[12:12] ;
assign n70 = ~ ( n69 ) ;
assign n71 = sp[12:12] ;
assign n72 =  ( n70 ) ^ ( n71 )  ;
assign n73 = ~ ( n72 ) ;
assign n74 = i_wb_data[11:11] ;
assign n75 =  ( n73 ) | ( n74 )  ;
assign n76 = sp[11:11] ;
assign n77 = ~ ( n76 ) ;
assign n78 =  ( n75 ) | ( n77 )  ;
assign n79 = ~ ( n78 ) ;
assign n80 =  ( n68 ) | ( n79 )  ;
assign n81 = i_wb_data[11:11] ;
assign n82 = ~ ( n81 ) ;
assign n83 = sp[11:11] ;
assign n84 =  ( n82 ) ^ ( n83 )  ;
assign n85 = ~ ( n84 ) ;
assign n86 =  ( n73 ) | ( n85 )  ;
assign n87 = i_wb_data[10:10] ;
assign n88 = sp[10:10] ;
assign n89 = ~ ( n88 ) ;
assign n90 =  ( n87 ) | ( n89 )  ;
assign n91 = ~ ( n90 ) ;
assign n92 = i_wb_data[10:10] ;
assign n93 = ~ ( n92 ) ;
assign n94 = sp[10:10] ;
assign n95 =  ( n93 ) ^ ( n94 )  ;
assign n96 = ~ ( n95 ) ;
assign n97 = i_wb_data[9:9] ;
assign n98 =  ( n96 ) | ( n97 )  ;
assign n99 = sp[9:9] ;
assign n100 = ~ ( n99 ) ;
assign n101 =  ( n98 ) | ( n100 )  ;
assign n102 = ~ ( n101 ) ;
assign n103 =  ( n91 ) | ( n102 )  ;
assign n104 = ~ ( n103 ) ;
assign n105 =  ( n86 ) | ( n104 )  ;
assign n106 = ~ ( n105 ) ;
assign n107 =  ( n80 ) | ( n106 )  ;
assign n108 =  ( n73 ) | ( n85 )  ;
assign n109 =  ( n108 ) | ( n96 )  ;
assign n110 = i_wb_data[9:9] ;
assign n111 = ~ ( n110 ) ;
assign n112 = sp[9:9] ;
assign n113 =  ( n111 ) ^ ( n112 )  ;
assign n114 = ~ ( n113 ) ;
assign n115 =  ( n109 ) | ( n114 )  ;
assign n116 = i_wb_data[8:8] ;
assign n117 = sp[8:8] ;
assign n118 = ~ ( n117 ) ;
assign n119 =  ( n116 ) | ( n118 )  ;
assign n120 = ~ ( n119 ) ;
assign n121 = i_wb_data[8:8] ;
assign n122 = ~ ( n121 ) ;
assign n123 = sp[8:8] ;
assign n124 =  ( n122 ) ^ ( n123 )  ;
assign n125 = ~ ( n124 ) ;
assign n126 = i_wb_data[7:7] ;
assign n127 =  ( n125 ) | ( n126 )  ;
assign n128 = sp[7:7] ;
assign n129 = ~ ( n128 ) ;
assign n130 =  ( n127 ) | ( n129 )  ;
assign n131 = ~ ( n130 ) ;
assign n132 =  ( n120 ) | ( n131 )  ;
assign n133 = i_wb_data[7:7] ;
assign n134 = ~ ( n133 ) ;
assign n135 = sp[7:7] ;
assign n136 =  ( n134 ) ^ ( n135 )  ;
assign n137 = ~ ( n136 ) ;
assign n138 =  ( n125 ) | ( n137 )  ;
assign n139 = i_wb_data[6:6] ;
assign n140 = sp[6:6] ;
assign n141 = ~ ( n140 ) ;
assign n142 =  ( n139 ) | ( n141 )  ;
assign n143 = ~ ( n142 ) ;
assign n144 = i_wb_data[6:6] ;
assign n145 = ~ ( n144 ) ;
assign n146 = sp[6:6] ;
assign n147 =  ( n145 ) ^ ( n146 )  ;
assign n148 = ~ ( n147 ) ;
assign n149 = i_wb_data[5:5] ;
assign n150 =  ( n148 ) | ( n149 )  ;
assign n151 = sp[5:5] ;
assign n152 = ~ ( n151 ) ;
assign n153 =  ( n150 ) | ( n152 )  ;
assign n154 = ~ ( n153 ) ;
assign n155 =  ( n143 ) | ( n154 )  ;
assign n156 = ~ ( n155 ) ;
assign n157 =  ( n138 ) | ( n156 )  ;
assign n158 = ~ ( n157 ) ;
assign n159 =  ( n132 ) | ( n158 )  ;
assign n160 = ~ ( n159 ) ;
assign n161 =  ( n115 ) | ( n160 )  ;
assign n162 = ~ ( n161 ) ;
assign n163 =  ( n107 ) | ( n162 )  ;
assign n164 =  ( n73 ) | ( n85 )  ;
assign n165 =  ( n164 ) | ( n96 )  ;
assign n166 =  ( n165 ) | ( n114 )  ;
assign n167 =  ( n166 ) | ( n125 )  ;
assign n168 =  ( n167 ) | ( n137 )  ;
assign n169 =  ( n168 ) | ( n148 )  ;
assign n170 = i_wb_data[5:5] ;
assign n171 = ~ ( n170 ) ;
assign n172 = sp[5:5] ;
assign n173 =  ( n171 ) ^ ( n172 )  ;
assign n174 = ~ ( n173 ) ;
assign n175 =  ( n169 ) | ( n174 )  ;
assign n176 = i_wb_data[4:4] ;
assign n177 = sp[4:4] ;
assign n178 = ~ ( n177 ) ;
assign n179 =  ( n176 ) | ( n178 )  ;
assign n180 = ~ ( n179 ) ;
assign n181 = i_wb_data[4:4] ;
assign n182 = ~ ( n181 ) ;
assign n183 = sp[4:4] ;
assign n184 =  ( n182 ) ^ ( n183 )  ;
assign n185 = ~ ( n184 ) ;
assign n186 = i_wb_data[3:3] ;
assign n187 =  ( n185 ) | ( n186 )  ;
assign n188 = sp[3:3] ;
assign n189 = ~ ( n188 ) ;
assign n190 =  ( n187 ) | ( n189 )  ;
assign n191 = ~ ( n190 ) ;
assign n192 =  ( n180 ) | ( n191 )  ;
assign n193 = i_wb_data[3:3] ;
assign n194 = ~ ( n193 ) ;
assign n195 = sp[3:3] ;
assign n196 =  ( n194 ) ^ ( n195 )  ;
assign n197 = ~ ( n196 ) ;
assign n198 =  ( n185 ) | ( n197 )  ;
assign n199 = i_wb_data[2:2] ;
assign n200 = sp[2:2] ;
assign n201 = ~ ( n200 ) ;
assign n202 =  ( n199 ) | ( n201 )  ;
assign n203 = ~ ( n202 ) ;
assign n204 = i_wb_data[2:2] ;
assign n205 = ~ ( n204 ) ;
assign n206 = sp[2:2] ;
assign n207 =  ( n205 ) ^ ( n206 )  ;
assign n208 = ~ ( n207 ) ;
assign n209 = i_wb_data[1:1] ;
assign n210 =  ( n208 ) | ( n209 )  ;
assign n211 = sp[1:1] ;
assign n212 = ~ ( n211 ) ;
assign n213 =  ( n210 ) | ( n212 )  ;
assign n214 = ~ ( n213 ) ;
assign n215 =  ( n203 ) | ( n214 )  ;
assign n216 = ~ ( n215 ) ;
assign n217 =  ( n198 ) | ( n216 )  ;
assign n218 = ~ ( n217 ) ;
assign n219 =  ( n192 ) | ( n218 )  ;
assign n220 =  ( n185 ) | ( n197 )  ;
assign n221 =  ( n220 ) | ( n208 )  ;
assign n222 = i_wb_data[1:1] ;
assign n223 = ~ ( n222 ) ;
assign n224 = sp[1:1] ;
assign n225 =  ( n223 ) ^ ( n224 )  ;
assign n226 = ~ ( n225 ) ;
assign n227 =  ( n221 ) | ( n226 )  ;
assign n228 = i_wb_data[0:0] ;
assign n229 = sp[0:0] ;
assign n230 = ~ ( n229 ) ;
assign n231 =  ( n228 ) | ( n230 )  ;
assign n232 = ~ ( n231 ) ;
assign n233 = i_wb_data[0:0] ;
assign n234 = ~ ( n233 ) ;
assign n235 = sp[0:0] ;
assign n236 =  ( n234 ) ^ ( n235 )  ;
assign n237 =  ( n232 ) | ( n236 )  ;
assign n238 = ~ ( n237 ) ;
assign n239 =  ( n227 ) | ( n238 )  ;
assign n240 = ~ ( n239 ) ;
assign n241 =  ( n219 ) | ( n240 )  ;
assign n242 = ~ ( n241 ) ;
assign n243 =  ( n175 ) | ( n242 )  ;
assign n244 = ~ ( n243 ) ;
assign n245 =  ( n163 ) | ( n244 )  ;
assign n246 = ~ ( n245 ) ;
assign n247 =  ( n63 ) | ( n246 )  ;
assign n248 = ~ ( n247 ) ;
assign n249 =  ( n58 ) | ( n248 )  ;
assign n250 =  ( n53 ) ^ ( n249 )  ;
assign n251 = i_wb_data[14:14] ;
assign n252 = ~ ( n251 ) ;
assign n253 = sp[14:14] ;
assign n254 =  ( n252 ) ^ ( n253 )  ;
assign n255 =  ( n254 ) ^ ( n249 )  ;
assign n256 = ~ ( n255 ) ;
assign n257 =  ( n49 ) ? ( n250 ) : ( n256 ) ;
assign n258 =  ( n40 ) ? ( bv_1_0_n2 ) : ( n257 ) ;
assign n259 =  ( n30 ) | ( n39 )  ;
assign n260 = ki[13:13] ;
assign n261 =  ( n260 ) == ( bv_1_0_n2 )  ;
assign n262 =  ( n261 ) | ( n48 )  ;
assign n263 = i_wb_data[15:15] ;
assign n264 = ~ ( n263 ) ;
assign n265 = sp[15:15] ;
assign n266 =  ( n264 ) ^ ( n265 )  ;
assign n267 = i_wb_data[14:14] ;
assign n268 = sp[14:14] ;
assign n269 = ~ ( n268 ) ;
assign n270 =  ( n267 ) | ( n269 )  ;
assign n271 = ~ ( n270 ) ;
assign n272 = i_wb_data[14:14] ;
assign n273 = ~ ( n272 ) ;
assign n274 = sp[14:14] ;
assign n275 =  ( n273 ) ^ ( n274 )  ;
assign n276 = ~ ( n275 ) ;
assign n277 = i_wb_data[13:13] ;
assign n278 =  ( n276 ) | ( n277 )  ;
assign n279 = sp[13:13] ;
assign n280 = ~ ( n279 ) ;
assign n281 =  ( n278 ) | ( n280 )  ;
assign n282 = ~ ( n281 ) ;
assign n283 =  ( n271 ) | ( n282 )  ;
assign n284 =  ( n276 ) | ( n63 )  ;
assign n285 =  ( n68 ) | ( n79 )  ;
assign n286 = ~ ( n285 ) ;
assign n287 =  ( n284 ) | ( n286 )  ;
assign n288 = ~ ( n287 ) ;
assign n289 =  ( n283 ) | ( n288 )  ;
assign n290 =  ( n276 ) | ( n63 )  ;
assign n291 =  ( n290 ) | ( n73 )  ;
assign n292 =  ( n291 ) | ( n85 )  ;
assign n293 =  ( n91 ) | ( n102 )  ;
assign n294 =  ( n96 ) | ( n114 )  ;
assign n295 =  ( n120 ) | ( n131 )  ;
assign n296 = ~ ( n295 ) ;
assign n297 =  ( n294 ) | ( n296 )  ;
assign n298 = ~ ( n297 ) ;
assign n299 =  ( n293 ) | ( n298 )  ;
assign n300 = ~ ( n299 ) ;
assign n301 =  ( n292 ) | ( n300 )  ;
assign n302 = ~ ( n301 ) ;
assign n303 =  ( n289 ) | ( n302 )  ;
assign n304 =  ( n276 ) | ( n63 )  ;
assign n305 =  ( n304 ) | ( n73 )  ;
assign n306 =  ( n305 ) | ( n85 )  ;
assign n307 =  ( n306 ) | ( n96 )  ;
assign n308 =  ( n307 ) | ( n114 )  ;
assign n309 =  ( n308 ) | ( n125 )  ;
assign n310 =  ( n309 ) | ( n137 )  ;
assign n311 =  ( n143 ) | ( n154 )  ;
assign n312 =  ( n148 ) | ( n174 )  ;
assign n313 =  ( n180 ) | ( n191 )  ;
assign n314 = ~ ( n313 ) ;
assign n315 =  ( n312 ) | ( n314 )  ;
assign n316 = ~ ( n315 ) ;
assign n317 =  ( n311 ) | ( n316 )  ;
assign n318 =  ( n148 ) | ( n174 )  ;
assign n319 =  ( n318 ) | ( n185 )  ;
assign n320 =  ( n319 ) | ( n197 )  ;
assign n321 =  ( n203 ) | ( n214 )  ;
assign n322 =  ( n208 ) | ( n226 )  ;
assign n323 = ~ ( n237 ) ;
assign n324 =  ( n322 ) | ( n323 )  ;
assign n325 = ~ ( n324 ) ;
assign n326 =  ( n321 ) | ( n325 )  ;
assign n327 = ~ ( n326 ) ;
assign n328 =  ( n320 ) | ( n327 )  ;
assign n329 = ~ ( n328 ) ;
assign n330 =  ( n317 ) | ( n329 )  ;
assign n331 = ~ ( n330 ) ;
assign n332 =  ( n310 ) | ( n331 )  ;
assign n333 = ~ ( n332 ) ;
assign n334 =  ( n303 ) | ( n333 )  ;
assign n335 =  ( n266 ) ^ ( n334 )  ;
assign n336 = i_wb_data[15:15] ;
assign n337 = ~ ( n336 ) ;
assign n338 = sp[15:15] ;
assign n339 =  ( n337 ) ^ ( n338 )  ;
assign n340 =  ( n339 ) ^ ( n334 )  ;
assign n341 = ~ ( n340 ) ;
assign n342 =  ( n262 ) ? ( n335 ) : ( n341 ) ;
assign n343 =  ( n259 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n344 =  ( n21 ) ? ( n258 ) : ( n343 ) ;
assign n345 = ~ ( n344 ) ;
assign n346 = ki[14:14] ;
assign n347 =  ( n346 ) == ( bv_1_1_n5 )  ;
assign n348 = ki[13:13] ;
assign n349 =  ( n348 ) == ( bv_1_1_n5 )  ;
assign n350 =  ( n347 ) | ( n349 )  ;
assign n351 = ki[15:15] ;
assign n352 =  ( n351 ) == ( bv_1_0_n2 )  ;
assign n353 =  ( n350 ) | ( n352 )  ;
assign n354 = ~ ( n353 )  ;
assign n355 = ki[15:15] ;
assign n356 =  ( n355 ) == ( bv_1_1_n5 )  ;
assign n357 = ki[14:14] ;
assign n358 =  ( n357 ) == ( bv_1_0_n2 )  ;
assign n359 =  ( n356 ) | ( n358 )  ;
assign n360 = ki[13:13] ;
assign n361 =  ( n360 ) == ( bv_1_0_n2 )  ;
assign n362 =  ( n359 ) | ( n361 )  ;
assign n363 = ~ ( n362 )  ;
assign n364 =  ( n354 ) | ( n363 )  ;
assign n365 = ki[15:15] ;
assign n366 =  ( n365 ) == ( bv_1_0_n2 )  ;
assign n367 = ki[14:14] ;
assign n368 =  ( n367 ) == ( bv_1_0_n2 )  ;
assign n369 =  ( n366 ) | ( n368 )  ;
assign n370 = ki[13:13] ;
assign n371 =  ( n370 ) == ( bv_1_0_n2 )  ;
assign n372 =  ( n369 ) | ( n371 )  ;
assign n373 = ~ ( n372 )  ;
assign n374 = ki[14:14] ;
assign n375 =  ( n374 ) == ( bv_1_1_n5 )  ;
assign n376 = ki[13:13] ;
assign n377 =  ( n376 ) == ( bv_1_1_n5 )  ;
assign n378 =  ( n375 ) | ( n377 )  ;
assign n379 = ki[15:15] ;
assign n380 =  ( n379 ) == ( bv_1_1_n5 )  ;
assign n381 =  ( n378 ) | ( n380 )  ;
assign n382 = ~ ( n381 )  ;
assign n383 =  ( n373 ) | ( n382 )  ;
assign n384 = ki[15:15] ;
assign n385 =  ( n384 ) == ( bv_1_0_n2 )  ;
assign n386 = ki[14:14] ;
assign n387 =  ( n386 ) == ( bv_1_0_n2 )  ;
assign n388 = ki[13:13] ;
assign n389 =  ( n388 ) == ( bv_1_0_n2 )  ;
assign n390 =  ( n387 ) | ( n389 )  ;
assign n391 = ~ ( n390 )  ;
assign n392 =  ( n385 ) | ( n391 )  ;
assign n393 = i_wb_data[12:12] ;
assign n394 = ~ ( n393 ) ;
assign n395 = sp[12:12] ;
assign n396 =  ( n394 ) ^ ( n395 )  ;
assign n397 = i_wb_data[11:11] ;
assign n398 = sp[11:11] ;
assign n399 = ~ ( n398 ) ;
assign n400 =  ( n397 ) | ( n399 )  ;
assign n401 = ~ ( n400 ) ;
assign n402 =  ( n91 ) | ( n102 )  ;
assign n403 =  ( n402 ) | ( n298 )  ;
assign n404 =  ( n96 ) | ( n114 )  ;
assign n405 =  ( n404 ) | ( n125 )  ;
assign n406 =  ( n405 ) | ( n137 )  ;
assign n407 =  ( n143 ) | ( n154 )  ;
assign n408 =  ( n407 ) | ( n316 )  ;
assign n409 = ~ ( n408 ) ;
assign n410 =  ( n406 ) | ( n409 )  ;
assign n411 = ~ ( n410 ) ;
assign n412 =  ( n403 ) | ( n411 )  ;
assign n413 =  ( n96 ) | ( n114 )  ;
assign n414 =  ( n413 ) | ( n125 )  ;
assign n415 =  ( n414 ) | ( n137 )  ;
assign n416 =  ( n415 ) | ( n148 )  ;
assign n417 =  ( n416 ) | ( n174 )  ;
assign n418 =  ( n417 ) | ( n185 )  ;
assign n419 =  ( n418 ) | ( n197 )  ;
assign n420 = ~ ( n326 ) ;
assign n421 =  ( n419 ) | ( n420 )  ;
assign n422 = ~ ( n421 ) ;
assign n423 =  ( n412 ) | ( n422 )  ;
assign n424 = ~ ( n423 ) ;
assign n425 =  ( n85 ) | ( n424 )  ;
assign n426 = ~ ( n425 ) ;
assign n427 =  ( n401 ) | ( n426 )  ;
assign n428 =  ( n396 ) ^ ( n427 )  ;
assign n429 = i_wb_data[12:12] ;
assign n430 = ~ ( n429 ) ;
assign n431 = sp[12:12] ;
assign n432 =  ( n430 ) ^ ( n431 )  ;
assign n433 =  ( n432 ) ^ ( n427 )  ;
assign n434 = ~ ( n433 ) ;
assign n435 =  ( n392 ) ? ( n428 ) : ( n434 ) ;
assign n436 =  ( n383 ) ? ( bv_1_0_n2 ) : ( n435 ) ;
assign n437 =  ( n373 ) | ( n382 )  ;
assign n438 = ki[15:15] ;
assign n439 =  ( n438 ) == ( bv_1_0_n2 )  ;
assign n440 =  ( n439 ) | ( n391 )  ;
assign n441 = i_wb_data[13:13] ;
assign n442 = ~ ( n441 ) ;
assign n443 = sp[13:13] ;
assign n444 =  ( n442 ) ^ ( n443 )  ;
assign n445 =  ( n444 ) ^ ( n245 )  ;
assign n446 = i_wb_data[13:13] ;
assign n447 = ~ ( n446 ) ;
assign n448 = sp[13:13] ;
assign n449 =  ( n447 ) ^ ( n448 )  ;
assign n450 =  ( n449 ) ^ ( n245 )  ;
assign n451 = ~ ( n450 ) ;
assign n452 =  ( n440 ) ? ( n445 ) : ( n451 ) ;
assign n453 =  ( n437 ) ? ( bv_1_0_n2 ) : ( n452 ) ;
assign n454 =  ( n364 ) ? ( n436 ) : ( n453 ) ;
assign n455 = ~ ( n454 ) ;
assign n456 =  ( n345 ) | ( n455 )  ;
assign n457 = ~ ( n456 ) ;
assign n458 =  ( n344 ) ^ ( n454 )  ;
assign n459 =  ( n457 ) | ( n458 )  ;
assign n460 = ~ ( n459 ) ;
assign n461 =  ( n30 ) | ( n39 )  ;
assign n462 =  ( n461 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n463 =  ( n460 ) | ( n462 )  ;
assign n464 = ~ ( n463 ) ;
assign n465 =  ( n30 ) | ( n39 )  ;
assign n466 =  ( n465 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n467 = ~ ( n466 ) ;
assign n468 =  ( n459 ) ^ ( n467 )  ;
assign n469 = ~ ( n468 ) ;
assign n470 =  ( n354 ) | ( n363 )  ;
assign n471 =  ( n373 ) | ( n382 )  ;
assign n472 =  ( n471 ) ? ( bv_1_0_n2 ) : ( n452 ) ;
assign n473 =  ( n373 ) | ( n382 )  ;
assign n474 = ki[15:15] ;
assign n475 =  ( n474 ) == ( bv_1_0_n2 )  ;
assign n476 =  ( n475 ) | ( n391 )  ;
assign n477 = i_wb_data[14:14] ;
assign n478 = ~ ( n477 ) ;
assign n479 = sp[14:14] ;
assign n480 =  ( n478 ) ^ ( n479 )  ;
assign n481 =  ( n480 ) ^ ( n249 )  ;
assign n482 =  ( n476 ) ? ( n481 ) : ( n256 ) ;
assign n483 =  ( n473 ) ? ( bv_1_0_n2 ) : ( n482 ) ;
assign n484 =  ( n470 ) ? ( n472 ) : ( n483 ) ;
assign n485 = ~ ( n484 ) ;
assign n486 =  ( n469 ) | ( n485 )  ;
assign n487 = ~ ( n486 ) ;
assign n488 =  ( n464 ) | ( n487 )  ;
assign n489 = ~ ( n488 ) ;
assign n490 =  ( n354 ) | ( n363 )  ;
assign n491 =  ( n373 ) | ( n382 )  ;
assign n492 =  ( n491 ) ? ( bv_1_0_n2 ) : ( n482 ) ;
assign n493 =  ( n373 ) | ( n382 )  ;
assign n494 = ki[15:15] ;
assign n495 =  ( n494 ) == ( bv_1_0_n2 )  ;
assign n496 =  ( n495 ) | ( n391 )  ;
assign n497 = i_wb_data[15:15] ;
assign n498 = ~ ( n497 ) ;
assign n499 = sp[15:15] ;
assign n500 =  ( n498 ) ^ ( n499 )  ;
assign n501 =  ( n500 ) ^ ( n334 )  ;
assign n502 =  ( n496 ) ? ( n501 ) : ( n341 ) ;
assign n503 =  ( n493 ) ? ( bv_1_0_n2 ) : ( n502 ) ;
assign n504 =  ( n490 ) ? ( n492 ) : ( n503 ) ;
assign n505 = ~ ( n504 ) ;
assign n506 =  ( n489 ) | ( n505 )  ;
assign n507 = ~ ( n506 ) ;
assign n508 =  ( n488 ) ^ ( n504 )  ;
assign n509 =  ( n507 ) | ( n508 )  ;
assign n510 = ~ ( n509 ) ;
assign n511 =  ( n373 ) | ( n382 )  ;
assign n512 =  ( n511 ) ? ( bv_1_0_n2 ) : ( n502 ) ;
assign n513 =  ( n510 ) | ( n512 )  ;
assign n514 = ~ ( n513 ) ;
assign n515 =  ( n373 ) | ( n382 )  ;
assign n516 =  ( n515 ) ? ( bv_1_0_n2 ) : ( n502 ) ;
assign n517 = ~ ( n516 ) ;
assign n518 =  ( n509 ) ^ ( n517 )  ;
assign n519 = ~ ( n518 ) ;
assign n520 =  ( bv_1_1_n5 ) ^ ( n488 )  ;
assign n521 =  ( n520 ) ^ ( n504 )  ;
assign n522 = ~ ( n521 ) ;
assign n523 =  ( n519 ) | ( n522 )  ;
assign n524 = ki[9:9] ;
assign n525 =  ( n524 ) == ( bv_1_0_n2 )  ;
assign n526 = ki[8:8] ;
assign n527 =  ( n526 ) == ( bv_1_0_n2 )  ;
assign n528 =  ( n525 ) | ( n527 )  ;
assign n529 = ki[7:7] ;
assign n530 =  ( n529 ) == ( bv_1_0_n2 )  ;
assign n531 =  ( n528 ) | ( n530 )  ;
assign n532 = ~ ( n531 )  ;
assign n533 = ki[9:9] ;
assign n534 =  ( n533 ) == ( bv_1_1_n5 )  ;
assign n535 = ki[8:8] ;
assign n536 =  ( n535 ) == ( bv_1_1_n5 )  ;
assign n537 =  ( n534 ) | ( n536 )  ;
assign n538 = ki[7:7] ;
assign n539 =  ( n538 ) == ( bv_1_1_n5 )  ;
assign n540 =  ( n537 ) | ( n539 )  ;
assign n541 = ~ ( n540 )  ;
assign n542 =  ( n532 ) | ( n541 )  ;
assign n543 = ki[9:9] ;
assign n544 =  ( n543 ) == ( bv_1_0_n2 )  ;
assign n545 = ki[8:8] ;
assign n546 =  ( n545 ) == ( bv_1_0_n2 )  ;
assign n547 = ki[7:7] ;
assign n548 =  ( n547 ) == ( bv_1_0_n2 )  ;
assign n549 =  ( n546 ) | ( n548 )  ;
assign n550 = ~ ( n549 )  ;
assign n551 =  ( n544 ) | ( n550 )  ;
assign n552 = i_wb_data[15:15] ;
assign n553 = ~ ( n552 ) ;
assign n554 = sp[15:15] ;
assign n555 =  ( n553 ) ^ ( n554 )  ;
assign n556 =  ( n555 ) ^ ( n334 )  ;
assign n557 =  ( n551 ) ? ( n556 ) : ( n341 ) ;
assign n558 =  ( n542 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n559 = ki[11:11] ;
assign n560 =  ( n559 ) == ( bv_1_0_n2 )  ;
assign n561 = ki[10:10] ;
assign n562 =  ( n561 ) == ( bv_1_1_n5 )  ;
assign n563 =  ( n560 ) | ( n562 )  ;
assign n564 = ki[9:9] ;
assign n565 =  ( n564 ) == ( bv_1_1_n5 )  ;
assign n566 =  ( n563 ) | ( n565 )  ;
assign n567 = ~ ( n566 )  ;
assign n568 = ki[11:11] ;
assign n569 =  ( n568 ) == ( bv_1_1_n5 )  ;
assign n570 = ki[10:10] ;
assign n571 =  ( n570 ) == ( bv_1_0_n2 )  ;
assign n572 =  ( n569 ) | ( n571 )  ;
assign n573 = ki[9:9] ;
assign n574 =  ( n573 ) == ( bv_1_0_n2 )  ;
assign n575 =  ( n572 ) | ( n574 )  ;
assign n576 = ~ ( n575 )  ;
assign n577 =  ( n567 ) | ( n576 )  ;
assign n578 = ki[11:11] ;
assign n579 =  ( n578 ) == ( bv_1_0_n2 )  ;
assign n580 = ki[10:10] ;
assign n581 =  ( n580 ) == ( bv_1_0_n2 )  ;
assign n582 =  ( n579 ) | ( n581 )  ;
assign n583 = ki[9:9] ;
assign n584 =  ( n583 ) == ( bv_1_0_n2 )  ;
assign n585 =  ( n582 ) | ( n584 )  ;
assign n586 = ~ ( n585 )  ;
assign n587 = ki[11:11] ;
assign n588 =  ( n587 ) == ( bv_1_1_n5 )  ;
assign n589 = ki[10:10] ;
assign n590 =  ( n589 ) == ( bv_1_1_n5 )  ;
assign n591 =  ( n588 ) | ( n590 )  ;
assign n592 = ki[9:9] ;
assign n593 =  ( n592 ) == ( bv_1_1_n5 )  ;
assign n594 =  ( n591 ) | ( n593 )  ;
assign n595 = ~ ( n594 )  ;
assign n596 =  ( n586 ) | ( n595 )  ;
assign n597 = ki[11:11] ;
assign n598 =  ( n597 ) == ( bv_1_0_n2 )  ;
assign n599 = ki[10:10] ;
assign n600 =  ( n599 ) == ( bv_1_0_n2 )  ;
assign n601 = ki[9:9] ;
assign n602 =  ( n601 ) == ( bv_1_0_n2 )  ;
assign n603 =  ( n600 ) | ( n602 )  ;
assign n604 = ~ ( n603 )  ;
assign n605 =  ( n598 ) | ( n604 )  ;
assign n606 = i_wb_data[13:13] ;
assign n607 = ~ ( n606 ) ;
assign n608 = sp[13:13] ;
assign n609 =  ( n607 ) ^ ( n608 )  ;
assign n610 =  ( n609 ) ^ ( n245 )  ;
assign n611 =  ( n605 ) ? ( n610 ) : ( n451 ) ;
assign n612 =  ( n596 ) ? ( bv_1_0_n2 ) : ( n611 ) ;
assign n613 =  ( n586 ) | ( n595 )  ;
assign n614 = ki[11:11] ;
assign n615 =  ( n614 ) == ( bv_1_0_n2 )  ;
assign n616 =  ( n615 ) | ( n604 )  ;
assign n617 = i_wb_data[14:14] ;
assign n618 = ~ ( n617 ) ;
assign n619 = sp[14:14] ;
assign n620 =  ( n618 ) ^ ( n619 )  ;
assign n621 =  ( n620 ) ^ ( n249 )  ;
assign n622 =  ( n616 ) ? ( n621 ) : ( n256 ) ;
assign n623 =  ( n613 ) ? ( bv_1_0_n2 ) : ( n622 ) ;
assign n624 =  ( n577 ) ? ( n612 ) : ( n623 ) ;
assign n625 = ~ ( n624 ) ;
assign n626 =  ( n558 ) | ( n625 )  ;
assign n627 = ~ ( n626 ) ;
assign n628 =  ( n532 ) | ( n541 )  ;
assign n629 =  ( n628 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n630 = ~ ( n629 ) ;
assign n631 =  ( n630 ) ^ ( n624 )  ;
assign n632 = ~ ( n631 ) ;
assign n633 =  ( n11 ) | ( n20 )  ;
assign n634 =  ( n30 ) | ( n39 )  ;
assign n635 = ki[13:13] ;
assign n636 =  ( n635 ) == ( bv_1_0_n2 )  ;
assign n637 =  ( n636 ) | ( n48 )  ;
assign n638 = i_wb_data[11:11] ;
assign n639 = ~ ( n638 ) ;
assign n640 = sp[11:11] ;
assign n641 =  ( n639 ) ^ ( n640 )  ;
assign n642 =  ( n641 ) ^ ( n423 )  ;
assign n643 = i_wb_data[11:11] ;
assign n644 = ~ ( n643 ) ;
assign n645 = sp[11:11] ;
assign n646 =  ( n644 ) ^ ( n645 )  ;
assign n647 =  ( n646 ) ^ ( n423 )  ;
assign n648 = ~ ( n647 ) ;
assign n649 =  ( n637 ) ? ( n642 ) : ( n648 ) ;
assign n650 =  ( n634 ) ? ( bv_1_0_n2 ) : ( n649 ) ;
assign n651 =  ( n30 ) | ( n39 )  ;
assign n652 = ki[13:13] ;
assign n653 =  ( n652 ) == ( bv_1_0_n2 )  ;
assign n654 =  ( n653 ) | ( n48 )  ;
assign n655 = i_wb_data[12:12] ;
assign n656 = ~ ( n655 ) ;
assign n657 = sp[12:12] ;
assign n658 =  ( n656 ) ^ ( n657 )  ;
assign n659 =  ( n658 ) ^ ( n427 )  ;
assign n660 =  ( n654 ) ? ( n659 ) : ( n434 ) ;
assign n661 =  ( n651 ) ? ( bv_1_0_n2 ) : ( n660 ) ;
assign n662 =  ( n633 ) ? ( n650 ) : ( n661 ) ;
assign n663 = ~ ( n662 ) ;
assign n664 =  ( n632 ) | ( n663 )  ;
assign n665 = ~ ( n664 ) ;
assign n666 =  ( n627 ) | ( n665 )  ;
assign n667 = ~ ( n666 ) ;
assign n668 =  ( n567 ) | ( n576 )  ;
assign n669 =  ( n586 ) | ( n595 )  ;
assign n670 =  ( n669 ) ? ( bv_1_0_n2 ) : ( n622 ) ;
assign n671 =  ( n586 ) | ( n595 )  ;
assign n672 = ki[11:11] ;
assign n673 =  ( n672 ) == ( bv_1_0_n2 )  ;
assign n674 =  ( n673 ) | ( n604 )  ;
assign n675 = i_wb_data[15:15] ;
assign n676 = ~ ( n675 ) ;
assign n677 = sp[15:15] ;
assign n678 =  ( n676 ) ^ ( n677 )  ;
assign n679 =  ( n678 ) ^ ( n334 )  ;
assign n680 =  ( n674 ) ? ( n679 ) : ( n341 ) ;
assign n681 =  ( n671 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n682 =  ( n668 ) ? ( n670 ) : ( n681 ) ;
assign n683 =  ( n11 ) | ( n20 )  ;
assign n684 =  ( n30 ) | ( n39 )  ;
assign n685 =  ( n684 ) ? ( bv_1_0_n2 ) : ( n660 ) ;
assign n686 =  ( n30 ) | ( n39 )  ;
assign n687 = ki[13:13] ;
assign n688 =  ( n687 ) == ( bv_1_0_n2 )  ;
assign n689 =  ( n688 ) | ( n48 )  ;
assign n690 = i_wb_data[13:13] ;
assign n691 = ~ ( n690 ) ;
assign n692 = sp[13:13] ;
assign n693 =  ( n691 ) ^ ( n692 )  ;
assign n694 =  ( n693 ) ^ ( n245 )  ;
assign n695 =  ( n689 ) ? ( n694 ) : ( n451 ) ;
assign n696 =  ( n686 ) ? ( bv_1_0_n2 ) : ( n695 ) ;
assign n697 =  ( n683 ) ? ( n685 ) : ( n696 ) ;
assign n698 =  ( n682 ) ^ ( n697 )  ;
assign n699 =  ( n354 ) | ( n363 )  ;
assign n700 =  ( n373 ) | ( n382 )  ;
assign n701 = ki[15:15] ;
assign n702 =  ( n701 ) == ( bv_1_0_n2 )  ;
assign n703 =  ( n702 ) | ( n391 )  ;
assign n704 = i_wb_data[10:10] ;
assign n705 = ~ ( n704 ) ;
assign n706 = sp[10:10] ;
assign n707 =  ( n705 ) ^ ( n706 )  ;
assign n708 = i_wb_data[9:9] ;
assign n709 = sp[9:9] ;
assign n710 = ~ ( n709 ) ;
assign n711 =  ( n708 ) | ( n710 )  ;
assign n712 = ~ ( n711 ) ;
assign n713 =  ( n120 ) | ( n131 )  ;
assign n714 =  ( n713 ) | ( n158 )  ;
assign n715 =  ( n125 ) | ( n137 )  ;
assign n716 =  ( n715 ) | ( n148 )  ;
assign n717 =  ( n716 ) | ( n174 )  ;
assign n718 =  ( n180 ) | ( n191 )  ;
assign n719 =  ( n718 ) | ( n218 )  ;
assign n720 = ~ ( n719 ) ;
assign n721 =  ( n717 ) | ( n720 )  ;
assign n722 = ~ ( n721 ) ;
assign n723 =  ( n714 ) | ( n722 )  ;
assign n724 =  ( n125 ) | ( n137 )  ;
assign n725 =  ( n724 ) | ( n148 )  ;
assign n726 =  ( n725 ) | ( n174 )  ;
assign n727 =  ( n726 ) | ( n185 )  ;
assign n728 =  ( n727 ) | ( n197 )  ;
assign n729 =  ( n728 ) | ( n208 )  ;
assign n730 =  ( n729 ) | ( n226 )  ;
assign n731 = ~ ( n237 ) ;
assign n732 =  ( n730 ) | ( n731 )  ;
assign n733 = ~ ( n732 ) ;
assign n734 =  ( n723 ) | ( n733 )  ;
assign n735 = ~ ( n734 ) ;
assign n736 =  ( n114 ) | ( n735 )  ;
assign n737 = ~ ( n736 ) ;
assign n738 =  ( n712 ) | ( n737 )  ;
assign n739 =  ( n707 ) ^ ( n738 )  ;
assign n740 = i_wb_data[10:10] ;
assign n741 = ~ ( n740 ) ;
assign n742 = sp[10:10] ;
assign n743 =  ( n741 ) ^ ( n742 )  ;
assign n744 =  ( n743 ) ^ ( n738 )  ;
assign n745 = ~ ( n744 ) ;
assign n746 =  ( n703 ) ? ( n739 ) : ( n745 ) ;
assign n747 =  ( n700 ) ? ( bv_1_0_n2 ) : ( n746 ) ;
assign n748 =  ( n373 ) | ( n382 )  ;
assign n749 = ki[15:15] ;
assign n750 =  ( n749 ) == ( bv_1_0_n2 )  ;
assign n751 =  ( n750 ) | ( n391 )  ;
assign n752 = i_wb_data[11:11] ;
assign n753 = ~ ( n752 ) ;
assign n754 = sp[11:11] ;
assign n755 =  ( n753 ) ^ ( n754 )  ;
assign n756 =  ( n755 ) ^ ( n423 )  ;
assign n757 =  ( n751 ) ? ( n756 ) : ( n648 ) ;
assign n758 =  ( n748 ) ? ( bv_1_0_n2 ) : ( n757 ) ;
assign n759 =  ( n699 ) ? ( n747 ) : ( n758 ) ;
assign n760 =  ( n698 ) ^ ( n759 )  ;
assign n761 = ~ ( n760 ) ;
assign n762 =  ( n667 ) | ( n761 )  ;
assign n763 = ~ ( n762 ) ;
assign n764 =  ( n666 ) ^ ( n682 )  ;
assign n765 =  ( n764 ) ^ ( n697 )  ;
assign n766 =  ( n765 ) ^ ( n759 )  ;
assign n767 =  ( n763 ) | ( n766 )  ;
assign n768 = ~ ( n767 ) ;
assign n769 = ~ ( n682 ) ;
assign n770 = ~ ( n697 ) ;
assign n771 =  ( n769 ) | ( n770 )  ;
assign n772 = ~ ( n771 ) ;
assign n773 =  ( n682 ) ^ ( n697 )  ;
assign n774 = ~ ( n773 ) ;
assign n775 = ~ ( n759 ) ;
assign n776 =  ( n774 ) | ( n775 )  ;
assign n777 = ~ ( n776 ) ;
assign n778 =  ( n772 ) | ( n777 )  ;
assign n779 = ~ ( n778 ) ;
assign n780 =  ( n768 ) | ( n779 )  ;
assign n781 = ~ ( n780 ) ;
assign n782 =  ( n666 ) ^ ( n682 )  ;
assign n783 =  ( n782 ) ^ ( n697 )  ;
assign n784 =  ( n783 ) ^ ( n759 )  ;
assign n785 =  ( n763 ) | ( n784 )  ;
assign n786 =  ( n785 ) ^ ( n778 )  ;
assign n787 = ~ ( n786 ) ;
assign n788 =  ( n586 ) | ( n595 )  ;
assign n789 =  ( n788 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n790 = ~ ( n789 ) ;
assign n791 =  ( n11 ) | ( n20 )  ;
assign n792 =  ( n30 ) | ( n39 )  ;
assign n793 =  ( n792 ) ? ( bv_1_0_n2 ) : ( n695 ) ;
assign n794 =  ( n30 ) | ( n39 )  ;
assign n795 =  ( n794 ) ? ( bv_1_0_n2 ) : ( n257 ) ;
assign n796 =  ( n791 ) ? ( n793 ) : ( n795 ) ;
assign n797 =  ( n790 ) ^ ( n796 )  ;
assign n798 =  ( n354 ) | ( n363 )  ;
assign n799 =  ( n373 ) | ( n382 )  ;
assign n800 =  ( n799 ) ? ( bv_1_0_n2 ) : ( n757 ) ;
assign n801 =  ( n373 ) | ( n382 )  ;
assign n802 =  ( n801 ) ? ( bv_1_0_n2 ) : ( n435 ) ;
assign n803 =  ( n798 ) ? ( n800 ) : ( n802 ) ;
assign n804 =  ( n797 ) ^ ( n803 )  ;
assign n805 = ~ ( n804 ) ;
assign n806 =  ( n787 ) | ( n805 )  ;
assign n807 = ~ ( n806 ) ;
assign n808 =  ( n781 ) | ( n807 )  ;
assign n809 = ~ ( n808 ) ;
assign n810 =  ( n586 ) | ( n595 )  ;
assign n811 =  ( n810 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n812 = ~ ( n796 ) ;
assign n813 =  ( n811 ) | ( n812 )  ;
assign n814 = ~ ( n813 ) ;
assign n815 =  ( n586 ) | ( n595 )  ;
assign n816 =  ( n815 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n817 = ~ ( n816 ) ;
assign n818 =  ( n817 ) ^ ( n796 )  ;
assign n819 = ~ ( n818 ) ;
assign n820 = ~ ( n803 ) ;
assign n821 =  ( n819 ) | ( n820 )  ;
assign n822 = ~ ( n821 ) ;
assign n823 =  ( n814 ) | ( n822 )  ;
assign n824 = ~ ( n823 ) ;
assign n825 =  ( n809 ) | ( n824 )  ;
assign n826 = ~ ( n825 ) ;
assign n827 =  ( n808 ) ^ ( n823 )  ;
assign n828 = ~ ( n827 ) ;
assign n829 =  ( bv_1_1_n5 ) ^ ( n344 )  ;
assign n830 =  ( n829 ) ^ ( n454 )  ;
assign n831 = ~ ( n830 ) ;
assign n832 =  ( n828 ) | ( n831 )  ;
assign n833 = ~ ( n832 ) ;
assign n834 =  ( n826 ) | ( n833 )  ;
assign n835 = ~ ( n834 ) ;
assign n836 =  ( n523 ) | ( n835 )  ;
assign n837 =  ( n30 ) | ( n39 )  ;
assign n838 =  ( n837 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n839 = ~ ( n838 ) ;
assign n840 =  ( n459 ) ^ ( n839 )  ;
assign n841 =  ( n840 ) ^ ( n484 )  ;
assign n842 = ~ ( n841 ) ;
assign n843 =  ( n836 ) | ( n842 )  ;
assign n844 = ~ ( n843 ) ;
assign n845 =  ( n514 ) | ( n844 )  ;
assign n846 = ~ ( n518 ) ;
assign n847 =  ( bv_1_1_n5 ) ^ ( n488 )  ;
assign n848 =  ( n847 ) ^ ( n504 )  ;
assign n849 = ~ ( n848 ) ;
assign n850 =  ( n846 ) | ( n849 )  ;
assign n851 =  ( n834 ) ^ ( n459 )  ;
assign n852 =  ( n30 ) | ( n39 )  ;
assign n853 =  ( n852 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n854 = ~ ( n853 ) ;
assign n855 =  ( n851 ) ^ ( n854 )  ;
assign n856 =  ( n855 ) ^ ( n484 )  ;
assign n857 = ~ ( n856 ) ;
assign n858 =  ( n850 ) | ( n857 )  ;
assign n859 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n860 =  ( n859 ) ^ ( n823 )  ;
assign n861 =  ( n860 ) ^ ( n344 )  ;
assign n862 =  ( n861 ) ^ ( n454 )  ;
assign n863 = ~ ( n862 ) ;
assign n864 =  ( n858 ) | ( n863 )  ;
assign n865 = ki[7:7] ;
assign n866 =  ( n865 ) == ( bv_1_0_n2 )  ;
assign n867 = ki[6:6] ;
assign n868 =  ( n867 ) == ( bv_1_0_n2 )  ;
assign n869 =  ( n866 ) | ( n868 )  ;
assign n870 = ki[5:5] ;
assign n871 =  ( n870 ) == ( bv_1_0_n2 )  ;
assign n872 =  ( n869 ) | ( n871 )  ;
assign n873 = ~ ( n872 )  ;
assign n874 = ki[7:7] ;
assign n875 =  ( n874 ) == ( bv_1_1_n5 )  ;
assign n876 = ki[6:6] ;
assign n877 =  ( n876 ) == ( bv_1_1_n5 )  ;
assign n878 =  ( n875 ) | ( n877 )  ;
assign n879 = ki[5:5] ;
assign n880 =  ( n879 ) == ( bv_1_1_n5 )  ;
assign n881 =  ( n878 ) | ( n880 )  ;
assign n882 = ~ ( n881 )  ;
assign n883 =  ( n873 ) | ( n882 )  ;
assign n884 = ki[7:7] ;
assign n885 =  ( n884 ) == ( bv_1_0_n2 )  ;
assign n886 = ki[6:6] ;
assign n887 =  ( n886 ) == ( bv_1_0_n2 )  ;
assign n888 = ki[5:5] ;
assign n889 =  ( n888 ) == ( bv_1_0_n2 )  ;
assign n890 =  ( n887 ) | ( n889 )  ;
assign n891 = ~ ( n890 )  ;
assign n892 =  ( n885 ) | ( n891 )  ;
assign n893 = i_wb_data[15:15] ;
assign n894 = ~ ( n893 ) ;
assign n895 = sp[15:15] ;
assign n896 =  ( n894 ) ^ ( n895 )  ;
assign n897 =  ( n896 ) ^ ( n334 )  ;
assign n898 =  ( n892 ) ? ( n897 ) : ( n341 ) ;
assign n899 =  ( n883 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n900 = ki[9:9] ;
assign n901 =  ( n900 ) == ( bv_1_0_n2 )  ;
assign n902 = ki[8:8] ;
assign n903 =  ( n902 ) == ( bv_1_1_n5 )  ;
assign n904 =  ( n901 ) | ( n903 )  ;
assign n905 = ki[7:7] ;
assign n906 =  ( n905 ) == ( bv_1_1_n5 )  ;
assign n907 =  ( n904 ) | ( n906 )  ;
assign n908 = ~ ( n907 )  ;
assign n909 = ki[9:9] ;
assign n910 =  ( n909 ) == ( bv_1_1_n5 )  ;
assign n911 = ki[8:8] ;
assign n912 =  ( n911 ) == ( bv_1_0_n2 )  ;
assign n913 =  ( n910 ) | ( n912 )  ;
assign n914 = ki[7:7] ;
assign n915 =  ( n914 ) == ( bv_1_0_n2 )  ;
assign n916 =  ( n913 ) | ( n915 )  ;
assign n917 = ~ ( n916 )  ;
assign n918 =  ( n908 ) | ( n917 )  ;
assign n919 =  ( n532 ) | ( n541 )  ;
assign n920 = ki[9:9] ;
assign n921 =  ( n920 ) == ( bv_1_0_n2 )  ;
assign n922 =  ( n921 ) | ( n550 )  ;
assign n923 = i_wb_data[13:13] ;
assign n924 = ~ ( n923 ) ;
assign n925 = sp[13:13] ;
assign n926 =  ( n924 ) ^ ( n925 )  ;
assign n927 =  ( n926 ) ^ ( n245 )  ;
assign n928 =  ( n922 ) ? ( n927 ) : ( n451 ) ;
assign n929 =  ( n919 ) ? ( bv_1_0_n2 ) : ( n928 ) ;
assign n930 =  ( n532 ) | ( n541 )  ;
assign n931 = ki[9:9] ;
assign n932 =  ( n931 ) == ( bv_1_0_n2 )  ;
assign n933 =  ( n932 ) | ( n550 )  ;
assign n934 = i_wb_data[14:14] ;
assign n935 = ~ ( n934 ) ;
assign n936 = sp[14:14] ;
assign n937 =  ( n935 ) ^ ( n936 )  ;
assign n938 =  ( n937 ) ^ ( n249 )  ;
assign n939 =  ( n933 ) ? ( n938 ) : ( n256 ) ;
assign n940 =  ( n930 ) ? ( bv_1_0_n2 ) : ( n939 ) ;
assign n941 =  ( n918 ) ? ( n929 ) : ( n940 ) ;
assign n942 = ~ ( n941 ) ;
assign n943 =  ( n899 ) | ( n942 )  ;
assign n944 =  ( n567 ) | ( n576 )  ;
assign n945 =  ( n586 ) | ( n595 )  ;
assign n946 = ki[11:11] ;
assign n947 =  ( n946 ) == ( bv_1_0_n2 )  ;
assign n948 =  ( n947 ) | ( n604 )  ;
assign n949 = i_wb_data[11:11] ;
assign n950 = ~ ( n949 ) ;
assign n951 = sp[11:11] ;
assign n952 =  ( n950 ) ^ ( n951 )  ;
assign n953 =  ( n952 ) ^ ( n423 )  ;
assign n954 =  ( n948 ) ? ( n953 ) : ( n648 ) ;
assign n955 =  ( n945 ) ? ( bv_1_0_n2 ) : ( n954 ) ;
assign n956 =  ( n586 ) | ( n595 )  ;
assign n957 = ki[11:11] ;
assign n958 =  ( n957 ) == ( bv_1_0_n2 )  ;
assign n959 =  ( n958 ) | ( n604 )  ;
assign n960 = i_wb_data[12:12] ;
assign n961 = ~ ( n960 ) ;
assign n962 = sp[12:12] ;
assign n963 =  ( n961 ) ^ ( n962 )  ;
assign n964 =  ( n963 ) ^ ( n427 )  ;
assign n965 =  ( n959 ) ? ( n964 ) : ( n434 ) ;
assign n966 =  ( n956 ) ? ( bv_1_0_n2 ) : ( n965 ) ;
assign n967 =  ( n944 ) ? ( n955 ) : ( n966 ) ;
assign n968 = ~ ( n967 ) ;
assign n969 =  ( n943 ) | ( n968 )  ;
assign n970 =  ( n11 ) | ( n20 )  ;
assign n971 =  ( n30 ) | ( n39 )  ;
assign n972 = ki[13:13] ;
assign n973 =  ( n972 ) == ( bv_1_0_n2 )  ;
assign n974 =  ( n973 ) | ( n48 )  ;
assign n975 = i_wb_data[9:9] ;
assign n976 = ~ ( n975 ) ;
assign n977 = sp[9:9] ;
assign n978 =  ( n976 ) ^ ( n977 )  ;
assign n979 =  ( n978 ) ^ ( n734 )  ;
assign n980 = i_wb_data[9:9] ;
assign n981 = ~ ( n980 ) ;
assign n982 = sp[9:9] ;
assign n983 =  ( n981 ) ^ ( n982 )  ;
assign n984 =  ( n983 ) ^ ( n734 )  ;
assign n985 = ~ ( n984 ) ;
assign n986 =  ( n974 ) ? ( n979 ) : ( n985 ) ;
assign n987 =  ( n971 ) ? ( bv_1_0_n2 ) : ( n986 ) ;
assign n988 =  ( n30 ) | ( n39 )  ;
assign n989 = ki[13:13] ;
assign n990 =  ( n989 ) == ( bv_1_0_n2 )  ;
assign n991 =  ( n990 ) | ( n48 )  ;
assign n992 = i_wb_data[10:10] ;
assign n993 = ~ ( n992 ) ;
assign n994 = sp[10:10] ;
assign n995 =  ( n993 ) ^ ( n994 )  ;
assign n996 =  ( n995 ) ^ ( n738 )  ;
assign n997 =  ( n991 ) ? ( n996 ) : ( n745 ) ;
assign n998 =  ( n988 ) ? ( bv_1_0_n2 ) : ( n997 ) ;
assign n999 =  ( n970 ) ? ( n987 ) : ( n998 ) ;
assign n1000 = ~ ( n999 ) ;
assign n1001 =  ( n969 ) | ( n1000 )  ;
assign n1002 = ~ ( n1001 ) ;
assign n1003 =  ( n873 ) | ( n882 )  ;
assign n1004 =  ( n1003 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n1005 = ~ ( n1004 ) ;
assign n1006 =  ( n1005 ) ^ ( n941 )  ;
assign n1007 = ~ ( n1006 ) ;
assign n1008 =  ( n967 ) ^ ( n999 )  ;
assign n1009 = ~ ( n1008 ) ;
assign n1010 =  ( n1007 ) | ( n1009 )  ;
assign n1011 = ~ ( n1010 ) ;
assign n1012 =  ( n1002 ) | ( n1011 )  ;
assign n1013 =  ( n873 ) | ( n882 )  ;
assign n1014 =  ( n1013 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n1015 = ~ ( n1014 ) ;
assign n1016 =  ( n1015 ) ^ ( n941 )  ;
assign n1017 =  ( n1016 ) ^ ( n967 )  ;
assign n1018 =  ( n1017 ) ^ ( n999 )  ;
assign n1019 = ~ ( n1018 ) ;
assign n1020 =  ( n354 ) | ( n363 )  ;
assign n1021 =  ( n373 ) | ( n382 )  ;
assign n1022 = ki[15:15] ;
assign n1023 =  ( n1022 ) == ( bv_1_0_n2 )  ;
assign n1024 =  ( n1023 ) | ( n391 )  ;
assign n1025 = i_wb_data[7:7] ;
assign n1026 = ~ ( n1025 ) ;
assign n1027 = sp[7:7] ;
assign n1028 =  ( n1026 ) ^ ( n1027 )  ;
assign n1029 =  ( n1028 ) ^ ( n330 )  ;
assign n1030 = i_wb_data[7:7] ;
assign n1031 = ~ ( n1030 ) ;
assign n1032 = sp[7:7] ;
assign n1033 =  ( n1031 ) ^ ( n1032 )  ;
assign n1034 =  ( n1033 ) ^ ( n330 )  ;
assign n1035 = ~ ( n1034 ) ;
assign n1036 =  ( n1024 ) ? ( n1029 ) : ( n1035 ) ;
assign n1037 =  ( n1021 ) ? ( bv_1_0_n2 ) : ( n1036 ) ;
assign n1038 =  ( n373 ) | ( n382 )  ;
assign n1039 = ki[15:15] ;
assign n1040 =  ( n1039 ) == ( bv_1_0_n2 )  ;
assign n1041 =  ( n1040 ) | ( n391 )  ;
assign n1042 = i_wb_data[8:8] ;
assign n1043 = ~ ( n1042 ) ;
assign n1044 = sp[8:8] ;
assign n1045 =  ( n1043 ) ^ ( n1044 )  ;
assign n1046 = i_wb_data[7:7] ;
assign n1047 = sp[7:7] ;
assign n1048 = ~ ( n1047 ) ;
assign n1049 =  ( n1046 ) | ( n1048 )  ;
assign n1050 = ~ ( n1049 ) ;
assign n1051 = ~ ( n330 ) ;
assign n1052 =  ( n137 ) | ( n1051 )  ;
assign n1053 = ~ ( n1052 ) ;
assign n1054 =  ( n1050 ) | ( n1053 )  ;
assign n1055 =  ( n1045 ) ^ ( n1054 )  ;
assign n1056 = i_wb_data[8:8] ;
assign n1057 = ~ ( n1056 ) ;
assign n1058 = sp[8:8] ;
assign n1059 =  ( n1057 ) ^ ( n1058 )  ;
assign n1060 =  ( n1059 ) ^ ( n1054 )  ;
assign n1061 = ~ ( n1060 ) ;
assign n1062 =  ( n1041 ) ? ( n1055 ) : ( n1061 ) ;
assign n1063 =  ( n1038 ) ? ( bv_1_0_n2 ) : ( n1062 ) ;
assign n1064 =  ( n1020 ) ? ( n1037 ) : ( n1063 ) ;
assign n1065 = ~ ( n1064 ) ;
assign n1066 =  ( n1019 ) | ( n1065 )  ;
assign n1067 = ~ ( n1066 ) ;
assign n1068 =  ( n1012 ) | ( n1067 )  ;
assign n1069 = ~ ( n1068 ) ;
assign n1070 =  ( n873 ) | ( n882 )  ;
assign n1071 =  ( n1070 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n1072 = ~ ( n941 ) ;
assign n1073 =  ( n1071 ) | ( n1072 )  ;
assign n1074 = ~ ( n1073 ) ;
assign n1075 = ~ ( n967 ) ;
assign n1076 = ~ ( n999 ) ;
assign n1077 =  ( n1075 ) | ( n1076 )  ;
assign n1078 = ~ ( n1077 ) ;
assign n1079 =  ( n1074 ) | ( n1078 )  ;
assign n1080 = ~ ( n1079 ) ;
assign n1081 =  ( n1069 ) | ( n1080 )  ;
assign n1082 = ~ ( n1081 ) ;
assign n1083 =  ( n1068 ) ^ ( n1079 )  ;
assign n1084 = ~ ( n1083 ) ;
assign n1085 =  ( n908 ) | ( n917 )  ;
assign n1086 =  ( n532 ) | ( n541 )  ;
assign n1087 =  ( n1086 ) ? ( bv_1_0_n2 ) : ( n939 ) ;
assign n1088 =  ( n532 ) | ( n541 )  ;
assign n1089 =  ( n1088 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n1090 =  ( n1085 ) ? ( n1087 ) : ( n1089 ) ;
assign n1091 =  ( bv_1_1_n5 ) ^ ( n1090 )  ;
assign n1092 =  ( n567 ) | ( n576 )  ;
assign n1093 =  ( n586 ) | ( n595 )  ;
assign n1094 =  ( n1093 ) ? ( bv_1_0_n2 ) : ( n965 ) ;
assign n1095 =  ( n586 ) | ( n595 )  ;
assign n1096 =  ( n1095 ) ? ( bv_1_0_n2 ) : ( n611 ) ;
assign n1097 =  ( n1092 ) ? ( n1094 ) : ( n1096 ) ;
assign n1098 =  ( n1091 ) ^ ( n1097 )  ;
assign n1099 =  ( n11 ) | ( n20 )  ;
assign n1100 =  ( n30 ) | ( n39 )  ;
assign n1101 =  ( n1100 ) ? ( bv_1_0_n2 ) : ( n997 ) ;
assign n1102 =  ( n30 ) | ( n39 )  ;
assign n1103 =  ( n1102 ) ? ( bv_1_0_n2 ) : ( n649 ) ;
assign n1104 =  ( n1099 ) ? ( n1101 ) : ( n1103 ) ;
assign n1105 =  ( n1098 ) ^ ( n1104 )  ;
assign n1106 =  ( n354 ) | ( n363 )  ;
assign n1107 =  ( n373 ) | ( n382 )  ;
assign n1108 =  ( n1107 ) ? ( bv_1_0_n2 ) : ( n1062 ) ;
assign n1109 =  ( n373 ) | ( n382 )  ;
assign n1110 = ki[15:15] ;
assign n1111 =  ( n1110 ) == ( bv_1_0_n2 )  ;
assign n1112 =  ( n1111 ) | ( n391 )  ;
assign n1113 = i_wb_data[9:9] ;
assign n1114 = ~ ( n1113 ) ;
assign n1115 = sp[9:9] ;
assign n1116 =  ( n1114 ) ^ ( n1115 )  ;
assign n1117 =  ( n1116 ) ^ ( n734 )  ;
assign n1118 =  ( n1112 ) ? ( n1117 ) : ( n985 ) ;
assign n1119 =  ( n1109 ) ? ( bv_1_0_n2 ) : ( n1118 ) ;
assign n1120 =  ( n1106 ) ? ( n1108 ) : ( n1119 ) ;
assign n1121 =  ( n1105 ) ^ ( n1120 )  ;
assign n1122 = ~ ( n1121 ) ;
assign n1123 =  ( n1084 ) | ( n1122 )  ;
assign n1124 = ~ ( n1123 ) ;
assign n1125 =  ( n1082 ) | ( n1124 )  ;
assign n1126 = ~ ( n1125 ) ;
assign n1127 = ~ ( n1090 ) ;
assign n1128 = ~ ( n1097 ) ;
assign n1129 =  ( n1127 ) | ( n1128 )  ;
assign n1130 = ~ ( n1104 ) ;
assign n1131 =  ( n1129 ) | ( n1130 )  ;
assign n1132 = ~ ( n1120 ) ;
assign n1133 =  ( n1131 ) | ( n1132 )  ;
assign n1134 = ~ ( n1133 ) ;
assign n1135 =  ( n1090 ) ^ ( n1097 )  ;
assign n1136 = ~ ( n1135 ) ;
assign n1137 =  ( n1104 ) ^ ( n1120 )  ;
assign n1138 = ~ ( n1137 ) ;
assign n1139 =  ( n1136 ) | ( n1138 )  ;
assign n1140 = ~ ( n1139 ) ;
assign n1141 =  ( n1134 ) | ( n1140 )  ;
assign n1142 =  ( n1090 ) ^ ( n1097 )  ;
assign n1143 =  ( n1142 ) ^ ( n1104 )  ;
assign n1144 =  ( n1143 ) ^ ( n1120 )  ;
assign n1145 =  ( n1141 ) | ( n1144 )  ;
assign n1146 = ~ ( n1090 ) ;
assign n1147 = ~ ( n1097 ) ;
assign n1148 =  ( n1146 ) | ( n1147 )  ;
assign n1149 = ~ ( n1148 ) ;
assign n1150 = ~ ( n1104 ) ;
assign n1151 = ~ ( n1120 ) ;
assign n1152 =  ( n1150 ) | ( n1151 )  ;
assign n1153 = ~ ( n1152 ) ;
assign n1154 =  ( n1149 ) | ( n1153 )  ;
assign n1155 =  ( n1145 ) ^ ( n1154 )  ;
assign n1156 =  ( n532 ) | ( n541 )  ;
assign n1157 =  ( n1156 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n1158 = ~ ( n1157 ) ;
assign n1159 =  ( n1155 ) ^ ( n1158 )  ;
assign n1160 =  ( n1159 ) ^ ( n624 )  ;
assign n1161 =  ( n1160 ) ^ ( n662 )  ;
assign n1162 = ~ ( n1161 ) ;
assign n1163 =  ( n1126 ) | ( n1162 )  ;
assign n1164 = ~ ( n1163 ) ;
assign n1165 =  ( n1125 ) ^ ( n1145 )  ;
assign n1166 =  ( n1165 ) ^ ( n1154 )  ;
assign n1167 =  ( n532 ) | ( n541 )  ;
assign n1168 =  ( n1167 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n1169 = ~ ( n1168 ) ;
assign n1170 =  ( n1166 ) ^ ( n1169 )  ;
assign n1171 =  ( n1170 ) ^ ( n624 )  ;
assign n1172 =  ( n1171 ) ^ ( n662 )  ;
assign n1173 = ~ ( n1172 ) ;
assign n1174 =  ( n354 ) | ( n363 )  ;
assign n1175 =  ( n373 ) | ( n382 )  ;
assign n1176 =  ( n1175 ) ? ( bv_1_0_n2 ) : ( n1118 ) ;
assign n1177 =  ( n373 ) | ( n382 )  ;
assign n1178 =  ( n1177 ) ? ( bv_1_0_n2 ) : ( n746 ) ;
assign n1179 =  ( n1174 ) ? ( n1176 ) : ( n1178 ) ;
assign n1180 = ~ ( n1179 ) ;
assign n1181 =  ( n1173 ) | ( n1180 )  ;
assign n1182 = ~ ( n1181 ) ;
assign n1183 =  ( n1164 ) | ( n1182 )  ;
assign n1184 = ~ ( n1183 ) ;
assign n1185 = ~ ( n1145 ) ;
assign n1186 = ~ ( n1154 ) ;
assign n1187 =  ( n1185 ) | ( n1186 )  ;
assign n1188 = ~ ( n1187 ) ;
assign n1189 =  ( n1145 ) ^ ( n1154 )  ;
assign n1190 = ~ ( n1189 ) ;
assign n1191 =  ( n532 ) | ( n541 )  ;
assign n1192 =  ( n1191 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n1193 = ~ ( n1192 ) ;
assign n1194 =  ( n1193 ) ^ ( n624 )  ;
assign n1195 =  ( n1194 ) ^ ( n662 )  ;
assign n1196 = ~ ( n1195 ) ;
assign n1197 =  ( n1190 ) | ( n1196 )  ;
assign n1198 = ~ ( n1197 ) ;
assign n1199 =  ( n1188 ) | ( n1198 )  ;
assign n1200 = ~ ( n1199 ) ;
assign n1201 =  ( n1184 ) | ( n1200 )  ;
assign n1202 = ~ ( n1201 ) ;
assign n1203 =  ( n1183 ) ^ ( n1199 )  ;
assign n1204 = ~ ( n1203 ) ;
assign n1205 =  ( bv_1_1_n5 ) ^ ( n666 )  ;
assign n1206 =  ( n1205 ) ^ ( n682 )  ;
assign n1207 =  ( n1206 ) ^ ( n697 )  ;
assign n1208 =  ( n1207 ) ^ ( n759 )  ;
assign n1209 = ~ ( n1208 ) ;
assign n1210 =  ( n1204 ) | ( n1209 )  ;
assign n1211 = ~ ( n1210 ) ;
assign n1212 =  ( n1202 ) | ( n1211 )  ;
assign n1213 = ~ ( n1212 ) ;
assign n1214 =  ( n666 ) ^ ( n682 )  ;
assign n1215 =  ( n1214 ) ^ ( n697 )  ;
assign n1216 =  ( n1215 ) ^ ( n759 )  ;
assign n1217 =  ( n763 ) | ( n1216 )  ;
assign n1218 =  ( n1217 ) ^ ( n778 )  ;
assign n1219 =  ( n586 ) | ( n595 )  ;
assign n1220 =  ( n1219 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n1221 = ~ ( n1220 ) ;
assign n1222 =  ( n1218 ) ^ ( n1221 )  ;
assign n1223 =  ( n1222 ) ^ ( n796 )  ;
assign n1224 =  ( n1223 ) ^ ( n803 )  ;
assign n1225 = ~ ( n1224 ) ;
assign n1226 =  ( n1213 ) | ( n1225 )  ;
assign n1227 = ~ ( n1226 ) ;
assign n1228 =  ( n666 ) ^ ( n682 )  ;
assign n1229 =  ( n1228 ) ^ ( n697 )  ;
assign n1230 =  ( n1229 ) ^ ( n759 )  ;
assign n1231 =  ( n763 ) | ( n1230 )  ;
assign n1232 =  ( n1212 ) ^ ( n1231 )  ;
assign n1233 =  ( n1232 ) ^ ( n778 )  ;
assign n1234 =  ( n586 ) | ( n595 )  ;
assign n1235 =  ( n1234 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n1236 = ~ ( n1235 ) ;
assign n1237 =  ( n1233 ) ^ ( n1236 )  ;
assign n1238 =  ( n1237 ) ^ ( n796 )  ;
assign n1239 =  ( n1238 ) ^ ( n803 )  ;
assign n1240 = ~ ( n1239 ) ;
assign n1241 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n1242 =  ( n1241 ) ^ ( n1199 )  ;
assign n1243 =  ( n1242 ) ^ ( n666 )  ;
assign n1244 =  ( n1243 ) ^ ( n682 )  ;
assign n1245 =  ( n1244 ) ^ ( n697 )  ;
assign n1246 =  ( n1245 ) ^ ( n759 )  ;
assign n1247 = ~ ( n1246 ) ;
assign n1248 =  ( n1240 ) | ( n1247 )  ;
assign n1249 = ki[7:7] ;
assign n1250 =  ( n1249 ) == ( bv_1_0_n2 )  ;
assign n1251 = ki[6:6] ;
assign n1252 =  ( n1251 ) == ( bv_1_1_n5 )  ;
assign n1253 =  ( n1250 ) | ( n1252 )  ;
assign n1254 = ki[5:5] ;
assign n1255 =  ( n1254 ) == ( bv_1_1_n5 )  ;
assign n1256 =  ( n1253 ) | ( n1255 )  ;
assign n1257 = ~ ( n1256 )  ;
assign n1258 = ki[7:7] ;
assign n1259 =  ( n1258 ) == ( bv_1_1_n5 )  ;
assign n1260 = ki[6:6] ;
assign n1261 =  ( n1260 ) == ( bv_1_0_n2 )  ;
assign n1262 =  ( n1259 ) | ( n1261 )  ;
assign n1263 = ki[5:5] ;
assign n1264 =  ( n1263 ) == ( bv_1_0_n2 )  ;
assign n1265 =  ( n1262 ) | ( n1264 )  ;
assign n1266 = ~ ( n1265 )  ;
assign n1267 =  ( n1257 ) | ( n1266 )  ;
assign n1268 =  ( n873 ) | ( n882 )  ;
assign n1269 = ki[7:7] ;
assign n1270 =  ( n1269 ) == ( bv_1_0_n2 )  ;
assign n1271 =  ( n1270 ) | ( n891 )  ;
assign n1272 = i_wb_data[14:14] ;
assign n1273 = ~ ( n1272 ) ;
assign n1274 = sp[14:14] ;
assign n1275 =  ( n1273 ) ^ ( n1274 )  ;
assign n1276 =  ( n1275 ) ^ ( n249 )  ;
assign n1277 =  ( n1271 ) ? ( n1276 ) : ( n256 ) ;
assign n1278 =  ( n1268 ) ? ( bv_1_0_n2 ) : ( n1277 ) ;
assign n1279 =  ( n873 ) | ( n882 )  ;
assign n1280 =  ( n1279 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n1281 =  ( n1267 ) ? ( n1278 ) : ( n1280 ) ;
assign n1282 = ~ ( n1281 ) ;
assign n1283 =  ( n908 ) | ( n917 )  ;
assign n1284 =  ( n532 ) | ( n541 )  ;
assign n1285 = ki[9:9] ;
assign n1286 =  ( n1285 ) == ( bv_1_0_n2 )  ;
assign n1287 =  ( n1286 ) | ( n550 )  ;
assign n1288 = i_wb_data[12:12] ;
assign n1289 = ~ ( n1288 ) ;
assign n1290 = sp[12:12] ;
assign n1291 =  ( n1289 ) ^ ( n1290 )  ;
assign n1292 =  ( n1291 ) ^ ( n427 )  ;
assign n1293 =  ( n1287 ) ? ( n1292 ) : ( n434 ) ;
assign n1294 =  ( n1284 ) ? ( bv_1_0_n2 ) : ( n1293 ) ;
assign n1295 =  ( n532 ) | ( n541 )  ;
assign n1296 =  ( n1295 ) ? ( bv_1_0_n2 ) : ( n928 ) ;
assign n1297 =  ( n1283 ) ? ( n1294 ) : ( n1296 ) ;
assign n1298 = ~ ( n1297 ) ;
assign n1299 =  ( n1282 ) | ( n1298 )  ;
assign n1300 =  ( n567 ) | ( n576 )  ;
assign n1301 =  ( n586 ) | ( n595 )  ;
assign n1302 = ki[11:11] ;
assign n1303 =  ( n1302 ) == ( bv_1_0_n2 )  ;
assign n1304 =  ( n1303 ) | ( n604 )  ;
assign n1305 = i_wb_data[10:10] ;
assign n1306 = ~ ( n1305 ) ;
assign n1307 = sp[10:10] ;
assign n1308 =  ( n1306 ) ^ ( n1307 )  ;
assign n1309 =  ( n1308 ) ^ ( n738 )  ;
assign n1310 =  ( n1304 ) ? ( n1309 ) : ( n745 ) ;
assign n1311 =  ( n1301 ) ? ( bv_1_0_n2 ) : ( n1310 ) ;
assign n1312 =  ( n586 ) | ( n595 )  ;
assign n1313 =  ( n1312 ) ? ( bv_1_0_n2 ) : ( n954 ) ;
assign n1314 =  ( n1300 ) ? ( n1311 ) : ( n1313 ) ;
assign n1315 = ~ ( n1314 ) ;
assign n1316 =  ( n1299 ) | ( n1315 )  ;
assign n1317 =  ( n11 ) | ( n20 )  ;
assign n1318 =  ( n30 ) | ( n39 )  ;
assign n1319 = ki[13:13] ;
assign n1320 =  ( n1319 ) == ( bv_1_0_n2 )  ;
assign n1321 =  ( n1320 ) | ( n48 )  ;
assign n1322 = i_wb_data[8:8] ;
assign n1323 = ~ ( n1322 ) ;
assign n1324 = sp[8:8] ;
assign n1325 =  ( n1323 ) ^ ( n1324 )  ;
assign n1326 =  ( n1325 ) ^ ( n1054 )  ;
assign n1327 =  ( n1321 ) ? ( n1326 ) : ( n1061 ) ;
assign n1328 =  ( n1318 ) ? ( bv_1_0_n2 ) : ( n1327 ) ;
assign n1329 =  ( n30 ) | ( n39 )  ;
assign n1330 =  ( n1329 ) ? ( bv_1_0_n2 ) : ( n986 ) ;
assign n1331 =  ( n1317 ) ? ( n1328 ) : ( n1330 ) ;
assign n1332 = ~ ( n1331 ) ;
assign n1333 =  ( n1316 ) | ( n1332 )  ;
assign n1334 = ~ ( n1333 ) ;
assign n1335 =  ( n1281 ) ^ ( n1297 )  ;
assign n1336 = ~ ( n1335 ) ;
assign n1337 =  ( n1314 ) ^ ( n1331 )  ;
assign n1338 = ~ ( n1337 ) ;
assign n1339 =  ( n1336 ) | ( n1338 )  ;
assign n1340 = ~ ( n1339 ) ;
assign n1341 =  ( n1334 ) | ( n1340 )  ;
assign n1342 =  ( n1281 ) ^ ( n1297 )  ;
assign n1343 =  ( n1342 ) ^ ( n1314 )  ;
assign n1344 =  ( n1343 ) ^ ( n1331 )  ;
assign n1345 = ~ ( n1344 ) ;
assign n1346 =  ( n354 ) | ( n363 )  ;
assign n1347 =  ( n373 ) | ( n382 )  ;
assign n1348 = ki[15:15] ;
assign n1349 =  ( n1348 ) == ( bv_1_0_n2 )  ;
assign n1350 =  ( n1349 ) | ( n391 )  ;
assign n1351 = i_wb_data[6:6] ;
assign n1352 = ~ ( n1351 ) ;
assign n1353 = sp[6:6] ;
assign n1354 =  ( n1352 ) ^ ( n1353 )  ;
assign n1355 = i_wb_data[5:5] ;
assign n1356 = sp[5:5] ;
assign n1357 = ~ ( n1356 ) ;
assign n1358 =  ( n1355 ) | ( n1357 )  ;
assign n1359 = ~ ( n1358 ) ;
assign n1360 = ~ ( n241 ) ;
assign n1361 =  ( n174 ) | ( n1360 )  ;
assign n1362 = ~ ( n1361 ) ;
assign n1363 =  ( n1359 ) | ( n1362 )  ;
assign n1364 =  ( n1354 ) ^ ( n1363 )  ;
assign n1365 = i_wb_data[6:6] ;
assign n1366 = ~ ( n1365 ) ;
assign n1367 = sp[6:6] ;
assign n1368 =  ( n1366 ) ^ ( n1367 )  ;
assign n1369 =  ( n1368 ) ^ ( n1363 )  ;
assign n1370 = ~ ( n1369 ) ;
assign n1371 =  ( n1350 ) ? ( n1364 ) : ( n1370 ) ;
assign n1372 =  ( n1347 ) ? ( bv_1_0_n2 ) : ( n1371 ) ;
assign n1373 =  ( n373 ) | ( n382 )  ;
assign n1374 =  ( n1373 ) ? ( bv_1_0_n2 ) : ( n1036 ) ;
assign n1375 =  ( n1346 ) ? ( n1372 ) : ( n1374 ) ;
assign n1376 = ~ ( n1375 ) ;
assign n1377 =  ( n1345 ) | ( n1376 )  ;
assign n1378 = ~ ( n1377 ) ;
assign n1379 =  ( n1341 ) | ( n1378 )  ;
assign n1380 = ~ ( n1379 ) ;
assign n1381 = ~ ( n1281 ) ;
assign n1382 = ~ ( n1297 ) ;
assign n1383 =  ( n1381 ) | ( n1382 )  ;
assign n1384 = ~ ( n1383 ) ;
assign n1385 = ~ ( n1314 ) ;
assign n1386 = ~ ( n1331 ) ;
assign n1387 =  ( n1385 ) | ( n1386 )  ;
assign n1388 = ~ ( n1387 ) ;
assign n1389 =  ( n1384 ) | ( n1388 )  ;
assign n1390 = ~ ( n1389 ) ;
assign n1391 =  ( n1380 ) | ( n1390 )  ;
assign n1392 = ~ ( n1391 ) ;
assign n1393 =  ( n1379 ) ^ ( n1389 )  ;
assign n1394 = ~ ( n1393 ) ;
assign n1395 =  ( n873 ) | ( n882 )  ;
assign n1396 =  ( n1395 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n1397 = ~ ( n1396 ) ;
assign n1398 =  ( n1397 ) ^ ( n941 )  ;
assign n1399 =  ( n1398 ) ^ ( n967 )  ;
assign n1400 =  ( n1399 ) ^ ( n999 )  ;
assign n1401 =  ( n1400 ) ^ ( n1064 )  ;
assign n1402 = ~ ( n1401 ) ;
assign n1403 =  ( n1394 ) | ( n1402 )  ;
assign n1404 = ~ ( n1403 ) ;
assign n1405 =  ( n1392 ) | ( n1404 )  ;
assign n1406 = ~ ( n1405 ) ;
assign n1407 =  ( bv_1_1_n5 ) ^ ( n1068 )  ;
assign n1408 =  ( n1407 ) ^ ( n1079 )  ;
assign n1409 =  ( n1408 ) ^ ( n1090 )  ;
assign n1410 =  ( n1409 ) ^ ( n1097 )  ;
assign n1411 =  ( n1410 ) ^ ( n1104 )  ;
assign n1412 =  ( n1411 ) ^ ( n1120 )  ;
assign n1413 = ~ ( n1412 ) ;
assign n1414 =  ( n1406 ) | ( n1413 )  ;
assign n1415 =  ( n1125 ) ^ ( n1145 )  ;
assign n1416 =  ( n1415 ) ^ ( n1154 )  ;
assign n1417 =  ( n532 ) | ( n541 )  ;
assign n1418 =  ( n1417 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n1419 = ~ ( n1418 ) ;
assign n1420 =  ( n1416 ) ^ ( n1419 )  ;
assign n1421 =  ( n1420 ) ^ ( n624 )  ;
assign n1422 =  ( n1421 ) ^ ( n662 )  ;
assign n1423 =  ( n1422 ) ^ ( n1179 )  ;
assign n1424 = ~ ( n1423 ) ;
assign n1425 =  ( n1414 ) | ( n1424 )  ;
assign n1426 = ~ ( n1425 ) ;
assign n1427 = ~ ( n1405 ) ;
assign n1428 =  ( bv_1_1_n5 ) ^ ( n1068 )  ;
assign n1429 =  ( n1428 ) ^ ( n1079 )  ;
assign n1430 =  ( n1429 ) ^ ( n1090 )  ;
assign n1431 =  ( n1430 ) ^ ( n1097 )  ;
assign n1432 =  ( n1431 ) ^ ( n1104 )  ;
assign n1433 =  ( n1432 ) ^ ( n1120 )  ;
assign n1434 = ~ ( n1433 ) ;
assign n1435 =  ( n1427 ) | ( n1434 )  ;
assign n1436 = ~ ( n1435 ) ;
assign n1437 =  ( n1436 ) ^ ( n1125 )  ;
assign n1438 =  ( n1437 ) ^ ( n1145 )  ;
assign n1439 =  ( n1438 ) ^ ( n1154 )  ;
assign n1440 =  ( n532 ) | ( n541 )  ;
assign n1441 =  ( n1440 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n1442 = ~ ( n1441 ) ;
assign n1443 =  ( n1439 ) ^ ( n1442 )  ;
assign n1444 =  ( n1443 ) ^ ( n624 )  ;
assign n1445 =  ( n1444 ) ^ ( n662 )  ;
assign n1446 =  ( n1445 ) ^ ( n1179 )  ;
assign n1447 = ~ ( n1446 ) ;
assign n1448 = ki[5:5] ;
assign n1449 =  ( n1448 ) == ( bv_1_0_n2 )  ;
assign n1450 = ki[4:4] ;
assign n1451 =  ( n1450 ) == ( bv_1_1_n5 )  ;
assign n1452 =  ( n1449 ) | ( n1451 )  ;
assign n1453 = ki[3:3] ;
assign n1454 =  ( n1453 ) == ( bv_1_1_n5 )  ;
assign n1455 =  ( n1452 ) | ( n1454 )  ;
assign n1456 = ~ ( n1455 )  ;
assign n1457 = ki[5:5] ;
assign n1458 =  ( n1457 ) == ( bv_1_1_n5 )  ;
assign n1459 = ki[4:4] ;
assign n1460 =  ( n1459 ) == ( bv_1_0_n2 )  ;
assign n1461 =  ( n1458 ) | ( n1460 )  ;
assign n1462 = ki[3:3] ;
assign n1463 =  ( n1462 ) == ( bv_1_0_n2 )  ;
assign n1464 =  ( n1461 ) | ( n1463 )  ;
assign n1465 = ~ ( n1464 )  ;
assign n1466 =  ( n1456 ) | ( n1465 )  ;
assign n1467 = ki[5:5] ;
assign n1468 =  ( n1467 ) == ( bv_1_0_n2 )  ;
assign n1469 = ki[4:4] ;
assign n1470 =  ( n1469 ) == ( bv_1_0_n2 )  ;
assign n1471 =  ( n1468 ) | ( n1470 )  ;
assign n1472 = ki[3:3] ;
assign n1473 =  ( n1472 ) == ( bv_1_0_n2 )  ;
assign n1474 =  ( n1471 ) | ( n1473 )  ;
assign n1475 = ~ ( n1474 )  ;
assign n1476 = ki[5:5] ;
assign n1477 =  ( n1476 ) == ( bv_1_1_n5 )  ;
assign n1478 = ki[4:4] ;
assign n1479 =  ( n1478 ) == ( bv_1_1_n5 )  ;
assign n1480 =  ( n1477 ) | ( n1479 )  ;
assign n1481 = ki[3:3] ;
assign n1482 =  ( n1481 ) == ( bv_1_1_n5 )  ;
assign n1483 =  ( n1480 ) | ( n1482 )  ;
assign n1484 = ~ ( n1483 )  ;
assign n1485 =  ( n1475 ) | ( n1484 )  ;
assign n1486 = ki[5:5] ;
assign n1487 =  ( n1486 ) == ( bv_1_0_n2 )  ;
assign n1488 = ki[4:4] ;
assign n1489 =  ( n1488 ) == ( bv_1_0_n2 )  ;
assign n1490 = ki[3:3] ;
assign n1491 =  ( n1490 ) == ( bv_1_0_n2 )  ;
assign n1492 =  ( n1489 ) | ( n1491 )  ;
assign n1493 = ~ ( n1492 )  ;
assign n1494 =  ( n1487 ) | ( n1493 )  ;
assign n1495 = i_wb_data[14:14] ;
assign n1496 = ~ ( n1495 ) ;
assign n1497 = sp[14:14] ;
assign n1498 =  ( n1496 ) ^ ( n1497 )  ;
assign n1499 =  ( n1498 ) ^ ( n249 )  ;
assign n1500 =  ( n1494 ) ? ( n1499 ) : ( n256 ) ;
assign n1501 =  ( n1485 ) ? ( bv_1_0_n2 ) : ( n1500 ) ;
assign n1502 =  ( n1475 ) | ( n1484 )  ;
assign n1503 = ki[5:5] ;
assign n1504 =  ( n1503 ) == ( bv_1_0_n2 )  ;
assign n1505 =  ( n1504 ) | ( n1493 )  ;
assign n1506 = i_wb_data[15:15] ;
assign n1507 = ~ ( n1506 ) ;
assign n1508 = sp[15:15] ;
assign n1509 =  ( n1507 ) ^ ( n1508 )  ;
assign n1510 =  ( n1509 ) ^ ( n334 )  ;
assign n1511 =  ( n1505 ) ? ( n1510 ) : ( n341 ) ;
assign n1512 =  ( n1502 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n1513 =  ( n1466 ) ? ( n1501 ) : ( n1512 ) ;
assign n1514 = ~ ( n1513 ) ;
assign n1515 =  ( n1257 ) | ( n1266 )  ;
assign n1516 =  ( n873 ) | ( n882 )  ;
assign n1517 = ki[7:7] ;
assign n1518 =  ( n1517 ) == ( bv_1_0_n2 )  ;
assign n1519 =  ( n1518 ) | ( n891 )  ;
assign n1520 = i_wb_data[12:12] ;
assign n1521 = ~ ( n1520 ) ;
assign n1522 = sp[12:12] ;
assign n1523 =  ( n1521 ) ^ ( n1522 )  ;
assign n1524 =  ( n1523 ) ^ ( n427 )  ;
assign n1525 =  ( n1519 ) ? ( n1524 ) : ( n434 ) ;
assign n1526 =  ( n1516 ) ? ( bv_1_0_n2 ) : ( n1525 ) ;
assign n1527 =  ( n873 ) | ( n882 )  ;
assign n1528 = ki[7:7] ;
assign n1529 =  ( n1528 ) == ( bv_1_0_n2 )  ;
assign n1530 =  ( n1529 ) | ( n891 )  ;
assign n1531 = i_wb_data[13:13] ;
assign n1532 = ~ ( n1531 ) ;
assign n1533 = sp[13:13] ;
assign n1534 =  ( n1532 ) ^ ( n1533 )  ;
assign n1535 =  ( n1534 ) ^ ( n245 )  ;
assign n1536 =  ( n1530 ) ? ( n1535 ) : ( n451 ) ;
assign n1537 =  ( n1527 ) ? ( bv_1_0_n2 ) : ( n1536 ) ;
assign n1538 =  ( n1515 ) ? ( n1526 ) : ( n1537 ) ;
assign n1539 = ~ ( n1538 ) ;
assign n1540 =  ( n1514 ) | ( n1539 )  ;
assign n1541 =  ( n908 ) | ( n917 )  ;
assign n1542 =  ( n532 ) | ( n541 )  ;
assign n1543 = ki[9:9] ;
assign n1544 =  ( n1543 ) == ( bv_1_0_n2 )  ;
assign n1545 =  ( n1544 ) | ( n550 )  ;
assign n1546 = i_wb_data[10:10] ;
assign n1547 = ~ ( n1546 ) ;
assign n1548 = sp[10:10] ;
assign n1549 =  ( n1547 ) ^ ( n1548 )  ;
assign n1550 =  ( n1549 ) ^ ( n738 )  ;
assign n1551 =  ( n1545 ) ? ( n1550 ) : ( n745 ) ;
assign n1552 =  ( n1542 ) ? ( bv_1_0_n2 ) : ( n1551 ) ;
assign n1553 =  ( n532 ) | ( n541 )  ;
assign n1554 = ki[9:9] ;
assign n1555 =  ( n1554 ) == ( bv_1_0_n2 )  ;
assign n1556 =  ( n1555 ) | ( n550 )  ;
assign n1557 = i_wb_data[11:11] ;
assign n1558 = ~ ( n1557 ) ;
assign n1559 = sp[11:11] ;
assign n1560 =  ( n1558 ) ^ ( n1559 )  ;
assign n1561 =  ( n1560 ) ^ ( n423 )  ;
assign n1562 =  ( n1556 ) ? ( n1561 ) : ( n648 ) ;
assign n1563 =  ( n1553 ) ? ( bv_1_0_n2 ) : ( n1562 ) ;
assign n1564 =  ( n1541 ) ? ( n1552 ) : ( n1563 ) ;
assign n1565 = ~ ( n1564 ) ;
assign n1566 =  ( n1540 ) | ( n1565 )  ;
assign n1567 =  ( n567 ) | ( n576 )  ;
assign n1568 =  ( n586 ) | ( n595 )  ;
assign n1569 = ki[11:11] ;
assign n1570 =  ( n1569 ) == ( bv_1_0_n2 )  ;
assign n1571 =  ( n1570 ) | ( n604 )  ;
assign n1572 = i_wb_data[8:8] ;
assign n1573 = ~ ( n1572 ) ;
assign n1574 = sp[8:8] ;
assign n1575 =  ( n1573 ) ^ ( n1574 )  ;
assign n1576 =  ( n1575 ) ^ ( n1054 )  ;
assign n1577 =  ( n1571 ) ? ( n1576 ) : ( n1061 ) ;
assign n1578 =  ( n1568 ) ? ( bv_1_0_n2 ) : ( n1577 ) ;
assign n1579 =  ( n586 ) | ( n595 )  ;
assign n1580 = ki[11:11] ;
assign n1581 =  ( n1580 ) == ( bv_1_0_n2 )  ;
assign n1582 =  ( n1581 ) | ( n604 )  ;
assign n1583 = i_wb_data[9:9] ;
assign n1584 = ~ ( n1583 ) ;
assign n1585 = sp[9:9] ;
assign n1586 =  ( n1584 ) ^ ( n1585 )  ;
assign n1587 =  ( n1586 ) ^ ( n734 )  ;
assign n1588 =  ( n1582 ) ? ( n1587 ) : ( n985 ) ;
assign n1589 =  ( n1579 ) ? ( bv_1_0_n2 ) : ( n1588 ) ;
assign n1590 =  ( n1567 ) ? ( n1578 ) : ( n1589 ) ;
assign n1591 = ~ ( n1590 ) ;
assign n1592 =  ( n1566 ) | ( n1591 )  ;
assign n1593 = ~ ( n1592 ) ;
assign n1594 =  ( n1513 ) ^ ( n1538 )  ;
assign n1595 = ~ ( n1594 ) ;
assign n1596 =  ( n1564 ) ^ ( n1590 )  ;
assign n1597 = ~ ( n1596 ) ;
assign n1598 =  ( n1595 ) | ( n1597 )  ;
assign n1599 = ~ ( n1598 ) ;
assign n1600 =  ( n1593 ) | ( n1599 )  ;
assign n1601 =  ( n1513 ) ^ ( n1538 )  ;
assign n1602 =  ( n1601 ) ^ ( n1564 )  ;
assign n1603 =  ( n1602 ) ^ ( n1590 )  ;
assign n1604 = ~ ( n1603 ) ;
assign n1605 =  ( n11 ) | ( n20 )  ;
assign n1606 =  ( n30 ) | ( n39 )  ;
assign n1607 = ki[13:13] ;
assign n1608 =  ( n1607 ) == ( bv_1_0_n2 )  ;
assign n1609 =  ( n1608 ) | ( n48 )  ;
assign n1610 = i_wb_data[6:6] ;
assign n1611 = ~ ( n1610 ) ;
assign n1612 = sp[6:6] ;
assign n1613 =  ( n1611 ) ^ ( n1612 )  ;
assign n1614 =  ( n1613 ) ^ ( n1363 )  ;
assign n1615 =  ( n1609 ) ? ( n1614 ) : ( n1370 ) ;
assign n1616 =  ( n1606 ) ? ( bv_1_0_n2 ) : ( n1615 ) ;
assign n1617 =  ( n30 ) | ( n39 )  ;
assign n1618 = ki[13:13] ;
assign n1619 =  ( n1618 ) == ( bv_1_0_n2 )  ;
assign n1620 =  ( n1619 ) | ( n48 )  ;
assign n1621 = i_wb_data[7:7] ;
assign n1622 = ~ ( n1621 ) ;
assign n1623 = sp[7:7] ;
assign n1624 =  ( n1622 ) ^ ( n1623 )  ;
assign n1625 =  ( n1624 ) ^ ( n330 )  ;
assign n1626 =  ( n1620 ) ? ( n1625 ) : ( n1035 ) ;
assign n1627 =  ( n1617 ) ? ( bv_1_0_n2 ) : ( n1626 ) ;
assign n1628 =  ( n1605 ) ? ( n1616 ) : ( n1627 ) ;
assign n1629 = ~ ( n1628 ) ;
assign n1630 =  ( n1604 ) | ( n1629 )  ;
assign n1631 = ~ ( n1630 ) ;
assign n1632 =  ( n1600 ) | ( n1631 )  ;
assign n1633 = ~ ( n1632 ) ;
assign n1634 = ~ ( n1513 ) ;
assign n1635 = ~ ( n1538 ) ;
assign n1636 =  ( n1634 ) | ( n1635 )  ;
assign n1637 = ~ ( n1636 ) ;
assign n1638 = ~ ( n1564 ) ;
assign n1639 = ~ ( n1590 ) ;
assign n1640 =  ( n1638 ) | ( n1639 )  ;
assign n1641 = ~ ( n1640 ) ;
assign n1642 =  ( n1637 ) | ( n1641 )  ;
assign n1643 = ~ ( n1642 ) ;
assign n1644 =  ( n1633 ) | ( n1643 )  ;
assign n1645 = ~ ( n1644 ) ;
assign n1646 =  ( n1632 ) ^ ( n1642 )  ;
assign n1647 = ~ ( n1646 ) ;
assign n1648 =  ( n1475 ) | ( n1484 )  ;
assign n1649 =  ( n1648 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n1650 = ~ ( n1649 ) ;
assign n1651 =  ( n1257 ) | ( n1266 )  ;
assign n1652 =  ( n873 ) | ( n882 )  ;
assign n1653 =  ( n1652 ) ? ( bv_1_0_n2 ) : ( n1536 ) ;
assign n1654 =  ( n873 ) | ( n882 )  ;
assign n1655 =  ( n1654 ) ? ( bv_1_0_n2 ) : ( n1277 ) ;
assign n1656 =  ( n1651 ) ? ( n1653 ) : ( n1655 ) ;
assign n1657 =  ( n1650 ) ^ ( n1656 )  ;
assign n1658 =  ( n908 ) | ( n917 )  ;
assign n1659 =  ( n532 ) | ( n541 )  ;
assign n1660 =  ( n1659 ) ? ( bv_1_0_n2 ) : ( n1562 ) ;
assign n1661 =  ( n532 ) | ( n541 )  ;
assign n1662 =  ( n1661 ) ? ( bv_1_0_n2 ) : ( n1293 ) ;
assign n1663 =  ( n1658 ) ? ( n1660 ) : ( n1662 ) ;
assign n1664 =  ( n1657 ) ^ ( n1663 )  ;
assign n1665 =  ( n567 ) | ( n576 )  ;
assign n1666 =  ( n586 ) | ( n595 )  ;
assign n1667 =  ( n1666 ) ? ( bv_1_0_n2 ) : ( n1588 ) ;
assign n1668 =  ( n586 ) | ( n595 )  ;
assign n1669 =  ( n1668 ) ? ( bv_1_0_n2 ) : ( n1310 ) ;
assign n1670 =  ( n1665 ) ? ( n1667 ) : ( n1669 ) ;
assign n1671 =  ( n1664 ) ^ ( n1670 )  ;
assign n1672 =  ( n11 ) | ( n20 )  ;
assign n1673 =  ( n30 ) | ( n39 )  ;
assign n1674 =  ( n1673 ) ? ( bv_1_0_n2 ) : ( n1626 ) ;
assign n1675 =  ( n30 ) | ( n39 )  ;
assign n1676 =  ( n1675 ) ? ( bv_1_0_n2 ) : ( n1327 ) ;
assign n1677 =  ( n1672 ) ? ( n1674 ) : ( n1676 ) ;
assign n1678 =  ( n1671 ) ^ ( n1677 )  ;
assign n1679 = ~ ( n1678 ) ;
assign n1680 =  ( n1647 ) | ( n1679 )  ;
assign n1681 = ~ ( n1680 ) ;
assign n1682 =  ( n1645 ) | ( n1681 )  ;
assign n1683 = ~ ( n1682 ) ;
assign n1684 =  ( n1475 ) | ( n1484 )  ;
assign n1685 =  ( n1684 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n1686 = ~ ( n1656 ) ;
assign n1687 =  ( n1685 ) | ( n1686 )  ;
assign n1688 = ~ ( n1663 ) ;
assign n1689 =  ( n1687 ) | ( n1688 )  ;
assign n1690 = ~ ( n1670 ) ;
assign n1691 =  ( n1689 ) | ( n1690 )  ;
assign n1692 = ~ ( n1691 ) ;
assign n1693 =  ( n1475 ) | ( n1484 )  ;
assign n1694 =  ( n1693 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n1695 = ~ ( n1694 ) ;
assign n1696 =  ( n1695 ) ^ ( n1656 )  ;
assign n1697 = ~ ( n1696 ) ;
assign n1698 =  ( n1663 ) ^ ( n1670 )  ;
assign n1699 = ~ ( n1698 ) ;
assign n1700 =  ( n1697 ) | ( n1699 )  ;
assign n1701 = ~ ( n1700 ) ;
assign n1702 =  ( n1692 ) | ( n1701 )  ;
assign n1703 =  ( n1475 ) | ( n1484 )  ;
assign n1704 =  ( n1703 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n1705 = ~ ( n1704 ) ;
assign n1706 =  ( n1705 ) ^ ( n1656 )  ;
assign n1707 =  ( n1706 ) ^ ( n1663 )  ;
assign n1708 =  ( n1707 ) ^ ( n1670 )  ;
assign n1709 = ~ ( n1708 ) ;
assign n1710 = ~ ( n1677 ) ;
assign n1711 =  ( n1709 ) | ( n1710 )  ;
assign n1712 = ~ ( n1711 ) ;
assign n1713 =  ( n1702 ) | ( n1712 )  ;
assign n1714 =  ( n1475 ) | ( n1484 )  ;
assign n1715 =  ( n1714 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n1716 = ~ ( n1656 ) ;
assign n1717 =  ( n1715 ) | ( n1716 )  ;
assign n1718 = ~ ( n1717 ) ;
assign n1719 = ~ ( n1663 ) ;
assign n1720 = ~ ( n1670 ) ;
assign n1721 =  ( n1719 ) | ( n1720 )  ;
assign n1722 = ~ ( n1721 ) ;
assign n1723 =  ( n1718 ) | ( n1722 )  ;
assign n1724 =  ( n1713 ) ^ ( n1723 )  ;
assign n1725 =  ( n1724 ) ^ ( n1281 )  ;
assign n1726 =  ( n1725 ) ^ ( n1297 )  ;
assign n1727 =  ( n1726 ) ^ ( n1314 )  ;
assign n1728 =  ( n1727 ) ^ ( n1331 )  ;
assign n1729 =  ( n1728 ) ^ ( n1375 )  ;
assign n1730 = ~ ( n1729 ) ;
assign n1731 =  ( n1683 ) | ( n1730 )  ;
assign n1732 = ~ ( n1731 ) ;
assign n1733 =  ( n1682 ) ^ ( n1713 )  ;
assign n1734 =  ( n1733 ) ^ ( n1723 )  ;
assign n1735 =  ( n1734 ) ^ ( n1281 )  ;
assign n1736 =  ( n1735 ) ^ ( n1297 )  ;
assign n1737 =  ( n1736 ) ^ ( n1314 )  ;
assign n1738 =  ( n1737 ) ^ ( n1331 )  ;
assign n1739 =  ( n1738 ) ^ ( n1375 )  ;
assign n1740 =  ( n1732 ) | ( n1739 )  ;
assign n1741 = ~ ( n1740 ) ;
assign n1742 = ~ ( n1713 ) ;
assign n1743 = ~ ( n1723 ) ;
assign n1744 =  ( n1742 ) | ( n1743 )  ;
assign n1745 = ~ ( n1744 ) ;
assign n1746 =  ( n1713 ) ^ ( n1723 )  ;
assign n1747 = ~ ( n1746 ) ;
assign n1748 =  ( n1281 ) ^ ( n1297 )  ;
assign n1749 =  ( n1748 ) ^ ( n1314 )  ;
assign n1750 =  ( n1749 ) ^ ( n1331 )  ;
assign n1751 =  ( n1750 ) ^ ( n1375 )  ;
assign n1752 = ~ ( n1751 ) ;
assign n1753 =  ( n1747 ) | ( n1752 )  ;
assign n1754 = ~ ( n1753 ) ;
assign n1755 =  ( n1745 ) | ( n1754 )  ;
assign n1756 = ~ ( n1755 ) ;
assign n1757 =  ( n1741 ) | ( n1756 )  ;
assign n1758 = ~ ( n1757 ) ;
assign n1759 =  ( n1740 ) ^ ( n1755 )  ;
assign n1760 = ~ ( n1759 ) ;
assign n1761 =  ( n1379 ) ^ ( n1389 )  ;
assign n1762 =  ( n873 ) | ( n882 )  ;
assign n1763 =  ( n1762 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n1764 = ~ ( n1763 ) ;
assign n1765 =  ( n1761 ) ^ ( n1764 )  ;
assign n1766 =  ( n1765 ) ^ ( n941 )  ;
assign n1767 =  ( n1766 ) ^ ( n967 )  ;
assign n1768 =  ( n1767 ) ^ ( n999 )  ;
assign n1769 =  ( n1768 ) ^ ( n1064 )  ;
assign n1770 = ~ ( n1769 ) ;
assign n1771 =  ( n1760 ) | ( n1770 )  ;
assign n1772 = ~ ( n1771 ) ;
assign n1773 =  ( n1758 ) | ( n1772 )  ;
assign n1774 = ~ ( n1773 ) ;
assign n1775 =  ( n1447 ) | ( n1774 )  ;
assign n1776 =  ( bv_1_1_n5 ) ^ ( n1405 )  ;
assign n1777 =  ( n1776 ) ^ ( n1068 )  ;
assign n1778 =  ( n1777 ) ^ ( n1079 )  ;
assign n1779 =  ( n1778 ) ^ ( n1090 )  ;
assign n1780 =  ( n1779 ) ^ ( n1097 )  ;
assign n1781 =  ( n1780 ) ^ ( n1104 )  ;
assign n1782 =  ( n1781 ) ^ ( n1120 )  ;
assign n1783 = ~ ( n1782 ) ;
assign n1784 =  ( n1775 ) | ( n1783 )  ;
assign n1785 = ~ ( n1784 ) ;
assign n1786 =  ( n1426 ) | ( n1785 )  ;
assign n1787 = ~ ( n1786 ) ;
assign n1788 =  ( n1248 ) | ( n1787 )  ;
assign n1789 = ~ ( n1788 ) ;
assign n1790 =  ( n1227 ) | ( n1789 )  ;
assign n1791 = ~ ( n1790 ) ;
assign n1792 =  ( n864 ) | ( n1791 )  ;
assign n1793 = ~ ( n1792 ) ;
assign n1794 =  ( n845 ) | ( n1793 )  ;
assign n1795 = ~ ( n518 ) ;
assign n1796 =  ( bv_1_1_n5 ) ^ ( n488 )  ;
assign n1797 =  ( n1796 ) ^ ( n504 )  ;
assign n1798 = ~ ( n1797 ) ;
assign n1799 =  ( n1795 ) | ( n1798 )  ;
assign n1800 = ~ ( n856 ) ;
assign n1801 =  ( n1799 ) | ( n1800 )  ;
assign n1802 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n1803 =  ( n1802 ) ^ ( n823 )  ;
assign n1804 =  ( n1803 ) ^ ( n344 )  ;
assign n1805 =  ( n1804 ) ^ ( n454 )  ;
assign n1806 = ~ ( n1805 ) ;
assign n1807 =  ( n1801 ) | ( n1806 )  ;
assign n1808 = ~ ( n1239 ) ;
assign n1809 =  ( n1807 ) | ( n1808 )  ;
assign n1810 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n1811 =  ( n1810 ) ^ ( n1199 )  ;
assign n1812 =  ( n1811 ) ^ ( n666 )  ;
assign n1813 =  ( n1812 ) ^ ( n682 )  ;
assign n1814 =  ( n1813 ) ^ ( n697 )  ;
assign n1815 =  ( n1814 ) ^ ( n759 )  ;
assign n1816 = ~ ( n1815 ) ;
assign n1817 =  ( n1809 ) | ( n1816 )  ;
assign n1818 = ~ ( n1446 ) ;
assign n1819 =  ( n1817 ) | ( n1818 )  ;
assign n1820 =  ( bv_1_1_n5 ) ^ ( n1773 )  ;
assign n1821 =  ( n1820 ) ^ ( n1405 )  ;
assign n1822 =  ( n1821 ) ^ ( n1068 )  ;
assign n1823 =  ( n1822 ) ^ ( n1079 )  ;
assign n1824 =  ( n1823 ) ^ ( n1090 )  ;
assign n1825 =  ( n1824 ) ^ ( n1097 )  ;
assign n1826 =  ( n1825 ) ^ ( n1104 )  ;
assign n1827 =  ( n1826 ) ^ ( n1120 )  ;
assign n1828 = ~ ( n1827 ) ;
assign n1829 =  ( n1819 ) | ( n1828 )  ;
assign n1830 = ki[3:3] ;
assign n1831 =  ( n1830 ) == ( bv_1_0_n2 )  ;
assign n1832 = ki[2:2] ;
assign n1833 =  ( n1832 ) == ( bv_1_0_n2 )  ;
assign n1834 =  ( n1831 ) | ( n1833 )  ;
assign n1835 = ki[1:1] ;
assign n1836 =  ( n1835 ) == ( bv_1_0_n2 )  ;
assign n1837 =  ( n1834 ) | ( n1836 )  ;
assign n1838 = ~ ( n1837 )  ;
assign n1839 = ki[3:3] ;
assign n1840 =  ( n1839 ) == ( bv_1_1_n5 )  ;
assign n1841 = ki[2:2] ;
assign n1842 =  ( n1841 ) == ( bv_1_1_n5 )  ;
assign n1843 =  ( n1840 ) | ( n1842 )  ;
assign n1844 = ki[1:1] ;
assign n1845 =  ( n1844 ) == ( bv_1_1_n5 )  ;
assign n1846 =  ( n1843 ) | ( n1845 )  ;
assign n1847 = ~ ( n1846 )  ;
assign n1848 =  ( n1838 ) | ( n1847 )  ;
assign n1849 = ki[3:3] ;
assign n1850 =  ( n1849 ) == ( bv_1_0_n2 )  ;
assign n1851 = ki[2:2] ;
assign n1852 =  ( n1851 ) == ( bv_1_0_n2 )  ;
assign n1853 = ki[1:1] ;
assign n1854 =  ( n1853 ) == ( bv_1_0_n2 )  ;
assign n1855 =  ( n1852 ) | ( n1854 )  ;
assign n1856 = ~ ( n1855 )  ;
assign n1857 =  ( n1850 ) | ( n1856 )  ;
assign n1858 = i_wb_data[15:15] ;
assign n1859 = ~ ( n1858 ) ;
assign n1860 = sp[15:15] ;
assign n1861 =  ( n1859 ) ^ ( n1860 )  ;
assign n1862 =  ( n1861 ) ^ ( n334 )  ;
assign n1863 =  ( n1857 ) ? ( n1862 ) : ( n341 ) ;
assign n1864 =  ( n1848 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n1865 =  ( n1456 ) | ( n1465 )  ;
assign n1866 =  ( n1475 ) | ( n1484 )  ;
assign n1867 = ki[5:5] ;
assign n1868 =  ( n1867 ) == ( bv_1_0_n2 )  ;
assign n1869 =  ( n1868 ) | ( n1493 )  ;
assign n1870 = i_wb_data[13:13] ;
assign n1871 = ~ ( n1870 ) ;
assign n1872 = sp[13:13] ;
assign n1873 =  ( n1871 ) ^ ( n1872 )  ;
assign n1874 =  ( n1873 ) ^ ( n245 )  ;
assign n1875 =  ( n1869 ) ? ( n1874 ) : ( n451 ) ;
assign n1876 =  ( n1866 ) ? ( bv_1_0_n2 ) : ( n1875 ) ;
assign n1877 =  ( n1475 ) | ( n1484 )  ;
assign n1878 =  ( n1877 ) ? ( bv_1_0_n2 ) : ( n1500 ) ;
assign n1879 =  ( n1865 ) ? ( n1876 ) : ( n1878 ) ;
assign n1880 = ~ ( n1879 ) ;
assign n1881 =  ( n1864 ) | ( n1880 )  ;
assign n1882 =  ( n1257 ) | ( n1266 )  ;
assign n1883 =  ( n873 ) | ( n882 )  ;
assign n1884 = ki[7:7] ;
assign n1885 =  ( n1884 ) == ( bv_1_0_n2 )  ;
assign n1886 =  ( n1885 ) | ( n891 )  ;
assign n1887 = i_wb_data[11:11] ;
assign n1888 = ~ ( n1887 ) ;
assign n1889 = sp[11:11] ;
assign n1890 =  ( n1888 ) ^ ( n1889 )  ;
assign n1891 =  ( n1890 ) ^ ( n423 )  ;
assign n1892 =  ( n1886 ) ? ( n1891 ) : ( n648 ) ;
assign n1893 =  ( n1883 ) ? ( bv_1_0_n2 ) : ( n1892 ) ;
assign n1894 =  ( n873 ) | ( n882 )  ;
assign n1895 =  ( n1894 ) ? ( bv_1_0_n2 ) : ( n1525 ) ;
assign n1896 =  ( n1882 ) ? ( n1893 ) : ( n1895 ) ;
assign n1897 = ~ ( n1896 ) ;
assign n1898 =  ( n1881 ) | ( n1897 )  ;
assign n1899 =  ( n908 ) | ( n917 )  ;
assign n1900 =  ( n532 ) | ( n541 )  ;
assign n1901 = ki[9:9] ;
assign n1902 =  ( n1901 ) == ( bv_1_0_n2 )  ;
assign n1903 =  ( n1902 ) | ( n550 )  ;
assign n1904 = i_wb_data[9:9] ;
assign n1905 = ~ ( n1904 ) ;
assign n1906 = sp[9:9] ;
assign n1907 =  ( n1905 ) ^ ( n1906 )  ;
assign n1908 =  ( n1907 ) ^ ( n734 )  ;
assign n1909 =  ( n1903 ) ? ( n1908 ) : ( n985 ) ;
assign n1910 =  ( n1900 ) ? ( bv_1_0_n2 ) : ( n1909 ) ;
assign n1911 =  ( n532 ) | ( n541 )  ;
assign n1912 =  ( n1911 ) ? ( bv_1_0_n2 ) : ( n1551 ) ;
assign n1913 =  ( n1899 ) ? ( n1910 ) : ( n1912 ) ;
assign n1914 = ~ ( n1913 ) ;
assign n1915 =  ( n1898 ) | ( n1914 )  ;
assign n1916 = ~ ( n1915 ) ;
assign n1917 =  ( n1838 ) | ( n1847 )  ;
assign n1918 =  ( n1917 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n1919 = ~ ( n1918 ) ;
assign n1920 =  ( n1919 ) ^ ( n1879 )  ;
assign n1921 = ~ ( n1920 ) ;
assign n1922 =  ( n1896 ) ^ ( n1913 )  ;
assign n1923 = ~ ( n1922 ) ;
assign n1924 =  ( n1921 ) | ( n1923 )  ;
assign n1925 = ~ ( n1924 ) ;
assign n1926 =  ( n1916 ) | ( n1925 )  ;
assign n1927 =  ( n1838 ) | ( n1847 )  ;
assign n1928 =  ( n1927 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n1929 = ~ ( n1928 ) ;
assign n1930 =  ( n1929 ) ^ ( n1879 )  ;
assign n1931 =  ( n1930 ) ^ ( n1896 )  ;
assign n1932 =  ( n1931 ) ^ ( n1913 )  ;
assign n1933 = ~ ( n1932 ) ;
assign n1934 =  ( n567 ) | ( n576 )  ;
assign n1935 =  ( n586 ) | ( n595 )  ;
assign n1936 = ki[11:11] ;
assign n1937 =  ( n1936 ) == ( bv_1_0_n2 )  ;
assign n1938 =  ( n1937 ) | ( n604 )  ;
assign n1939 = i_wb_data[7:7] ;
assign n1940 = ~ ( n1939 ) ;
assign n1941 = sp[7:7] ;
assign n1942 =  ( n1940 ) ^ ( n1941 )  ;
assign n1943 =  ( n1942 ) ^ ( n330 )  ;
assign n1944 =  ( n1938 ) ? ( n1943 ) : ( n1035 ) ;
assign n1945 =  ( n1935 ) ? ( bv_1_0_n2 ) : ( n1944 ) ;
assign n1946 =  ( n586 ) | ( n595 )  ;
assign n1947 =  ( n1946 ) ? ( bv_1_0_n2 ) : ( n1577 ) ;
assign n1948 =  ( n1934 ) ? ( n1945 ) : ( n1947 ) ;
assign n1949 = ~ ( n1948 ) ;
assign n1950 =  ( n1933 ) | ( n1949 )  ;
assign n1951 = ~ ( n1950 ) ;
assign n1952 =  ( n1926 ) | ( n1951 )  ;
assign n1953 = ~ ( n1952 ) ;
assign n1954 =  ( n1838 ) | ( n1847 )  ;
assign n1955 =  ( n1954 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n1956 = ~ ( n1879 ) ;
assign n1957 =  ( n1955 ) | ( n1956 )  ;
assign n1958 = ~ ( n1957 ) ;
assign n1959 = ~ ( n1896 ) ;
assign n1960 = ~ ( n1913 ) ;
assign n1961 =  ( n1959 ) | ( n1960 )  ;
assign n1962 = ~ ( n1961 ) ;
assign n1963 =  ( n1958 ) | ( n1962 )  ;
assign n1964 = ~ ( n1963 ) ;
assign n1965 =  ( n1953 ) | ( n1964 )  ;
assign n1966 =  ( n1513 ) ^ ( n1538 )  ;
assign n1967 =  ( n1966 ) ^ ( n1564 )  ;
assign n1968 =  ( n1967 ) ^ ( n1590 )  ;
assign n1969 =  ( n1968 ) ^ ( n1628 )  ;
assign n1970 = ~ ( n1969 ) ;
assign n1971 =  ( n1965 ) | ( n1970 )  ;
assign n1972 =  ( n354 ) | ( n363 )  ;
assign n1973 =  ( n373 ) | ( n382 )  ;
assign n1974 = ki[15:15] ;
assign n1975 =  ( n1974 ) == ( bv_1_0_n2 )  ;
assign n1976 =  ( n1975 ) | ( n391 )  ;
assign n1977 = i_wb_data[4:4] ;
assign n1978 = ~ ( n1977 ) ;
assign n1979 = sp[4:4] ;
assign n1980 =  ( n1978 ) ^ ( n1979 )  ;
assign n1981 = i_wb_data[3:3] ;
assign n1982 = sp[3:3] ;
assign n1983 = ~ ( n1982 ) ;
assign n1984 =  ( n1981 ) | ( n1983 )  ;
assign n1985 = ~ ( n1984 ) ;
assign n1986 = ~ ( n326 ) ;
assign n1987 =  ( n197 ) | ( n1986 )  ;
assign n1988 = ~ ( n1987 ) ;
assign n1989 =  ( n1985 ) | ( n1988 )  ;
assign n1990 =  ( n1980 ) ^ ( n1989 )  ;
assign n1991 = i_wb_data[4:4] ;
assign n1992 = ~ ( n1991 ) ;
assign n1993 = sp[4:4] ;
assign n1994 =  ( n1992 ) ^ ( n1993 )  ;
assign n1995 =  ( n1994 ) ^ ( n1989 )  ;
assign n1996 = ~ ( n1995 ) ;
assign n1997 =  ( n1976 ) ? ( n1990 ) : ( n1996 ) ;
assign n1998 =  ( n1973 ) ? ( bv_1_0_n2 ) : ( n1997 ) ;
assign n1999 =  ( n373 ) | ( n382 )  ;
assign n2000 = ki[15:15] ;
assign n2001 =  ( n2000 ) == ( bv_1_0_n2 )  ;
assign n2002 =  ( n2001 ) | ( n391 )  ;
assign n2003 = i_wb_data[5:5] ;
assign n2004 = ~ ( n2003 ) ;
assign n2005 = sp[5:5] ;
assign n2006 =  ( n2004 ) ^ ( n2005 )  ;
assign n2007 =  ( n2006 ) ^ ( n241 )  ;
assign n2008 = i_wb_data[5:5] ;
assign n2009 = ~ ( n2008 ) ;
assign n2010 = sp[5:5] ;
assign n2011 =  ( n2009 ) ^ ( n2010 )  ;
assign n2012 =  ( n2011 ) ^ ( n241 )  ;
assign n2013 = ~ ( n2012 ) ;
assign n2014 =  ( n2002 ) ? ( n2007 ) : ( n2013 ) ;
assign n2015 =  ( n1999 ) ? ( bv_1_0_n2 ) : ( n2014 ) ;
assign n2016 =  ( n1972 ) ? ( n1998 ) : ( n2015 ) ;
assign n2017 = ~ ( n2016 ) ;
assign n2018 =  ( n1971 ) | ( n2017 )  ;
assign n2019 = ~ ( n2018 ) ;
assign n2020 =  ( n1952 ) ^ ( n1963 )  ;
assign n2021 = ~ ( n2020 ) ;
assign n2022 =  ( n1513 ) ^ ( n1538 )  ;
assign n2023 =  ( n2022 ) ^ ( n1564 )  ;
assign n2024 =  ( n2023 ) ^ ( n1590 )  ;
assign n2025 =  ( n2024 ) ^ ( n1628 )  ;
assign n2026 =  ( n2025 ) ^ ( n2016 )  ;
assign n2027 = ~ ( n2026 ) ;
assign n2028 =  ( n2021 ) | ( n2027 )  ;
assign n2029 = ~ ( n2028 ) ;
assign n2030 =  ( n2019 ) | ( n2029 )  ;
assign n2031 =  ( n1952 ) ^ ( n1963 )  ;
assign n2032 =  ( n2031 ) ^ ( n1513 )  ;
assign n2033 =  ( n2032 ) ^ ( n1538 )  ;
assign n2034 =  ( n2033 ) ^ ( n1564 )  ;
assign n2035 =  ( n2034 ) ^ ( n1590 )  ;
assign n2036 =  ( n2035 ) ^ ( n1628 )  ;
assign n2037 =  ( n2036 ) ^ ( n2016 )  ;
assign n2038 =  ( n2030 ) | ( n2037 )  ;
assign n2039 = ~ ( n2038 ) ;
assign n2040 = ~ ( n1952 ) ;
assign n2041 = ~ ( n1963 ) ;
assign n2042 =  ( n2040 ) | ( n2041 )  ;
assign n2043 = ~ ( n2042 ) ;
assign n2044 =  ( n1513 ) ^ ( n1538 )  ;
assign n2045 =  ( n2044 ) ^ ( n1564 )  ;
assign n2046 =  ( n2045 ) ^ ( n1590 )  ;
assign n2047 =  ( n2046 ) ^ ( n1628 )  ;
assign n2048 = ~ ( n2047 ) ;
assign n2049 = ~ ( n2016 ) ;
assign n2050 =  ( n2048 ) | ( n2049 )  ;
assign n2051 = ~ ( n2050 ) ;
assign n2052 =  ( n2043 ) | ( n2051 )  ;
assign n2053 = ~ ( n2052 ) ;
assign n2054 =  ( n2039 ) | ( n2053 )  ;
assign n2055 = ~ ( n2054 ) ;
assign n2056 =  ( n2038 ) ^ ( n2052 )  ;
assign n2057 = ~ ( n2056 ) ;
assign n2058 =  ( n1632 ) ^ ( n1642 )  ;
assign n2059 =  ( n1475 ) | ( n1484 )  ;
assign n2060 =  ( n2059 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n2061 = ~ ( n2060 ) ;
assign n2062 =  ( n2058 ) ^ ( n2061 )  ;
assign n2063 =  ( n2062 ) ^ ( n1656 )  ;
assign n2064 =  ( n2063 ) ^ ( n1663 )  ;
assign n2065 =  ( n2064 ) ^ ( n1670 )  ;
assign n2066 =  ( n2065 ) ^ ( n1677 )  ;
assign n2067 = ~ ( n2066 ) ;
assign n2068 =  ( n2057 ) | ( n2067 )  ;
assign n2069 = ~ ( n2068 ) ;
assign n2070 =  ( n2055 ) | ( n2069 )  ;
assign n2071 = ~ ( n2070 ) ;
assign n2072 =  ( bv_1_1_n5 ) ^ ( n1682 )  ;
assign n2073 =  ( n2072 ) ^ ( n1713 )  ;
assign n2074 =  ( n2073 ) ^ ( n1723 )  ;
assign n2075 =  ( n2074 ) ^ ( n1281 )  ;
assign n2076 =  ( n2075 ) ^ ( n1297 )  ;
assign n2077 =  ( n2076 ) ^ ( n1314 )  ;
assign n2078 =  ( n2077 ) ^ ( n1331 )  ;
assign n2079 =  ( n2078 ) ^ ( n1375 )  ;
assign n2080 = ~ ( n2079 ) ;
assign n2081 =  ( n2071 ) | ( n2080 )  ;
assign n2082 =  ( n1740 ) ^ ( n1755 )  ;
assign n2083 =  ( n2082 ) ^ ( n1379 )  ;
assign n2084 =  ( n2083 ) ^ ( n1389 )  ;
assign n2085 =  ( n873 ) | ( n882 )  ;
assign n2086 =  ( n2085 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n2087 = ~ ( n2086 ) ;
assign n2088 =  ( n2084 ) ^ ( n2087 )  ;
assign n2089 =  ( n2088 ) ^ ( n941 )  ;
assign n2090 =  ( n2089 ) ^ ( n967 )  ;
assign n2091 =  ( n2090 ) ^ ( n999 )  ;
assign n2092 =  ( n2091 ) ^ ( n1064 )  ;
assign n2093 = ~ ( n2092 ) ;
assign n2094 =  ( n2081 ) | ( n2093 )  ;
assign n2095 = ~ ( n2094 ) ;
assign n2096 = ~ ( n2070 ) ;
assign n2097 =  ( n2096 ) | ( n2080 )  ;
assign n2098 = ~ ( n2097 ) ;
assign n2099 =  ( n2098 ) ^ ( n1740 )  ;
assign n2100 =  ( n2099 ) ^ ( n1755 )  ;
assign n2101 =  ( n2100 ) ^ ( n1379 )  ;
assign n2102 =  ( n2101 ) ^ ( n1389 )  ;
assign n2103 =  ( n873 ) | ( n882 )  ;
assign n2104 =  ( n2103 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n2105 = ~ ( n2104 ) ;
assign n2106 =  ( n2102 ) ^ ( n2105 )  ;
assign n2107 =  ( n2106 ) ^ ( n941 )  ;
assign n2108 =  ( n2107 ) ^ ( n967 )  ;
assign n2109 =  ( n2108 ) ^ ( n999 )  ;
assign n2110 =  ( n2109 ) ^ ( n1064 )  ;
assign n2111 = ~ ( n2110 ) ;
assign n2112 = ki[3:3] ;
assign n2113 =  ( n2112 ) == ( bv_1_0_n2 )  ;
assign n2114 = ki[2:2] ;
assign n2115 =  ( n2114 ) == ( bv_1_1_n5 )  ;
assign n2116 =  ( n2113 ) | ( n2115 )  ;
assign n2117 = ki[1:1] ;
assign n2118 =  ( n2117 ) == ( bv_1_1_n5 )  ;
assign n2119 =  ( n2116 ) | ( n2118 )  ;
assign n2120 = ~ ( n2119 )  ;
assign n2121 = ki[3:3] ;
assign n2122 =  ( n2121 ) == ( bv_1_1_n5 )  ;
assign n2123 = ki[2:2] ;
assign n2124 =  ( n2123 ) == ( bv_1_0_n2 )  ;
assign n2125 =  ( n2122 ) | ( n2124 )  ;
assign n2126 = ki[1:1] ;
assign n2127 =  ( n2126 ) == ( bv_1_0_n2 )  ;
assign n2128 =  ( n2125 ) | ( n2127 )  ;
assign n2129 = ~ ( n2128 )  ;
assign n2130 =  ( n2120 ) | ( n2129 )  ;
assign n2131 =  ( n1838 ) | ( n1847 )  ;
assign n2132 = ki[3:3] ;
assign n2133 =  ( n2132 ) == ( bv_1_0_n2 )  ;
assign n2134 =  ( n2133 ) | ( n1856 )  ;
assign n2135 = i_wb_data[14:14] ;
assign n2136 = ~ ( n2135 ) ;
assign n2137 = sp[14:14] ;
assign n2138 =  ( n2136 ) ^ ( n2137 )  ;
assign n2139 =  ( n2138 ) ^ ( n249 )  ;
assign n2140 =  ( n2134 ) ? ( n2139 ) : ( n256 ) ;
assign n2141 =  ( n2131 ) ? ( bv_1_0_n2 ) : ( n2140 ) ;
assign n2142 =  ( n1838 ) | ( n1847 )  ;
assign n2143 =  ( n2142 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n2144 =  ( n2130 ) ? ( n2141 ) : ( n2143 ) ;
assign n2145 = ~ ( n2144 ) ;
assign n2146 =  ( n1456 ) | ( n1465 )  ;
assign n2147 =  ( n1475 ) | ( n1484 )  ;
assign n2148 = ki[5:5] ;
assign n2149 =  ( n2148 ) == ( bv_1_0_n2 )  ;
assign n2150 =  ( n2149 ) | ( n1493 )  ;
assign n2151 = i_wb_data[12:12] ;
assign n2152 = ~ ( n2151 ) ;
assign n2153 = sp[12:12] ;
assign n2154 =  ( n2152 ) ^ ( n2153 )  ;
assign n2155 =  ( n2154 ) ^ ( n427 )  ;
assign n2156 =  ( n2150 ) ? ( n2155 ) : ( n434 ) ;
assign n2157 =  ( n2147 ) ? ( bv_1_0_n2 ) : ( n2156 ) ;
assign n2158 =  ( n1475 ) | ( n1484 )  ;
assign n2159 =  ( n2158 ) ? ( bv_1_0_n2 ) : ( n1875 ) ;
assign n2160 =  ( n2146 ) ? ( n2157 ) : ( n2159 ) ;
assign n2161 = ~ ( n2160 ) ;
assign n2162 =  ( n2145 ) | ( n2161 )  ;
assign n2163 =  ( n1257 ) | ( n1266 )  ;
assign n2164 =  ( n873 ) | ( n882 )  ;
assign n2165 = ki[7:7] ;
assign n2166 =  ( n2165 ) == ( bv_1_0_n2 )  ;
assign n2167 =  ( n2166 ) | ( n891 )  ;
assign n2168 = i_wb_data[10:10] ;
assign n2169 = ~ ( n2168 ) ;
assign n2170 = sp[10:10] ;
assign n2171 =  ( n2169 ) ^ ( n2170 )  ;
assign n2172 =  ( n2171 ) ^ ( n738 )  ;
assign n2173 =  ( n2167 ) ? ( n2172 ) : ( n745 ) ;
assign n2174 =  ( n2164 ) ? ( bv_1_0_n2 ) : ( n2173 ) ;
assign n2175 =  ( n873 ) | ( n882 )  ;
assign n2176 =  ( n2175 ) ? ( bv_1_0_n2 ) : ( n1892 ) ;
assign n2177 =  ( n2163 ) ? ( n2174 ) : ( n2176 ) ;
assign n2178 = ~ ( n2177 ) ;
assign n2179 =  ( n2162 ) | ( n2178 )  ;
assign n2180 =  ( n908 ) | ( n917 )  ;
assign n2181 =  ( n532 ) | ( n541 )  ;
assign n2182 = ki[9:9] ;
assign n2183 =  ( n2182 ) == ( bv_1_0_n2 )  ;
assign n2184 =  ( n2183 ) | ( n550 )  ;
assign n2185 = i_wb_data[8:8] ;
assign n2186 = ~ ( n2185 ) ;
assign n2187 = sp[8:8] ;
assign n2188 =  ( n2186 ) ^ ( n2187 )  ;
assign n2189 =  ( n2188 ) ^ ( n1054 )  ;
assign n2190 =  ( n2184 ) ? ( n2189 ) : ( n1061 ) ;
assign n2191 =  ( n2181 ) ? ( bv_1_0_n2 ) : ( n2190 ) ;
assign n2192 =  ( n532 ) | ( n541 )  ;
assign n2193 =  ( n2192 ) ? ( bv_1_0_n2 ) : ( n1909 ) ;
assign n2194 =  ( n2180 ) ? ( n2191 ) : ( n2193 ) ;
assign n2195 = ~ ( n2194 ) ;
assign n2196 =  ( n2179 ) | ( n2195 )  ;
assign n2197 = ~ ( n2196 ) ;
assign n2198 =  ( n2144 ) ^ ( n2160 )  ;
assign n2199 = ~ ( n2198 ) ;
assign n2200 =  ( n2177 ) ^ ( n2194 )  ;
assign n2201 = ~ ( n2200 ) ;
assign n2202 =  ( n2199 ) | ( n2201 )  ;
assign n2203 = ~ ( n2202 ) ;
assign n2204 =  ( n2197 ) | ( n2203 )  ;
assign n2205 =  ( n2144 ) ^ ( n2160 )  ;
assign n2206 =  ( n2205 ) ^ ( n2177 )  ;
assign n2207 =  ( n2206 ) ^ ( n2194 )  ;
assign n2208 = ~ ( n2207 ) ;
assign n2209 =  ( n567 ) | ( n576 )  ;
assign n2210 =  ( n586 ) | ( n595 )  ;
assign n2211 = ki[11:11] ;
assign n2212 =  ( n2211 ) == ( bv_1_0_n2 )  ;
assign n2213 =  ( n2212 ) | ( n604 )  ;
assign n2214 = i_wb_data[6:6] ;
assign n2215 = ~ ( n2214 ) ;
assign n2216 = sp[6:6] ;
assign n2217 =  ( n2215 ) ^ ( n2216 )  ;
assign n2218 =  ( n2217 ) ^ ( n1363 )  ;
assign n2219 =  ( n2213 ) ? ( n2218 ) : ( n1370 ) ;
assign n2220 =  ( n2210 ) ? ( bv_1_0_n2 ) : ( n2219 ) ;
assign n2221 =  ( n586 ) | ( n595 )  ;
assign n2222 =  ( n2221 ) ? ( bv_1_0_n2 ) : ( n1944 ) ;
assign n2223 =  ( n2209 ) ? ( n2220 ) : ( n2222 ) ;
assign n2224 = ~ ( n2223 ) ;
assign n2225 =  ( n2208 ) | ( n2224 )  ;
assign n2226 = ~ ( n2225 ) ;
assign n2227 =  ( n2204 ) | ( n2226 )  ;
assign n2228 = ~ ( n2227 ) ;
assign n2229 = ~ ( n2144 ) ;
assign n2230 = ~ ( n2160 ) ;
assign n2231 =  ( n2229 ) | ( n2230 )  ;
assign n2232 = ~ ( n2231 ) ;
assign n2233 = ~ ( n2177 ) ;
assign n2234 = ~ ( n2194 ) ;
assign n2235 =  ( n2233 ) | ( n2234 )  ;
assign n2236 = ~ ( n2235 ) ;
assign n2237 =  ( n2232 ) | ( n2236 )  ;
assign n2238 = ~ ( n2237 ) ;
assign n2239 =  ( n2228 ) | ( n2238 )  ;
assign n2240 =  ( n11 ) | ( n20 )  ;
assign n2241 =  ( n30 ) | ( n39 )  ;
assign n2242 = ki[13:13] ;
assign n2243 =  ( n2242 ) == ( bv_1_0_n2 )  ;
assign n2244 =  ( n2243 ) | ( n48 )  ;
assign n2245 = i_wb_data[4:4] ;
assign n2246 = ~ ( n2245 ) ;
assign n2247 = sp[4:4] ;
assign n2248 =  ( n2246 ) ^ ( n2247 )  ;
assign n2249 =  ( n2248 ) ^ ( n1989 )  ;
assign n2250 =  ( n2244 ) ? ( n2249 ) : ( n1996 ) ;
assign n2251 =  ( n2241 ) ? ( bv_1_0_n2 ) : ( n2250 ) ;
assign n2252 =  ( n30 ) | ( n39 )  ;
assign n2253 = ki[13:13] ;
assign n2254 =  ( n2253 ) == ( bv_1_0_n2 )  ;
assign n2255 =  ( n2254 ) | ( n48 )  ;
assign n2256 = i_wb_data[5:5] ;
assign n2257 = ~ ( n2256 ) ;
assign n2258 = sp[5:5] ;
assign n2259 =  ( n2257 ) ^ ( n2258 )  ;
assign n2260 =  ( n2259 ) ^ ( n241 )  ;
assign n2261 =  ( n2255 ) ? ( n2260 ) : ( n2013 ) ;
assign n2262 =  ( n2252 ) ? ( bv_1_0_n2 ) : ( n2261 ) ;
assign n2263 =  ( n2240 ) ? ( n2251 ) : ( n2262 ) ;
assign n2264 = ~ ( n2263 ) ;
assign n2265 =  ( n354 ) | ( n363 )  ;
assign n2266 =  ( n373 ) | ( n382 )  ;
assign n2267 = ki[15:15] ;
assign n2268 =  ( n2267 ) == ( bv_1_0_n2 )  ;
assign n2269 =  ( n2268 ) | ( n391 )  ;
assign n2270 = i_wb_data[2:2] ;
assign n2271 = ~ ( n2270 ) ;
assign n2272 = sp[2:2] ;
assign n2273 =  ( n2271 ) ^ ( n2272 )  ;
assign n2274 = i_wb_data[1:1] ;
assign n2275 = sp[1:1] ;
assign n2276 = ~ ( n2275 ) ;
assign n2277 =  ( n2274 ) | ( n2276 )  ;
assign n2278 = ~ ( n2277 ) ;
assign n2279 = ~ ( n237 ) ;
assign n2280 =  ( n226 ) | ( n2279 )  ;
assign n2281 = ~ ( n2280 ) ;
assign n2282 =  ( n2278 ) | ( n2281 )  ;
assign n2283 =  ( n2273 ) ^ ( n2282 )  ;
assign n2284 = i_wb_data[2:2] ;
assign n2285 = ~ ( n2284 ) ;
assign n2286 = sp[2:2] ;
assign n2287 =  ( n2285 ) ^ ( n2286 )  ;
assign n2288 =  ( n2287 ) ^ ( n2282 )  ;
assign n2289 = ~ ( n2288 ) ;
assign n2290 =  ( n2269 ) ? ( n2283 ) : ( n2289 ) ;
assign n2291 =  ( n2266 ) ? ( bv_1_0_n2 ) : ( n2290 ) ;
assign n2292 =  ( n373 ) | ( n382 )  ;
assign n2293 = ki[15:15] ;
assign n2294 =  ( n2293 ) == ( bv_1_0_n2 )  ;
assign n2295 =  ( n2294 ) | ( n391 )  ;
assign n2296 = i_wb_data[3:3] ;
assign n2297 = ~ ( n2296 ) ;
assign n2298 = sp[3:3] ;
assign n2299 =  ( n2297 ) ^ ( n2298 )  ;
assign n2300 =  ( n2299 ) ^ ( n326 )  ;
assign n2301 = i_wb_data[3:3] ;
assign n2302 = ~ ( n2301 ) ;
assign n2303 = sp[3:3] ;
assign n2304 =  ( n2302 ) ^ ( n2303 )  ;
assign n2305 =  ( n2304 ) ^ ( n326 )  ;
assign n2306 = ~ ( n2305 ) ;
assign n2307 =  ( n2295 ) ? ( n2300 ) : ( n2306 ) ;
assign n2308 =  ( n2292 ) ? ( bv_1_0_n2 ) : ( n2307 ) ;
assign n2309 =  ( n2265 ) ? ( n2291 ) : ( n2308 ) ;
assign n2310 = ~ ( n2309 ) ;
assign n2311 =  ( n2264 ) | ( n2310 )  ;
assign n2312 = ~ ( n2311 ) ;
assign n2313 =  ( n2263 ) ^ ( n2309 )  ;
assign n2314 =  ( n2312 ) | ( n2313 )  ;
assign n2315 = ~ ( n2314 ) ;
assign n2316 =  ( n2239 ) | ( n2315 )  ;
assign n2317 =  ( n1838 ) | ( n1847 )  ;
assign n2318 =  ( n2317 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n2319 = ~ ( n2318 ) ;
assign n2320 =  ( n2319 ) ^ ( n1879 )  ;
assign n2321 =  ( n2320 ) ^ ( n1896 )  ;
assign n2322 =  ( n2321 ) ^ ( n1913 )  ;
assign n2323 =  ( n2322 ) ^ ( n1948 )  ;
assign n2324 = ~ ( n2323 ) ;
assign n2325 =  ( n2316 ) | ( n2324 )  ;
assign n2326 = ~ ( n2325 ) ;
assign n2327 =  ( n2227 ) ^ ( n2237 )  ;
assign n2328 = ~ ( n2327 ) ;
assign n2329 =  ( n1838 ) | ( n1847 )  ;
assign n2330 =  ( n2329 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n2331 = ~ ( n2330 ) ;
assign n2332 =  ( n2314 ) ^ ( n2331 )  ;
assign n2333 =  ( n2332 ) ^ ( n1879 )  ;
assign n2334 =  ( n2333 ) ^ ( n1896 )  ;
assign n2335 =  ( n2334 ) ^ ( n1913 )  ;
assign n2336 =  ( n2335 ) ^ ( n1948 )  ;
assign n2337 = ~ ( n2336 ) ;
assign n2338 =  ( n2328 ) | ( n2337 )  ;
assign n2339 = ~ ( n2338 ) ;
assign n2340 =  ( n2326 ) | ( n2339 )  ;
assign n2341 =  ( n2227 ) ^ ( n2237 )  ;
assign n2342 =  ( n2341 ) ^ ( n2314 )  ;
assign n2343 =  ( n1838 ) | ( n1847 )  ;
assign n2344 =  ( n2343 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n2345 = ~ ( n2344 ) ;
assign n2346 =  ( n2342 ) ^ ( n2345 )  ;
assign n2347 =  ( n2346 ) ^ ( n1879 )  ;
assign n2348 =  ( n2347 ) ^ ( n1896 )  ;
assign n2349 =  ( n2348 ) ^ ( n1913 )  ;
assign n2350 =  ( n2349 ) ^ ( n1948 )  ;
assign n2351 = ~ ( n2350 ) ;
assign n2352 =  ( n11 ) | ( n20 )  ;
assign n2353 =  ( n30 ) | ( n39 )  ;
assign n2354 =  ( n2353 ) ? ( bv_1_0_n2 ) : ( n2261 ) ;
assign n2355 =  ( n30 ) | ( n39 )  ;
assign n2356 =  ( n2355 ) ? ( bv_1_0_n2 ) : ( n1615 ) ;
assign n2357 =  ( n2352 ) ? ( n2354 ) : ( n2356 ) ;
assign n2358 = ~ ( n2357 ) ;
assign n2359 =  ( n2351 ) | ( n2358 )  ;
assign n2360 = ~ ( n2359 ) ;
assign n2361 =  ( n2340 ) | ( n2360 )  ;
assign n2362 = ~ ( n2361 ) ;
assign n2363 = ~ ( n2227 ) ;
assign n2364 = ~ ( n2237 ) ;
assign n2365 =  ( n2363 ) | ( n2364 )  ;
assign n2366 = ~ ( n2365 ) ;
assign n2367 = ~ ( n2314 ) ;
assign n2368 = ~ ( n2323 ) ;
assign n2369 =  ( n2367 ) | ( n2368 )  ;
assign n2370 = ~ ( n2369 ) ;
assign n2371 =  ( n2366 ) | ( n2370 )  ;
assign n2372 = ~ ( n2371 ) ;
assign n2373 =  ( n2362 ) | ( n2372 )  ;
assign n2374 = ~ ( n2373 ) ;
assign n2375 =  ( n2361 ) ^ ( n2371 )  ;
assign n2376 = ~ ( n2375 ) ;
assign n2377 =  ( bv_1_1_n5 ) ^ ( n1952 )  ;
assign n2378 =  ( n2377 ) ^ ( n1963 )  ;
assign n2379 =  ( n2378 ) ^ ( n1513 )  ;
assign n2380 =  ( n2379 ) ^ ( n1538 )  ;
assign n2381 =  ( n2380 ) ^ ( n1564 )  ;
assign n2382 =  ( n2381 ) ^ ( n1590 )  ;
assign n2383 =  ( n2382 ) ^ ( n1628 )  ;
assign n2384 =  ( n2383 ) ^ ( n2016 )  ;
assign n2385 = ~ ( n2384 ) ;
assign n2386 =  ( n2376 ) | ( n2385 )  ;
assign n2387 = ~ ( n2386 ) ;
assign n2388 =  ( n2374 ) | ( n2387 )  ;
assign n2389 = ~ ( n2388 ) ;
assign n2390 =  ( n2038 ) ^ ( n2052 )  ;
assign n2391 =  ( n2390 ) ^ ( n1632 )  ;
assign n2392 =  ( n2391 ) ^ ( n1642 )  ;
assign n2393 =  ( n1475 ) | ( n1484 )  ;
assign n2394 =  ( n2393 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n2395 = ~ ( n2394 ) ;
assign n2396 =  ( n2392 ) ^ ( n2395 )  ;
assign n2397 =  ( n2396 ) ^ ( n1656 )  ;
assign n2398 =  ( n2397 ) ^ ( n1663 )  ;
assign n2399 =  ( n2398 ) ^ ( n1670 )  ;
assign n2400 =  ( n2399 ) ^ ( n1677 )  ;
assign n2401 = ~ ( n2400 ) ;
assign n2402 =  ( n2389 ) | ( n2401 )  ;
assign n2403 = ~ ( n2402 ) ;
assign n2404 =  ( n2388 ) ^ ( n2038 )  ;
assign n2405 =  ( n2404 ) ^ ( n2052 )  ;
assign n2406 =  ( n2405 ) ^ ( n1632 )  ;
assign n2407 =  ( n2406 ) ^ ( n1642 )  ;
assign n2408 =  ( n1475 ) | ( n1484 )  ;
assign n2409 =  ( n2408 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n2410 = ~ ( n2409 ) ;
assign n2411 =  ( n2407 ) ^ ( n2410 )  ;
assign n2412 =  ( n2411 ) ^ ( n1656 )  ;
assign n2413 =  ( n2412 ) ^ ( n1663 )  ;
assign n2414 =  ( n2413 ) ^ ( n1670 )  ;
assign n2415 =  ( n2414 ) ^ ( n1677 )  ;
assign n2416 = ~ ( n2415 ) ;
assign n2417 =  ( n354 ) | ( n363 )  ;
assign n2418 =  ( n373 ) | ( n382 )  ;
assign n2419 =  ( n2418 ) ? ( bv_1_0_n2 ) : ( n2014 ) ;
assign n2420 =  ( n373 ) | ( n382 )  ;
assign n2421 =  ( n2420 ) ? ( bv_1_0_n2 ) : ( n1371 ) ;
assign n2422 =  ( n2417 ) ? ( n2419 ) : ( n2421 ) ;
assign n2423 = ~ ( n2422 ) ;
assign n2424 =  ( n2416 ) | ( n2423 )  ;
assign n2425 = ~ ( n2424 ) ;
assign n2426 =  ( n2403 ) | ( n2425 )  ;
assign n2427 = ~ ( n2426 ) ;
assign n2428 =  ( n2111 ) | ( n2427 )  ;
assign n2429 =  ( bv_1_1_n5 ) ^ ( n2070 )  ;
assign n2430 =  ( n2429 ) ^ ( n1682 )  ;
assign n2431 =  ( n2430 ) ^ ( n1713 )  ;
assign n2432 =  ( n2431 ) ^ ( n1723 )  ;
assign n2433 =  ( n2432 ) ^ ( n1281 )  ;
assign n2434 =  ( n2433 ) ^ ( n1297 )  ;
assign n2435 =  ( n2434 ) ^ ( n1314 )  ;
assign n2436 =  ( n2435 ) ^ ( n1331 )  ;
assign n2437 =  ( n2436 ) ^ ( n1375 )  ;
assign n2438 = ~ ( n2437 ) ;
assign n2439 =  ( n2428 ) | ( n2438 )  ;
assign n2440 = ~ ( n2439 ) ;
assign n2441 =  ( n2095 ) | ( n2440 )  ;
assign n2442 = ~ ( n2110 ) ;
assign n2443 =  ( bv_1_1_n5 ) ^ ( n2426 )  ;
assign n2444 =  ( n2443 ) ^ ( n2070 )  ;
assign n2445 =  ( n2444 ) ^ ( n1682 )  ;
assign n2446 =  ( n2445 ) ^ ( n1713 )  ;
assign n2447 =  ( n2446 ) ^ ( n1723 )  ;
assign n2448 =  ( n2447 ) ^ ( n1281 )  ;
assign n2449 =  ( n2448 ) ^ ( n1297 )  ;
assign n2450 =  ( n2449 ) ^ ( n1314 )  ;
assign n2451 =  ( n2450 ) ^ ( n1331 )  ;
assign n2452 =  ( n2451 ) ^ ( n1375 )  ;
assign n2453 = ~ ( n2452 ) ;
assign n2454 =  ( n2442 ) | ( n2453 )  ;
assign n2455 = ki[1:1] ;
assign n2456 =  ( n2455 ) == ( bv_1_1_n5 )  ;
assign n2457 = ki[0:0] ;
assign n2458 =  ( n2457 ) == ( bv_1_1_n5 )  ;
assign n2459 =  ( n2456 ) | ( n2458 )  ;
assign n2460 = ki[1:1] ;
assign n2461 =  ( n2460 ) == ( bv_1_1_n5 )  ;
assign n2462 = i_wb_data[15:15] ;
assign n2463 = ~ ( n2462 ) ;
assign n2464 = sp[15:15] ;
assign n2465 =  ( n2463 ) ^ ( n2464 )  ;
assign n2466 =  ( n2465 ) ^ ( n334 )  ;
assign n2467 =  ( n2461 ) ? ( n341 ) : ( n2466 ) ;
assign n2468 =  ( n2459 ) ? ( n2467 ) : ( bv_1_0_n2 ) ;
assign n2469 =  ( n2120 ) | ( n2129 )  ;
assign n2470 =  ( n1838 ) | ( n1847 )  ;
assign n2471 = ki[3:3] ;
assign n2472 =  ( n2471 ) == ( bv_1_0_n2 )  ;
assign n2473 =  ( n2472 ) | ( n1856 )  ;
assign n2474 = i_wb_data[13:13] ;
assign n2475 = ~ ( n2474 ) ;
assign n2476 = sp[13:13] ;
assign n2477 =  ( n2475 ) ^ ( n2476 )  ;
assign n2478 =  ( n2477 ) ^ ( n245 )  ;
assign n2479 =  ( n2473 ) ? ( n2478 ) : ( n451 ) ;
assign n2480 =  ( n2470 ) ? ( bv_1_0_n2 ) : ( n2479 ) ;
assign n2481 =  ( n1838 ) | ( n1847 )  ;
assign n2482 =  ( n2481 ) ? ( bv_1_0_n2 ) : ( n2140 ) ;
assign n2483 =  ( n2469 ) ? ( n2480 ) : ( n2482 ) ;
assign n2484 = ~ ( n2483 ) ;
assign n2485 =  ( n2468 ) | ( n2484 )  ;
assign n2486 =  ( n1456 ) | ( n1465 )  ;
assign n2487 =  ( n1475 ) | ( n1484 )  ;
assign n2488 = ki[5:5] ;
assign n2489 =  ( n2488 ) == ( bv_1_0_n2 )  ;
assign n2490 =  ( n2489 ) | ( n1493 )  ;
assign n2491 = i_wb_data[11:11] ;
assign n2492 = ~ ( n2491 ) ;
assign n2493 = sp[11:11] ;
assign n2494 =  ( n2492 ) ^ ( n2493 )  ;
assign n2495 =  ( n2494 ) ^ ( n423 )  ;
assign n2496 =  ( n2490 ) ? ( n2495 ) : ( n648 ) ;
assign n2497 =  ( n2487 ) ? ( bv_1_0_n2 ) : ( n2496 ) ;
assign n2498 =  ( n1475 ) | ( n1484 )  ;
assign n2499 =  ( n2498 ) ? ( bv_1_0_n2 ) : ( n2156 ) ;
assign n2500 =  ( n2486 ) ? ( n2497 ) : ( n2499 ) ;
assign n2501 = ~ ( n2500 ) ;
assign n2502 =  ( n2485 ) | ( n2501 )  ;
assign n2503 =  ( n1257 ) | ( n1266 )  ;
assign n2504 =  ( n873 ) | ( n882 )  ;
assign n2505 = ki[7:7] ;
assign n2506 =  ( n2505 ) == ( bv_1_0_n2 )  ;
assign n2507 =  ( n2506 ) | ( n891 )  ;
assign n2508 = i_wb_data[9:9] ;
assign n2509 = ~ ( n2508 ) ;
assign n2510 = sp[9:9] ;
assign n2511 =  ( n2509 ) ^ ( n2510 )  ;
assign n2512 =  ( n2511 ) ^ ( n734 )  ;
assign n2513 =  ( n2507 ) ? ( n2512 ) : ( n985 ) ;
assign n2514 =  ( n2504 ) ? ( bv_1_0_n2 ) : ( n2513 ) ;
assign n2515 =  ( n873 ) | ( n882 )  ;
assign n2516 =  ( n2515 ) ? ( bv_1_0_n2 ) : ( n2173 ) ;
assign n2517 =  ( n2503 ) ? ( n2514 ) : ( n2516 ) ;
assign n2518 = ~ ( n2517 ) ;
assign n2519 =  ( n2502 ) | ( n2518 )  ;
assign n2520 = ~ ( n2519 ) ;
assign n2521 = ~ ( n2468 ) ;
assign n2522 =  ( n2521 ) ^ ( n2483 )  ;
assign n2523 = ~ ( n2522 ) ;
assign n2524 =  ( n2500 ) ^ ( n2517 )  ;
assign n2525 = ~ ( n2524 ) ;
assign n2526 =  ( n2523 ) | ( n2525 )  ;
assign n2527 = ~ ( n2526 ) ;
assign n2528 =  ( n2520 ) | ( n2527 )  ;
assign n2529 = ~ ( n2468 ) ;
assign n2530 =  ( n2529 ) ^ ( n2483 )  ;
assign n2531 =  ( n2530 ) ^ ( n2500 )  ;
assign n2532 =  ( n2531 ) ^ ( n2517 )  ;
assign n2533 = ~ ( n2532 ) ;
assign n2534 =  ( n908 ) | ( n917 )  ;
assign n2535 =  ( n532 ) | ( n541 )  ;
assign n2536 = ki[9:9] ;
assign n2537 =  ( n2536 ) == ( bv_1_0_n2 )  ;
assign n2538 =  ( n2537 ) | ( n550 )  ;
assign n2539 = i_wb_data[7:7] ;
assign n2540 = ~ ( n2539 ) ;
assign n2541 = sp[7:7] ;
assign n2542 =  ( n2540 ) ^ ( n2541 )  ;
assign n2543 =  ( n2542 ) ^ ( n330 )  ;
assign n2544 =  ( n2538 ) ? ( n2543 ) : ( n1035 ) ;
assign n2545 =  ( n2535 ) ? ( bv_1_0_n2 ) : ( n2544 ) ;
assign n2546 =  ( n532 ) | ( n541 )  ;
assign n2547 =  ( n2546 ) ? ( bv_1_0_n2 ) : ( n2190 ) ;
assign n2548 =  ( n2534 ) ? ( n2545 ) : ( n2547 ) ;
assign n2549 = ~ ( n2548 ) ;
assign n2550 =  ( n2533 ) | ( n2549 )  ;
assign n2551 = ~ ( n2550 ) ;
assign n2552 =  ( n2528 ) | ( n2551 )  ;
assign n2553 = ~ ( n2552 ) ;
assign n2554 = ~ ( n2483 ) ;
assign n2555 =  ( n2468 ) | ( n2554 )  ;
assign n2556 = ~ ( n2555 ) ;
assign n2557 = ~ ( n2500 ) ;
assign n2558 = ~ ( n2517 ) ;
assign n2559 =  ( n2557 ) | ( n2558 )  ;
assign n2560 = ~ ( n2559 ) ;
assign n2561 =  ( n2556 ) | ( n2560 )  ;
assign n2562 = ~ ( n2561 ) ;
assign n2563 =  ( n2553 ) | ( n2562 )  ;
assign n2564 =  ( n567 ) | ( n576 )  ;
assign n2565 =  ( n586 ) | ( n595 )  ;
assign n2566 = ki[11:11] ;
assign n2567 =  ( n2566 ) == ( bv_1_0_n2 )  ;
assign n2568 =  ( n2567 ) | ( n604 )  ;
assign n2569 = i_wb_data[5:5] ;
assign n2570 = ~ ( n2569 ) ;
assign n2571 = sp[5:5] ;
assign n2572 =  ( n2570 ) ^ ( n2571 )  ;
assign n2573 =  ( n2572 ) ^ ( n241 )  ;
assign n2574 =  ( n2568 ) ? ( n2573 ) : ( n2013 ) ;
assign n2575 =  ( n2565 ) ? ( bv_1_0_n2 ) : ( n2574 ) ;
assign n2576 =  ( n586 ) | ( n595 )  ;
assign n2577 =  ( n2576 ) ? ( bv_1_0_n2 ) : ( n2219 ) ;
assign n2578 =  ( n2564 ) ? ( n2575 ) : ( n2577 ) ;
assign n2579 = ~ ( n2578 ) ;
assign n2580 =  ( n11 ) | ( n20 )  ;
assign n2581 =  ( n30 ) | ( n39 )  ;
assign n2582 = ki[13:13] ;
assign n2583 =  ( n2582 ) == ( bv_1_0_n2 )  ;
assign n2584 =  ( n2583 ) | ( n48 )  ;
assign n2585 = i_wb_data[3:3] ;
assign n2586 = ~ ( n2585 ) ;
assign n2587 = sp[3:3] ;
assign n2588 =  ( n2586 ) ^ ( n2587 )  ;
assign n2589 =  ( n2588 ) ^ ( n326 )  ;
assign n2590 =  ( n2584 ) ? ( n2589 ) : ( n2306 ) ;
assign n2591 =  ( n2581 ) ? ( bv_1_0_n2 ) : ( n2590 ) ;
assign n2592 =  ( n30 ) | ( n39 )  ;
assign n2593 =  ( n2592 ) ? ( bv_1_0_n2 ) : ( n2250 ) ;
assign n2594 =  ( n2580 ) ? ( n2591 ) : ( n2593 ) ;
assign n2595 = ~ ( n2594 ) ;
assign n2596 =  ( n2579 ) | ( n2595 )  ;
assign n2597 = ~ ( n2596 ) ;
assign n2598 =  ( n2578 ) ^ ( n2594 )  ;
assign n2599 = ~ ( n2598 ) ;
assign n2600 =  ( n354 ) | ( n363 )  ;
assign n2601 =  ( n373 ) | ( n382 )  ;
assign n2602 = ki[15:15] ;
assign n2603 =  ( n2602 ) == ( bv_1_0_n2 )  ;
assign n2604 =  ( n2603 ) | ( n391 )  ;
assign n2605 = i_wb_data[1:1] ;
assign n2606 = ~ ( n2605 ) ;
assign n2607 = sp[1:1] ;
assign n2608 =  ( n2606 ) ^ ( n2607 )  ;
assign n2609 =  ( n2608 ) ^ ( n237 )  ;
assign n2610 = i_wb_data[1:1] ;
assign n2611 = ~ ( n2610 ) ;
assign n2612 = sp[1:1] ;
assign n2613 =  ( n2611 ) ^ ( n2612 )  ;
assign n2614 =  ( n2613 ) ^ ( n237 )  ;
assign n2615 = ~ ( n2614 ) ;
assign n2616 =  ( n2604 ) ? ( n2609 ) : ( n2615 ) ;
assign n2617 =  ( n2601 ) ? ( bv_1_0_n2 ) : ( n2616 ) ;
assign n2618 =  ( n373 ) | ( n382 )  ;
assign n2619 =  ( n2618 ) ? ( bv_1_0_n2 ) : ( n2290 ) ;
assign n2620 =  ( n2600 ) ? ( n2617 ) : ( n2619 ) ;
assign n2621 = ~ ( n2620 ) ;
assign n2622 =  ( n2599 ) | ( n2621 )  ;
assign n2623 = ~ ( n2622 ) ;
assign n2624 =  ( n2597 ) | ( n2623 )  ;
assign n2625 = ~ ( n2624 ) ;
assign n2626 =  ( n2563 ) | ( n2625 )  ;
assign n2627 =  ( n2144 ) ^ ( n2160 )  ;
assign n2628 =  ( n2627 ) ^ ( n2177 )  ;
assign n2629 =  ( n2628 ) ^ ( n2194 )  ;
assign n2630 =  ( n2629 ) ^ ( n2223 )  ;
assign n2631 = ~ ( n2630 ) ;
assign n2632 =  ( n2626 ) | ( n2631 )  ;
assign n2633 = ~ ( n2632 ) ;
assign n2634 =  ( n2552 ) ^ ( n2561 )  ;
assign n2635 = ~ ( n2634 ) ;
assign n2636 =  ( n2624 ) ^ ( n2144 )  ;
assign n2637 =  ( n2636 ) ^ ( n2160 )  ;
assign n2638 =  ( n2637 ) ^ ( n2177 )  ;
assign n2639 =  ( n2638 ) ^ ( n2194 )  ;
assign n2640 =  ( n2639 ) ^ ( n2223 )  ;
assign n2641 = ~ ( n2640 ) ;
assign n2642 =  ( n2635 ) | ( n2641 )  ;
assign n2643 = ~ ( n2642 ) ;
assign n2644 =  ( n2633 ) | ( n2643 )  ;
assign n2645 =  ( n2552 ) ^ ( n2561 )  ;
assign n2646 =  ( n2645 ) ^ ( n2624 )  ;
assign n2647 =  ( n2646 ) ^ ( n2144 )  ;
assign n2648 =  ( n2647 ) ^ ( n2160 )  ;
assign n2649 =  ( n2648 ) ^ ( n2177 )  ;
assign n2650 =  ( n2649 ) ^ ( n2194 )  ;
assign n2651 =  ( n2650 ) ^ ( n2223 )  ;
assign n2652 = ~ ( n2651 ) ;
assign n2653 =  ( bv_1_1_n5 ) ^ ( n2263 )  ;
assign n2654 =  ( n2653 ) ^ ( n2309 )  ;
assign n2655 = ~ ( n2654 ) ;
assign n2656 =  ( n2652 ) | ( n2655 )  ;
assign n2657 = ~ ( n2656 ) ;
assign n2658 =  ( n2644 ) | ( n2657 )  ;
assign n2659 = ~ ( n2658 ) ;
assign n2660 = ~ ( n2552 ) ;
assign n2661 = ~ ( n2561 ) ;
assign n2662 =  ( n2660 ) | ( n2661 )  ;
assign n2663 = ~ ( n2662 ) ;
assign n2664 = ~ ( n2624 ) ;
assign n2665 =  ( n2144 ) ^ ( n2160 )  ;
assign n2666 =  ( n2665 ) ^ ( n2177 )  ;
assign n2667 =  ( n2666 ) ^ ( n2194 )  ;
assign n2668 =  ( n2667 ) ^ ( n2223 )  ;
assign n2669 = ~ ( n2668 ) ;
assign n2670 =  ( n2664 ) | ( n2669 )  ;
assign n2671 = ~ ( n2670 ) ;
assign n2672 =  ( n2663 ) | ( n2671 )  ;
assign n2673 = ~ ( n2672 ) ;
assign n2674 =  ( n2659 ) | ( n2673 )  ;
assign n2675 = ~ ( n2674 ) ;
assign n2676 =  ( n2633 ) | ( n2643 )  ;
assign n2677 =  ( n2676 ) | ( n2657 )  ;
assign n2678 =  ( n2677 ) ^ ( n2672 )  ;
assign n2679 = ~ ( n2678 ) ;
assign n2680 =  ( n2227 ) ^ ( n2237 )  ;
assign n2681 =  ( n2680 ) ^ ( n2314 )  ;
assign n2682 =  ( n1838 ) | ( n1847 )  ;
assign n2683 =  ( n2682 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n2684 = ~ ( n2683 ) ;
assign n2685 =  ( n2681 ) ^ ( n2684 )  ;
assign n2686 =  ( n2685 ) ^ ( n1879 )  ;
assign n2687 =  ( n2686 ) ^ ( n1896 )  ;
assign n2688 =  ( n2687 ) ^ ( n1913 )  ;
assign n2689 =  ( n2688 ) ^ ( n1948 )  ;
assign n2690 =  ( n2689 ) ^ ( n2357 )  ;
assign n2691 = ~ ( n2690 ) ;
assign n2692 =  ( n2679 ) | ( n2691 )  ;
assign n2693 = ~ ( n2692 ) ;
assign n2694 =  ( n2675 ) | ( n2693 )  ;
assign n2695 = ~ ( n2694 ) ;
assign n2696 =  ( bv_1_1_n5 ) ^ ( n2361 )  ;
assign n2697 =  ( n2696 ) ^ ( n2371 )  ;
assign n2698 =  ( n2697 ) ^ ( n1952 )  ;
assign n2699 =  ( n2698 ) ^ ( n1963 )  ;
assign n2700 =  ( n2699 ) ^ ( n1513 )  ;
assign n2701 =  ( n2700 ) ^ ( n1538 )  ;
assign n2702 =  ( n2701 ) ^ ( n1564 )  ;
assign n2703 =  ( n2702 ) ^ ( n1590 )  ;
assign n2704 =  ( n2703 ) ^ ( n1628 )  ;
assign n2705 =  ( n2704 ) ^ ( n2016 )  ;
assign n2706 = ~ ( n2705 ) ;
assign n2707 =  ( n2695 ) | ( n2706 )  ;
assign n2708 =  ( n2388 ) ^ ( n2038 )  ;
assign n2709 =  ( n2708 ) ^ ( n2052 )  ;
assign n2710 =  ( n2709 ) ^ ( n1632 )  ;
assign n2711 =  ( n2710 ) ^ ( n1642 )  ;
assign n2712 =  ( n1475 ) | ( n1484 )  ;
assign n2713 =  ( n2712 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n2714 = ~ ( n2713 ) ;
assign n2715 =  ( n2711 ) ^ ( n2714 )  ;
assign n2716 =  ( n2715 ) ^ ( n1656 )  ;
assign n2717 =  ( n2716 ) ^ ( n1663 )  ;
assign n2718 =  ( n2717 ) ^ ( n1670 )  ;
assign n2719 =  ( n2718 ) ^ ( n1677 )  ;
assign n2720 =  ( n2719 ) ^ ( n2422 )  ;
assign n2721 = ~ ( n2720 ) ;
assign n2722 =  ( n2707 ) | ( n2721 )  ;
assign n2723 = ~ ( n2722 ) ;
assign n2724 = ~ ( n2692 ) ;
assign n2725 =  ( n2675 ) | ( n2724 )  ;
assign n2726 = ~ ( n2725 ) ;
assign n2727 =  ( n2726 ) | ( n2706 )  ;
assign n2728 = ~ ( n2727 ) ;
assign n2729 =  ( n2728 ) ^ ( n2388 )  ;
assign n2730 =  ( n2729 ) ^ ( n2038 )  ;
assign n2731 =  ( n2730 ) ^ ( n2052 )  ;
assign n2732 =  ( n2731 ) ^ ( n1632 )  ;
assign n2733 =  ( n2732 ) ^ ( n1642 )  ;
assign n2734 =  ( n1475 ) | ( n1484 )  ;
assign n2735 =  ( n2734 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n2736 = ~ ( n2735 ) ;
assign n2737 =  ( n2733 ) ^ ( n2736 )  ;
assign n2738 =  ( n2737 ) ^ ( n1656 )  ;
assign n2739 =  ( n2738 ) ^ ( n1663 )  ;
assign n2740 =  ( n2739 ) ^ ( n1670 )  ;
assign n2741 =  ( n2740 ) ^ ( n1677 )  ;
assign n2742 =  ( n2741 ) ^ ( n2422 )  ;
assign n2743 = ~ ( n2742 ) ;
assign n2744 = ki[0:0] ;
assign n2745 =  ( n2744 ) == ( bv_1_1_n5 )  ;
assign n2746 = ki[1:1] ;
assign n2747 =  ( n2746 ) == ( bv_1_0_n2 )  ;
assign n2748 =  ( n2745 ) | ( n2747 )  ;
assign n2749 = ki[1:1] ;
assign n2750 =  ( n2749 ) == ( bv_1_1_n5 )  ;
assign n2751 = ki[0:0] ;
assign n2752 =  ( n2751 ) == ( bv_1_1_n5 )  ;
assign n2753 =  ( n2750 ) | ( n2752 )  ;
assign n2754 = ki[1:1] ;
assign n2755 =  ( n2754 ) == ( bv_1_1_n5 )  ;
assign n2756 = i_wb_data[14:14] ;
assign n2757 = ~ ( n2756 ) ;
assign n2758 = sp[14:14] ;
assign n2759 =  ( n2757 ) ^ ( n2758 )  ;
assign n2760 =  ( n2759 ) ^ ( n249 )  ;
assign n2761 =  ( n2755 ) ? ( n256 ) : ( n2760 ) ;
assign n2762 =  ( n2753 ) ? ( n2761 ) : ( bv_1_0_n2 ) ;
assign n2763 =  ( n2748 ) ? ( n2468 ) : ( n2762 ) ;
assign n2764 = ~ ( n2763 ) ;
assign n2765 =  ( n2120 ) | ( n2129 )  ;
assign n2766 =  ( n1838 ) | ( n1847 )  ;
assign n2767 = ki[3:3] ;
assign n2768 =  ( n2767 ) == ( bv_1_0_n2 )  ;
assign n2769 =  ( n2768 ) | ( n1856 )  ;
assign n2770 = i_wb_data[12:12] ;
assign n2771 = ~ ( n2770 ) ;
assign n2772 = sp[12:12] ;
assign n2773 =  ( n2771 ) ^ ( n2772 )  ;
assign n2774 =  ( n2773 ) ^ ( n427 )  ;
assign n2775 =  ( n2769 ) ? ( n2774 ) : ( n434 ) ;
assign n2776 =  ( n2766 ) ? ( bv_1_0_n2 ) : ( n2775 ) ;
assign n2777 =  ( n1838 ) | ( n1847 )  ;
assign n2778 =  ( n2777 ) ? ( bv_1_0_n2 ) : ( n2479 ) ;
assign n2779 =  ( n2765 ) ? ( n2776 ) : ( n2778 ) ;
assign n2780 = ~ ( n2779 ) ;
assign n2781 =  ( n2764 ) | ( n2780 )  ;
assign n2782 =  ( n1456 ) | ( n1465 )  ;
assign n2783 =  ( n1475 ) | ( n1484 )  ;
assign n2784 = ki[5:5] ;
assign n2785 =  ( n2784 ) == ( bv_1_0_n2 )  ;
assign n2786 =  ( n2785 ) | ( n1493 )  ;
assign n2787 = i_wb_data[10:10] ;
assign n2788 = ~ ( n2787 ) ;
assign n2789 = sp[10:10] ;
assign n2790 =  ( n2788 ) ^ ( n2789 )  ;
assign n2791 =  ( n2790 ) ^ ( n738 )  ;
assign n2792 =  ( n2786 ) ? ( n2791 ) : ( n745 ) ;
assign n2793 =  ( n2783 ) ? ( bv_1_0_n2 ) : ( n2792 ) ;
assign n2794 =  ( n1475 ) | ( n1484 )  ;
assign n2795 =  ( n2794 ) ? ( bv_1_0_n2 ) : ( n2496 ) ;
assign n2796 =  ( n2782 ) ? ( n2793 ) : ( n2795 ) ;
assign n2797 = ~ ( n2796 ) ;
assign n2798 =  ( n2781 ) | ( n2797 )  ;
assign n2799 =  ( n1257 ) | ( n1266 )  ;
assign n2800 =  ( n873 ) | ( n882 )  ;
assign n2801 = ki[7:7] ;
assign n2802 =  ( n2801 ) == ( bv_1_0_n2 )  ;
assign n2803 =  ( n2802 ) | ( n891 )  ;
assign n2804 = i_wb_data[8:8] ;
assign n2805 = ~ ( n2804 ) ;
assign n2806 = sp[8:8] ;
assign n2807 =  ( n2805 ) ^ ( n2806 )  ;
assign n2808 =  ( n2807 ) ^ ( n1054 )  ;
assign n2809 =  ( n2803 ) ? ( n2808 ) : ( n1061 ) ;
assign n2810 =  ( n2800 ) ? ( bv_1_0_n2 ) : ( n2809 ) ;
assign n2811 =  ( n873 ) | ( n882 )  ;
assign n2812 =  ( n2811 ) ? ( bv_1_0_n2 ) : ( n2513 ) ;
assign n2813 =  ( n2799 ) ? ( n2810 ) : ( n2812 ) ;
assign n2814 = ~ ( n2813 ) ;
assign n2815 =  ( n2798 ) | ( n2814 )  ;
assign n2816 = ~ ( n2815 ) ;
assign n2817 =  ( n2763 ) ^ ( n2779 )  ;
assign n2818 = ~ ( n2817 ) ;
assign n2819 =  ( n2796 ) ^ ( n2813 )  ;
assign n2820 = ~ ( n2819 ) ;
assign n2821 =  ( n2818 ) | ( n2820 )  ;
assign n2822 = ~ ( n2821 ) ;
assign n2823 =  ( n2816 ) | ( n2822 )  ;
assign n2824 =  ( n2763 ) ^ ( n2779 )  ;
assign n2825 =  ( n2824 ) ^ ( n2796 )  ;
assign n2826 =  ( n2825 ) ^ ( n2813 )  ;
assign n2827 = ~ ( n2826 ) ;
assign n2828 =  ( n908 ) | ( n917 )  ;
assign n2829 =  ( n532 ) | ( n541 )  ;
assign n2830 = ki[9:9] ;
assign n2831 =  ( n2830 ) == ( bv_1_0_n2 )  ;
assign n2832 =  ( n2831 ) | ( n550 )  ;
assign n2833 = i_wb_data[6:6] ;
assign n2834 = ~ ( n2833 ) ;
assign n2835 = sp[6:6] ;
assign n2836 =  ( n2834 ) ^ ( n2835 )  ;
assign n2837 =  ( n2836 ) ^ ( n1363 )  ;
assign n2838 =  ( n2832 ) ? ( n2837 ) : ( n1370 ) ;
assign n2839 =  ( n2829 ) ? ( bv_1_0_n2 ) : ( n2838 ) ;
assign n2840 =  ( n532 ) | ( n541 )  ;
assign n2841 =  ( n2840 ) ? ( bv_1_0_n2 ) : ( n2544 ) ;
assign n2842 =  ( n2828 ) ? ( n2839 ) : ( n2841 ) ;
assign n2843 = ~ ( n2842 ) ;
assign n2844 =  ( n2827 ) | ( n2843 )  ;
assign n2845 = ~ ( n2844 ) ;
assign n2846 =  ( n2823 ) | ( n2845 )  ;
assign n2847 = ~ ( n2846 ) ;
assign n2848 = ~ ( n2763 ) ;
assign n2849 = ~ ( n2779 ) ;
assign n2850 =  ( n2848 ) | ( n2849 )  ;
assign n2851 = ~ ( n2850 ) ;
assign n2852 = ~ ( n2796 ) ;
assign n2853 = ~ ( n2813 ) ;
assign n2854 =  ( n2852 ) | ( n2853 )  ;
assign n2855 = ~ ( n2854 ) ;
assign n2856 =  ( n2851 ) | ( n2855 )  ;
assign n2857 = ~ ( n2856 ) ;
assign n2858 =  ( n2847 ) | ( n2857 )  ;
assign n2859 =  ( n567 ) | ( n576 )  ;
assign n2860 =  ( n586 ) | ( n595 )  ;
assign n2861 = ki[11:11] ;
assign n2862 =  ( n2861 ) == ( bv_1_0_n2 )  ;
assign n2863 =  ( n2862 ) | ( n604 )  ;
assign n2864 = i_wb_data[4:4] ;
assign n2865 = ~ ( n2864 ) ;
assign n2866 = sp[4:4] ;
assign n2867 =  ( n2865 ) ^ ( n2866 )  ;
assign n2868 =  ( n2867 ) ^ ( n1989 )  ;
assign n2869 =  ( n2863 ) ? ( n2868 ) : ( n1996 ) ;
assign n2870 =  ( n2860 ) ? ( bv_1_0_n2 ) : ( n2869 ) ;
assign n2871 =  ( n586 ) | ( n595 )  ;
assign n2872 =  ( n2871 ) ? ( bv_1_0_n2 ) : ( n2574 ) ;
assign n2873 =  ( n2859 ) ? ( n2870 ) : ( n2872 ) ;
assign n2874 = ~ ( n2873 ) ;
assign n2875 =  ( n11 ) | ( n20 )  ;
assign n2876 =  ( n30 ) | ( n39 )  ;
assign n2877 = ki[13:13] ;
assign n2878 =  ( n2877 ) == ( bv_1_0_n2 )  ;
assign n2879 =  ( n2878 ) | ( n48 )  ;
assign n2880 = i_wb_data[2:2] ;
assign n2881 = ~ ( n2880 ) ;
assign n2882 = sp[2:2] ;
assign n2883 =  ( n2881 ) ^ ( n2882 )  ;
assign n2884 =  ( n2883 ) ^ ( n2282 )  ;
assign n2885 =  ( n2879 ) ? ( n2884 ) : ( n2289 ) ;
assign n2886 =  ( n2876 ) ? ( bv_1_0_n2 ) : ( n2885 ) ;
assign n2887 =  ( n30 ) | ( n39 )  ;
assign n2888 =  ( n2887 ) ? ( bv_1_0_n2 ) : ( n2590 ) ;
assign n2889 =  ( n2875 ) ? ( n2886 ) : ( n2888 ) ;
assign n2890 = ~ ( n2889 ) ;
assign n2891 =  ( n2874 ) | ( n2890 )  ;
assign n2892 = ~ ( n2891 ) ;
assign n2893 =  ( n2873 ) ^ ( n2889 )  ;
assign n2894 = ~ ( n2893 ) ;
assign n2895 =  ( n354 ) | ( n363 )  ;
assign n2896 =  ( n373 ) | ( n382 )  ;
assign n2897 = ki[15:15] ;
assign n2898 =  ( n2897 ) == ( bv_1_0_n2 )  ;
assign n2899 =  ( n2898 ) | ( n391 )  ;
assign n2900 = i_wb_data[0:0] ;
assign n2901 = ~ ( n2900 ) ;
assign n2902 =  ( bv_1_1_n5 ) ^ ( n2901 )  ;
assign n2903 = sp[0:0] ;
assign n2904 =  ( n2902 ) ^ ( n2903 )  ;
assign n2905 = i_wb_data[0:0] ;
assign n2906 = ~ ( n2905 ) ;
assign n2907 =  ( bv_1_1_n5 ) ^ ( n2906 )  ;
assign n2908 = sp[0:0] ;
assign n2909 =  ( n2907 ) ^ ( n2908 )  ;
assign n2910 = ~ ( n2909 ) ;
assign n2911 =  ( n2899 ) ? ( n2904 ) : ( n2910 ) ;
assign n2912 =  ( n2896 ) ? ( bv_1_0_n2 ) : ( n2911 ) ;
assign n2913 =  ( n373 ) | ( n382 )  ;
assign n2914 =  ( n2913 ) ? ( bv_1_0_n2 ) : ( n2616 ) ;
assign n2915 =  ( n2895 ) ? ( n2912 ) : ( n2914 ) ;
assign n2916 = ~ ( n2915 ) ;
assign n2917 =  ( n2894 ) | ( n2916 )  ;
assign n2918 = ~ ( n2917 ) ;
assign n2919 =  ( n2892 ) | ( n2918 )  ;
assign n2920 = ~ ( n2919 ) ;
assign n2921 =  ( n2858 ) | ( n2920 )  ;
assign n2922 = ~ ( n2468 ) ;
assign n2923 =  ( n2922 ) ^ ( n2483 )  ;
assign n2924 =  ( n2923 ) ^ ( n2500 )  ;
assign n2925 =  ( n2924 ) ^ ( n2517 )  ;
assign n2926 =  ( n2925 ) ^ ( n2548 )  ;
assign n2927 = ~ ( n2926 ) ;
assign n2928 =  ( n2921 ) | ( n2927 )  ;
assign n2929 = ~ ( n2928 ) ;
assign n2930 =  ( n2846 ) ^ ( n2856 )  ;
assign n2931 = ~ ( n2930 ) ;
assign n2932 = ~ ( n2468 ) ;
assign n2933 =  ( n2919 ) ^ ( n2932 )  ;
assign n2934 =  ( n2933 ) ^ ( n2483 )  ;
assign n2935 =  ( n2934 ) ^ ( n2500 )  ;
assign n2936 =  ( n2935 ) ^ ( n2517 )  ;
assign n2937 =  ( n2936 ) ^ ( n2548 )  ;
assign n2938 = ~ ( n2937 ) ;
assign n2939 =  ( n2931 ) | ( n2938 )  ;
assign n2940 = ~ ( n2939 ) ;
assign n2941 =  ( n2929 ) | ( n2940 )  ;
assign n2942 =  ( n2846 ) ^ ( n2856 )  ;
assign n2943 =  ( n2942 ) ^ ( n2919 )  ;
assign n2944 = ~ ( n2468 ) ;
assign n2945 =  ( n2943 ) ^ ( n2944 )  ;
assign n2946 =  ( n2945 ) ^ ( n2483 )  ;
assign n2947 =  ( n2946 ) ^ ( n2500 )  ;
assign n2948 =  ( n2947 ) ^ ( n2517 )  ;
assign n2949 =  ( n2948 ) ^ ( n2548 )  ;
assign n2950 = ~ ( n2949 ) ;
assign n2951 =  ( n2578 ) ^ ( n2594 )  ;
assign n2952 =  ( n2951 ) ^ ( n2620 )  ;
assign n2953 = ~ ( n2952 ) ;
assign n2954 =  ( n2950 ) | ( n2953 )  ;
assign n2955 = ~ ( n2954 ) ;
assign n2956 =  ( n2941 ) | ( n2955 )  ;
assign n2957 = ~ ( n2956 ) ;
assign n2958 = ~ ( n2846 ) ;
assign n2959 = ~ ( n2856 ) ;
assign n2960 =  ( n2958 ) | ( n2959 )  ;
assign n2961 = ~ ( n2960 ) ;
assign n2962 = ~ ( n2919 ) ;
assign n2963 = ~ ( n2468 ) ;
assign n2964 =  ( n2963 ) ^ ( n2483 )  ;
assign n2965 =  ( n2964 ) ^ ( n2500 )  ;
assign n2966 =  ( n2965 ) ^ ( n2517 )  ;
assign n2967 =  ( n2966 ) ^ ( n2548 )  ;
assign n2968 = ~ ( n2967 ) ;
assign n2969 =  ( n2962 ) | ( n2968 )  ;
assign n2970 = ~ ( n2969 ) ;
assign n2971 =  ( n2961 ) | ( n2970 )  ;
assign n2972 = ~ ( n2971 ) ;
assign n2973 =  ( n2957 ) | ( n2972 )  ;
assign n2974 = ~ ( n2973 ) ;
assign n2975 = ~ ( n2928 ) ;
assign n2976 = ~ ( n2939 ) ;
assign n2977 =  ( n2975 ) | ( n2976 )  ;
assign n2978 = ~ ( n2954 ) ;
assign n2979 =  ( n2977 ) | ( n2978 )  ;
assign n2980 =  ( n2979 ) ^ ( n2971 )  ;
assign n2981 = ~ ( n2980 ) ;
assign n2982 =  ( bv_1_1_n5 ) ^ ( n2552 )  ;
assign n2983 =  ( n2982 ) ^ ( n2561 )  ;
assign n2984 =  ( n2983 ) ^ ( n2624 )  ;
assign n2985 =  ( n2984 ) ^ ( n2144 )  ;
assign n2986 =  ( n2985 ) ^ ( n2160 )  ;
assign n2987 =  ( n2986 ) ^ ( n2177 )  ;
assign n2988 =  ( n2987 ) ^ ( n2194 )  ;
assign n2989 =  ( n2988 ) ^ ( n2223 )  ;
assign n2990 =  ( n2989 ) ^ ( n2263 )  ;
assign n2991 =  ( n2990 ) ^ ( n2309 )  ;
assign n2992 = ~ ( n2991 ) ;
assign n2993 =  ( n2981 ) | ( n2992 )  ;
assign n2994 = ~ ( n2993 ) ;
assign n2995 =  ( n2974 ) | ( n2994 )  ;
assign n2996 = ~ ( n2995 ) ;
assign n2997 =  ( n2633 ) | ( n2643 )  ;
assign n2998 =  ( n2997 ) | ( n2657 )  ;
assign n2999 =  ( n2998 ) ^ ( n2672 )  ;
assign n3000 =  ( n2999 ) ^ ( n2227 )  ;
assign n3001 =  ( n3000 ) ^ ( n2237 )  ;
assign n3002 =  ( n3001 ) ^ ( n2314 )  ;
assign n3003 =  ( n1838 ) | ( n1847 )  ;
assign n3004 =  ( n3003 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n3005 = ~ ( n3004 ) ;
assign n3006 =  ( n3002 ) ^ ( n3005 )  ;
assign n3007 =  ( n3006 ) ^ ( n1879 )  ;
assign n3008 =  ( n3007 ) ^ ( n1896 )  ;
assign n3009 =  ( n3008 ) ^ ( n1913 )  ;
assign n3010 =  ( n3009 ) ^ ( n1948 )  ;
assign n3011 =  ( n3010 ) ^ ( n2357 )  ;
assign n3012 = ~ ( n3011 ) ;
assign n3013 =  ( n2996 ) | ( n3012 )  ;
assign n3014 = ~ ( n3013 ) ;
assign n3015 = ~ ( n2973 ) ;
assign n3016 =  ( n3015 ) | ( n2994 )  ;
assign n3017 =  ( n2633 ) | ( n2643 )  ;
assign n3018 =  ( n3017 ) | ( n2657 )  ;
assign n3019 =  ( n3016 ) ^ ( n3018 )  ;
assign n3020 =  ( n3019 ) ^ ( n2672 )  ;
assign n3021 =  ( n3020 ) ^ ( n2227 )  ;
assign n3022 =  ( n3021 ) ^ ( n2237 )  ;
assign n3023 =  ( n3022 ) ^ ( n2314 )  ;
assign n3024 =  ( n1838 ) | ( n1847 )  ;
assign n3025 =  ( n3024 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n3026 = ~ ( n3025 ) ;
assign n3027 =  ( n3023 ) ^ ( n3026 )  ;
assign n3028 =  ( n3027 ) ^ ( n1879 )  ;
assign n3029 =  ( n3028 ) ^ ( n1896 )  ;
assign n3030 =  ( n3029 ) ^ ( n1913 )  ;
assign n3031 =  ( n3030 ) ^ ( n1948 )  ;
assign n3032 =  ( n3031 ) ^ ( n2357 )  ;
assign n3033 = ~ ( n3032 ) ;
assign n3034 =  ( n354 ) | ( n363 )  ;
assign n3035 =  ( n373 ) | ( n382 )  ;
assign n3036 =  ( n3035 ) ? ( bv_1_0_n2 ) : ( n2307 ) ;
assign n3037 =  ( n373 ) | ( n382 )  ;
assign n3038 =  ( n3037 ) ? ( bv_1_0_n2 ) : ( n1997 ) ;
assign n3039 =  ( n3034 ) ? ( n3036 ) : ( n3038 ) ;
assign n3040 = ~ ( n3039 ) ;
assign n3041 =  ( n3033 ) | ( n3040 )  ;
assign n3042 = ~ ( n3041 ) ;
assign n3043 =  ( n3014 ) | ( n3042 )  ;
assign n3044 = ~ ( n3043 ) ;
assign n3045 =  ( n2743 ) | ( n3044 )  ;
assign n3046 = ~ ( n2692 ) ;
assign n3047 =  ( n2675 ) | ( n3046 )  ;
assign n3048 =  ( bv_1_1_n5 ) ^ ( n3047 )  ;
assign n3049 =  ( n3048 ) ^ ( n2361 )  ;
assign n3050 =  ( n3049 ) ^ ( n2371 )  ;
assign n3051 =  ( n3050 ) ^ ( n1952 )  ;
assign n3052 =  ( n3051 ) ^ ( n1963 )  ;
assign n3053 =  ( n3052 ) ^ ( n1513 )  ;
assign n3054 =  ( n3053 ) ^ ( n1538 )  ;
assign n3055 =  ( n3054 ) ^ ( n1564 )  ;
assign n3056 =  ( n3055 ) ^ ( n1590 )  ;
assign n3057 =  ( n3056 ) ^ ( n1628 )  ;
assign n3058 =  ( n3057 ) ^ ( n2016 )  ;
assign n3059 = ~ ( n3058 ) ;
assign n3060 =  ( n3045 ) | ( n3059 )  ;
assign n3061 = ~ ( n3060 ) ;
assign n3062 =  ( n2723 ) | ( n3061 )  ;
assign n3063 = ~ ( n3062 ) ;
assign n3064 =  ( n2454 ) | ( n3063 )  ;
assign n3065 = ~ ( n3064 ) ;
assign n3066 =  ( n2441 ) | ( n3065 )  ;
assign n3067 = ~ ( n2110 ) ;
assign n3068 =  ( n3067 ) | ( n2453 )  ;
assign n3069 = ~ ( n2742 ) ;
assign n3070 =  ( n3068 ) | ( n3069 )  ;
assign n3071 =  ( bv_1_1_n5 ) ^ ( n3043 )  ;
assign n3072 = ~ ( n2692 ) ;
assign n3073 =  ( n2675 ) | ( n3072 )  ;
assign n3074 =  ( n3071 ) ^ ( n3073 )  ;
assign n3075 =  ( n3074 ) ^ ( n2361 )  ;
assign n3076 =  ( n3075 ) ^ ( n2371 )  ;
assign n3077 =  ( n3076 ) ^ ( n1952 )  ;
assign n3078 =  ( n3077 ) ^ ( n1963 )  ;
assign n3079 =  ( n3078 ) ^ ( n1513 )  ;
assign n3080 =  ( n3079 ) ^ ( n1538 )  ;
assign n3081 =  ( n3080 ) ^ ( n1564 )  ;
assign n3082 =  ( n3081 ) ^ ( n1590 )  ;
assign n3083 =  ( n3082 ) ^ ( n1628 )  ;
assign n3084 =  ( n3083 ) ^ ( n2016 )  ;
assign n3085 = ~ ( n3084 ) ;
assign n3086 =  ( n3070 ) | ( n3085 )  ;
assign n3087 = ki[0:0] ;
assign n3088 =  ( n3087 ) == ( bv_1_1_n5 )  ;
assign n3089 = ki[1:1] ;
assign n3090 =  ( n3089 ) == ( bv_1_0_n2 )  ;
assign n3091 =  ( n3088 ) | ( n3090 )  ;
assign n3092 = ki[1:1] ;
assign n3093 =  ( n3092 ) == ( bv_1_1_n5 )  ;
assign n3094 = ki[0:0] ;
assign n3095 =  ( n3094 ) == ( bv_1_1_n5 )  ;
assign n3096 =  ( n3093 ) | ( n3095 )  ;
assign n3097 = ki[1:1] ;
assign n3098 =  ( n3097 ) == ( bv_1_1_n5 )  ;
assign n3099 = i_wb_data[13:13] ;
assign n3100 = ~ ( n3099 ) ;
assign n3101 = sp[13:13] ;
assign n3102 =  ( n3100 ) ^ ( n3101 )  ;
assign n3103 =  ( n3102 ) ^ ( n245 )  ;
assign n3104 =  ( n3098 ) ? ( n451 ) : ( n3103 ) ;
assign n3105 =  ( n3096 ) ? ( n3104 ) : ( bv_1_0_n2 ) ;
assign n3106 =  ( n3091 ) ? ( n2762 ) : ( n3105 ) ;
assign n3107 = ~ ( n3106 ) ;
assign n3108 =  ( n2120 ) | ( n2129 )  ;
assign n3109 =  ( n1838 ) | ( n1847 )  ;
assign n3110 = ki[3:3] ;
assign n3111 =  ( n3110 ) == ( bv_1_0_n2 )  ;
assign n3112 =  ( n3111 ) | ( n1856 )  ;
assign n3113 = i_wb_data[11:11] ;
assign n3114 = ~ ( n3113 ) ;
assign n3115 = sp[11:11] ;
assign n3116 =  ( n3114 ) ^ ( n3115 )  ;
assign n3117 =  ( n3116 ) ^ ( n423 )  ;
assign n3118 =  ( n3112 ) ? ( n3117 ) : ( n648 ) ;
assign n3119 =  ( n3109 ) ? ( bv_1_0_n2 ) : ( n3118 ) ;
assign n3120 =  ( n1838 ) | ( n1847 )  ;
assign n3121 =  ( n3120 ) ? ( bv_1_0_n2 ) : ( n2775 ) ;
assign n3122 =  ( n3108 ) ? ( n3119 ) : ( n3121 ) ;
assign n3123 = ~ ( n3122 ) ;
assign n3124 =  ( n3107 ) | ( n3123 )  ;
assign n3125 =  ( n1456 ) | ( n1465 )  ;
assign n3126 =  ( n1475 ) | ( n1484 )  ;
assign n3127 = ki[5:5] ;
assign n3128 =  ( n3127 ) == ( bv_1_0_n2 )  ;
assign n3129 =  ( n3128 ) | ( n1493 )  ;
assign n3130 = i_wb_data[9:9] ;
assign n3131 = ~ ( n3130 ) ;
assign n3132 = sp[9:9] ;
assign n3133 =  ( n3131 ) ^ ( n3132 )  ;
assign n3134 =  ( n3133 ) ^ ( n734 )  ;
assign n3135 =  ( n3129 ) ? ( n3134 ) : ( n985 ) ;
assign n3136 =  ( n3126 ) ? ( bv_1_0_n2 ) : ( n3135 ) ;
assign n3137 =  ( n1475 ) | ( n1484 )  ;
assign n3138 =  ( n3137 ) ? ( bv_1_0_n2 ) : ( n2792 ) ;
assign n3139 =  ( n3125 ) ? ( n3136 ) : ( n3138 ) ;
assign n3140 = ~ ( n3139 ) ;
assign n3141 =  ( n3124 ) | ( n3140 )  ;
assign n3142 =  ( n1257 ) | ( n1266 )  ;
assign n3143 =  ( n873 ) | ( n882 )  ;
assign n3144 = ki[7:7] ;
assign n3145 =  ( n3144 ) == ( bv_1_0_n2 )  ;
assign n3146 =  ( n3145 ) | ( n891 )  ;
assign n3147 = i_wb_data[7:7] ;
assign n3148 = ~ ( n3147 ) ;
assign n3149 = sp[7:7] ;
assign n3150 =  ( n3148 ) ^ ( n3149 )  ;
assign n3151 =  ( n3150 ) ^ ( n330 )  ;
assign n3152 =  ( n3146 ) ? ( n3151 ) : ( n1035 ) ;
assign n3153 =  ( n3143 ) ? ( bv_1_0_n2 ) : ( n3152 ) ;
assign n3154 =  ( n873 ) | ( n882 )  ;
assign n3155 =  ( n3154 ) ? ( bv_1_0_n2 ) : ( n2809 ) ;
assign n3156 =  ( n3142 ) ? ( n3153 ) : ( n3155 ) ;
assign n3157 = ~ ( n3156 ) ;
assign n3158 =  ( n3141 ) | ( n3157 )  ;
assign n3159 = ~ ( n3158 ) ;
assign n3160 =  ( n3106 ) ^ ( n3122 )  ;
assign n3161 = ~ ( n3160 ) ;
assign n3162 =  ( n3139 ) ^ ( n3156 )  ;
assign n3163 = ~ ( n3162 ) ;
assign n3164 =  ( n3161 ) | ( n3163 )  ;
assign n3165 = ~ ( n3164 ) ;
assign n3166 =  ( n3159 ) | ( n3165 )  ;
assign n3167 =  ( n3106 ) ^ ( n3122 )  ;
assign n3168 =  ( n3167 ) ^ ( n3139 )  ;
assign n3169 =  ( n3168 ) ^ ( n3156 )  ;
assign n3170 = ~ ( n3169 ) ;
assign n3171 =  ( n908 ) | ( n917 )  ;
assign n3172 =  ( n532 ) | ( n541 )  ;
assign n3173 = ki[9:9] ;
assign n3174 =  ( n3173 ) == ( bv_1_0_n2 )  ;
assign n3175 =  ( n3174 ) | ( n550 )  ;
assign n3176 = i_wb_data[5:5] ;
assign n3177 = ~ ( n3176 ) ;
assign n3178 = sp[5:5] ;
assign n3179 =  ( n3177 ) ^ ( n3178 )  ;
assign n3180 =  ( n3179 ) ^ ( n241 )  ;
assign n3181 =  ( n3175 ) ? ( n3180 ) : ( n2013 ) ;
assign n3182 =  ( n3172 ) ? ( bv_1_0_n2 ) : ( n3181 ) ;
assign n3183 =  ( n532 ) | ( n541 )  ;
assign n3184 =  ( n3183 ) ? ( bv_1_0_n2 ) : ( n2838 ) ;
assign n3185 =  ( n3171 ) ? ( n3182 ) : ( n3184 ) ;
assign n3186 = ~ ( n3185 ) ;
assign n3187 =  ( n3170 ) | ( n3186 )  ;
assign n3188 = ~ ( n3187 ) ;
assign n3189 =  ( n3166 ) | ( n3188 )  ;
assign n3190 = ~ ( n3189 ) ;
assign n3191 = ~ ( n3106 ) ;
assign n3192 = ~ ( n3122 ) ;
assign n3193 =  ( n3191 ) | ( n3192 )  ;
assign n3194 = ~ ( n3193 ) ;
assign n3195 = ~ ( n3139 ) ;
assign n3196 = ~ ( n3156 ) ;
assign n3197 =  ( n3195 ) | ( n3196 )  ;
assign n3198 = ~ ( n3197 ) ;
assign n3199 =  ( n3194 ) | ( n3198 )  ;
assign n3200 = ~ ( n3199 ) ;
assign n3201 =  ( n3190 ) | ( n3200 )  ;
assign n3202 =  ( n567 ) | ( n576 )  ;
assign n3203 =  ( n586 ) | ( n595 )  ;
assign n3204 = ki[11:11] ;
assign n3205 =  ( n3204 ) == ( bv_1_0_n2 )  ;
assign n3206 =  ( n3205 ) | ( n604 )  ;
assign n3207 = i_wb_data[3:3] ;
assign n3208 = ~ ( n3207 ) ;
assign n3209 = sp[3:3] ;
assign n3210 =  ( n3208 ) ^ ( n3209 )  ;
assign n3211 =  ( n3210 ) ^ ( n326 )  ;
assign n3212 =  ( n3206 ) ? ( n3211 ) : ( n2306 ) ;
assign n3213 =  ( n3203 ) ? ( bv_1_0_n2 ) : ( n3212 ) ;
assign n3214 =  ( n586 ) | ( n595 )  ;
assign n3215 =  ( n3214 ) ? ( bv_1_0_n2 ) : ( n2869 ) ;
assign n3216 =  ( n3202 ) ? ( n3213 ) : ( n3215 ) ;
assign n3217 = ~ ( n3216 ) ;
assign n3218 =  ( n11 ) | ( n20 )  ;
assign n3219 =  ( n30 ) | ( n39 )  ;
assign n3220 = ki[13:13] ;
assign n3221 =  ( n3220 ) == ( bv_1_0_n2 )  ;
assign n3222 =  ( n3221 ) | ( n48 )  ;
assign n3223 = i_wb_data[1:1] ;
assign n3224 = ~ ( n3223 ) ;
assign n3225 = sp[1:1] ;
assign n3226 =  ( n3224 ) ^ ( n3225 )  ;
assign n3227 =  ( n3226 ) ^ ( n237 )  ;
assign n3228 =  ( n3222 ) ? ( n3227 ) : ( n2615 ) ;
assign n3229 =  ( n3219 ) ? ( bv_1_0_n2 ) : ( n3228 ) ;
assign n3230 =  ( n30 ) | ( n39 )  ;
assign n3231 =  ( n3230 ) ? ( bv_1_0_n2 ) : ( n2885 ) ;
assign n3232 =  ( n3218 ) ? ( n3229 ) : ( n3231 ) ;
assign n3233 = ~ ( n3232 ) ;
assign n3234 =  ( n3217 ) | ( n3233 )  ;
assign n3235 = ~ ( n3234 ) ;
assign n3236 =  ( n3216 ) ^ ( n3232 )  ;
assign n3237 = ~ ( n3236 ) ;
assign n3238 =  ( n354 ) | ( n363 )  ;
assign n3239 = ki[15:15] ;
assign n3240 = ~ ( n3239 ) ;
assign n3241 = ki[14:14] ;
assign n3242 = ~ ( n3241 ) ;
assign n3243 = ki[13:13] ;
assign n3244 = ~ ( n3243 ) ;
assign n3245 =  ( n3242 ) | ( n3244 )  ;
assign n3246 = ~ ( n3245 ) ;
assign n3247 =  ( n3240 ) | ( n3246 )  ;
assign n3248 = ~ ( n3247 ) ;
assign n3249 =  ( n373 ) | ( n382 )  ;
assign n3250 =  ( n3249 ) ? ( bv_1_0_n2 ) : ( n2911 ) ;
assign n3251 =  ( n3238 ) ? ( n3248 ) : ( n3250 ) ;
assign n3252 = ~ ( n3251 ) ;
assign n3253 =  ( n3237 ) | ( n3252 )  ;
assign n3254 = ~ ( n3253 ) ;
assign n3255 =  ( n3235 ) | ( n3254 )  ;
assign n3256 = ~ ( n3255 ) ;
assign n3257 =  ( n3201 ) | ( n3256 )  ;
assign n3258 =  ( n2763 ) ^ ( n2779 )  ;
assign n3259 =  ( n3258 ) ^ ( n2796 )  ;
assign n3260 =  ( n3259 ) ^ ( n2813 )  ;
assign n3261 =  ( n3260 ) ^ ( n2842 )  ;
assign n3262 = ~ ( n3261 ) ;
assign n3263 =  ( n3257 ) | ( n3262 )  ;
assign n3264 = ~ ( n3263 ) ;
assign n3265 =  ( n3189 ) ^ ( n3199 )  ;
assign n3266 = ~ ( n3265 ) ;
assign n3267 =  ( n3255 ) ^ ( n2763 )  ;
assign n3268 =  ( n3267 ) ^ ( n2779 )  ;
assign n3269 =  ( n3268 ) ^ ( n2796 )  ;
assign n3270 =  ( n3269 ) ^ ( n2813 )  ;
assign n3271 =  ( n3270 ) ^ ( n2842 )  ;
assign n3272 = ~ ( n3271 ) ;
assign n3273 =  ( n3266 ) | ( n3272 )  ;
assign n3274 = ~ ( n3273 ) ;
assign n3275 =  ( n3264 ) | ( n3274 )  ;
assign n3276 =  ( n3189 ) ^ ( n3199 )  ;
assign n3277 =  ( n3276 ) ^ ( n3255 )  ;
assign n3278 =  ( n3277 ) ^ ( n2763 )  ;
assign n3279 =  ( n3278 ) ^ ( n2779 )  ;
assign n3280 =  ( n3279 ) ^ ( n2796 )  ;
assign n3281 =  ( n3280 ) ^ ( n2813 )  ;
assign n3282 =  ( n3281 ) ^ ( n2842 )  ;
assign n3283 = ~ ( n3282 ) ;
assign n3284 =  ( n2873 ) ^ ( n2889 )  ;
assign n3285 =  ( n3284 ) ^ ( n2915 )  ;
assign n3286 = ~ ( n3285 ) ;
assign n3287 =  ( n3283 ) | ( n3286 )  ;
assign n3288 = ~ ( n3287 ) ;
assign n3289 =  ( n3275 ) | ( n3288 )  ;
assign n3290 = ~ ( n3289 ) ;
assign n3291 = ~ ( n3189 ) ;
assign n3292 = ~ ( n3199 ) ;
assign n3293 =  ( n3291 ) | ( n3292 )  ;
assign n3294 = ~ ( n3293 ) ;
assign n3295 = ~ ( n3255 ) ;
assign n3296 =  ( n2763 ) ^ ( n2779 )  ;
assign n3297 =  ( n3296 ) ^ ( n2796 )  ;
assign n3298 =  ( n3297 ) ^ ( n2813 )  ;
assign n3299 =  ( n3298 ) ^ ( n2842 )  ;
assign n3300 = ~ ( n3299 ) ;
assign n3301 =  ( n3295 ) | ( n3300 )  ;
assign n3302 = ~ ( n3301 ) ;
assign n3303 =  ( n3294 ) | ( n3302 )  ;
assign n3304 = ~ ( n3303 ) ;
assign n3305 =  ( n3290 ) | ( n3304 )  ;
assign n3306 = ~ ( n3305 ) ;
assign n3307 =  ( n3264 ) | ( n3274 )  ;
assign n3308 =  ( n3307 ) | ( n3288 )  ;
assign n3309 =  ( n3308 ) ^ ( n3303 )  ;
assign n3310 = ~ ( n3309 ) ;
assign n3311 =  ( n2846 ) ^ ( n2856 )  ;
assign n3312 =  ( n3311 ) ^ ( n2919 )  ;
assign n3313 = ~ ( n2468 ) ;
assign n3314 =  ( n3312 ) ^ ( n3313 )  ;
assign n3315 =  ( n3314 ) ^ ( n2483 )  ;
assign n3316 =  ( n3315 ) ^ ( n2500 )  ;
assign n3317 =  ( n3316 ) ^ ( n2517 )  ;
assign n3318 =  ( n3317 ) ^ ( n2548 )  ;
assign n3319 =  ( n3318 ) ^ ( n2578 )  ;
assign n3320 =  ( n3319 ) ^ ( n2594 )  ;
assign n3321 =  ( n3320 ) ^ ( n2620 )  ;
assign n3322 = ~ ( n3321 ) ;
assign n3323 =  ( n3310 ) | ( n3322 )  ;
assign n3324 = ~ ( n3323 ) ;
assign n3325 =  ( n3306 ) | ( n3324 )  ;
assign n3326 = ~ ( n3325 ) ;
assign n3327 = ~ ( n2928 ) ;
assign n3328 = ~ ( n2939 ) ;
assign n3329 =  ( n3327 ) | ( n3328 )  ;
assign n3330 = ~ ( n2954 ) ;
assign n3331 =  ( n3329 ) | ( n3330 )  ;
assign n3332 =  ( bv_1_1_n5 ) ^ ( n3331 )  ;
assign n3333 =  ( n3332 ) ^ ( n2971 )  ;
assign n3334 =  ( n3333 ) ^ ( n2552 )  ;
assign n3335 =  ( n3334 ) ^ ( n2561 )  ;
assign n3336 =  ( n3335 ) ^ ( n2624 )  ;
assign n3337 =  ( n3336 ) ^ ( n2144 )  ;
assign n3338 =  ( n3337 ) ^ ( n2160 )  ;
assign n3339 =  ( n3338 ) ^ ( n2177 )  ;
assign n3340 =  ( n3339 ) ^ ( n2194 )  ;
assign n3341 =  ( n3340 ) ^ ( n2223 )  ;
assign n3342 =  ( n3341 ) ^ ( n2263 )  ;
assign n3343 =  ( n3342 ) ^ ( n2309 )  ;
assign n3344 = ~ ( n3343 ) ;
assign n3345 =  ( n3326 ) | ( n3344 )  ;
assign n3346 = ~ ( n2973 ) ;
assign n3347 =  ( n3346 ) | ( n2994 )  ;
assign n3348 =  ( n2633 ) | ( n2643 )  ;
assign n3349 =  ( n3348 ) | ( n2657 )  ;
assign n3350 =  ( n3347 ) ^ ( n3349 )  ;
assign n3351 =  ( n3350 ) ^ ( n2672 )  ;
assign n3352 =  ( n3351 ) ^ ( n2227 )  ;
assign n3353 =  ( n3352 ) ^ ( n2237 )  ;
assign n3354 =  ( n3353 ) ^ ( n2314 )  ;
assign n3355 =  ( n1838 ) | ( n1847 )  ;
assign n3356 =  ( n3355 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n3357 = ~ ( n3356 ) ;
assign n3358 =  ( n3354 ) ^ ( n3357 )  ;
assign n3359 =  ( n3358 ) ^ ( n1879 )  ;
assign n3360 =  ( n3359 ) ^ ( n1896 )  ;
assign n3361 =  ( n3360 ) ^ ( n1913 )  ;
assign n3362 =  ( n3361 ) ^ ( n1948 )  ;
assign n3363 =  ( n3362 ) ^ ( n2357 )  ;
assign n3364 =  ( n3363 ) ^ ( n3039 )  ;
assign n3365 = ~ ( n3364 ) ;
assign n3366 =  ( n3345 ) | ( n3365 )  ;
assign n3367 = ~ ( n3366 ) ;
assign n3368 = ~ ( n3323 ) ;
assign n3369 =  ( n3306 ) | ( n3368 )  ;
assign n3370 = ~ ( n3369 ) ;
assign n3371 =  ( n3370 ) | ( n3344 )  ;
assign n3372 = ~ ( n3371 ) ;
assign n3373 = ~ ( n2973 ) ;
assign n3374 =  ( n3373 ) | ( n2994 )  ;
assign n3375 =  ( n3372 ) ^ ( n3374 )  ;
assign n3376 =  ( n2633 ) | ( n2643 )  ;
assign n3377 =  ( n3376 ) | ( n2657 )  ;
assign n3378 =  ( n3375 ) ^ ( n3377 )  ;
assign n3379 =  ( n3378 ) ^ ( n2672 )  ;
assign n3380 =  ( n3379 ) ^ ( n2227 )  ;
assign n3381 =  ( n3380 ) ^ ( n2237 )  ;
assign n3382 =  ( n3381 ) ^ ( n2314 )  ;
assign n3383 =  ( n1838 ) | ( n1847 )  ;
assign n3384 =  ( n3383 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n3385 = ~ ( n3384 ) ;
assign n3386 =  ( n3382 ) ^ ( n3385 )  ;
assign n3387 =  ( n3386 ) ^ ( n1879 )  ;
assign n3388 =  ( n3387 ) ^ ( n1896 )  ;
assign n3389 =  ( n3388 ) ^ ( n1913 )  ;
assign n3390 =  ( n3389 ) ^ ( n1948 )  ;
assign n3391 =  ( n3390 ) ^ ( n2357 )  ;
assign n3392 =  ( n3391 ) ^ ( n3039 )  ;
assign n3393 = ~ ( n3392 ) ;
assign n3394 = ki[0:0] ;
assign n3395 =  ( n3394 ) == ( bv_1_1_n5 )  ;
assign n3396 = ki[1:1] ;
assign n3397 =  ( n3396 ) == ( bv_1_0_n2 )  ;
assign n3398 =  ( n3395 ) | ( n3397 )  ;
assign n3399 = ki[1:1] ;
assign n3400 =  ( n3399 ) == ( bv_1_1_n5 )  ;
assign n3401 = ki[0:0] ;
assign n3402 =  ( n3401 ) == ( bv_1_1_n5 )  ;
assign n3403 =  ( n3400 ) | ( n3402 )  ;
assign n3404 = ki[1:1] ;
assign n3405 =  ( n3404 ) == ( bv_1_1_n5 )  ;
assign n3406 = i_wb_data[12:12] ;
assign n3407 = ~ ( n3406 ) ;
assign n3408 = sp[12:12] ;
assign n3409 =  ( n3407 ) ^ ( n3408 )  ;
assign n3410 =  ( n3409 ) ^ ( n427 )  ;
assign n3411 =  ( n3405 ) ? ( n434 ) : ( n3410 ) ;
assign n3412 =  ( n3403 ) ? ( n3411 ) : ( bv_1_0_n2 ) ;
assign n3413 =  ( n3398 ) ? ( n3105 ) : ( n3412 ) ;
assign n3414 = ~ ( n3413 ) ;
assign n3415 =  ( n2120 ) | ( n2129 )  ;
assign n3416 =  ( n1838 ) | ( n1847 )  ;
assign n3417 = ki[3:3] ;
assign n3418 =  ( n3417 ) == ( bv_1_0_n2 )  ;
assign n3419 =  ( n3418 ) | ( n1856 )  ;
assign n3420 = i_wb_data[10:10] ;
assign n3421 = ~ ( n3420 ) ;
assign n3422 = sp[10:10] ;
assign n3423 =  ( n3421 ) ^ ( n3422 )  ;
assign n3424 =  ( n3423 ) ^ ( n738 )  ;
assign n3425 =  ( n3419 ) ? ( n3424 ) : ( n745 ) ;
assign n3426 =  ( n3416 ) ? ( bv_1_0_n2 ) : ( n3425 ) ;
assign n3427 =  ( n1838 ) | ( n1847 )  ;
assign n3428 =  ( n3427 ) ? ( bv_1_0_n2 ) : ( n3118 ) ;
assign n3429 =  ( n3415 ) ? ( n3426 ) : ( n3428 ) ;
assign n3430 = ~ ( n3429 ) ;
assign n3431 =  ( n3414 ) | ( n3430 )  ;
assign n3432 =  ( n1456 ) | ( n1465 )  ;
assign n3433 =  ( n1475 ) | ( n1484 )  ;
assign n3434 = ki[5:5] ;
assign n3435 =  ( n3434 ) == ( bv_1_0_n2 )  ;
assign n3436 =  ( n3435 ) | ( n1493 )  ;
assign n3437 = i_wb_data[8:8] ;
assign n3438 = ~ ( n3437 ) ;
assign n3439 = sp[8:8] ;
assign n3440 =  ( n3438 ) ^ ( n3439 )  ;
assign n3441 =  ( n3440 ) ^ ( n1054 )  ;
assign n3442 =  ( n3436 ) ? ( n3441 ) : ( n1061 ) ;
assign n3443 =  ( n3433 ) ? ( bv_1_0_n2 ) : ( n3442 ) ;
assign n3444 =  ( n1475 ) | ( n1484 )  ;
assign n3445 =  ( n3444 ) ? ( bv_1_0_n2 ) : ( n3135 ) ;
assign n3446 =  ( n3432 ) ? ( n3443 ) : ( n3445 ) ;
assign n3447 = ~ ( n3446 ) ;
assign n3448 =  ( n3431 ) | ( n3447 )  ;
assign n3449 =  ( n1257 ) | ( n1266 )  ;
assign n3450 =  ( n873 ) | ( n882 )  ;
assign n3451 = ki[7:7] ;
assign n3452 =  ( n3451 ) == ( bv_1_0_n2 )  ;
assign n3453 =  ( n3452 ) | ( n891 )  ;
assign n3454 = i_wb_data[6:6] ;
assign n3455 = ~ ( n3454 ) ;
assign n3456 = sp[6:6] ;
assign n3457 =  ( n3455 ) ^ ( n3456 )  ;
assign n3458 =  ( n3457 ) ^ ( n1363 )  ;
assign n3459 =  ( n3453 ) ? ( n3458 ) : ( n1370 ) ;
assign n3460 =  ( n3450 ) ? ( bv_1_0_n2 ) : ( n3459 ) ;
assign n3461 =  ( n873 ) | ( n882 )  ;
assign n3462 =  ( n3461 ) ? ( bv_1_0_n2 ) : ( n3152 ) ;
assign n3463 =  ( n3449 ) ? ( n3460 ) : ( n3462 ) ;
assign n3464 = ~ ( n3463 ) ;
assign n3465 =  ( n3448 ) | ( n3464 )  ;
assign n3466 = ~ ( n3465 ) ;
assign n3467 =  ( n3413 ) ^ ( n3429 )  ;
assign n3468 = ~ ( n3467 ) ;
assign n3469 =  ( n3446 ) ^ ( n3463 )  ;
assign n3470 = ~ ( n3469 ) ;
assign n3471 =  ( n3468 ) | ( n3470 )  ;
assign n3472 = ~ ( n3471 ) ;
assign n3473 =  ( n3466 ) | ( n3472 )  ;
assign n3474 =  ( n3413 ) ^ ( n3429 )  ;
assign n3475 =  ( n3474 ) ^ ( n3446 )  ;
assign n3476 =  ( n3475 ) ^ ( n3463 )  ;
assign n3477 = ~ ( n3476 ) ;
assign n3478 =  ( n908 ) | ( n917 )  ;
assign n3479 =  ( n532 ) | ( n541 )  ;
assign n3480 = ki[9:9] ;
assign n3481 =  ( n3480 ) == ( bv_1_0_n2 )  ;
assign n3482 =  ( n3481 ) | ( n550 )  ;
assign n3483 = i_wb_data[4:4] ;
assign n3484 = ~ ( n3483 ) ;
assign n3485 = sp[4:4] ;
assign n3486 =  ( n3484 ) ^ ( n3485 )  ;
assign n3487 =  ( n3486 ) ^ ( n1989 )  ;
assign n3488 =  ( n3482 ) ? ( n3487 ) : ( n1996 ) ;
assign n3489 =  ( n3479 ) ? ( bv_1_0_n2 ) : ( n3488 ) ;
assign n3490 =  ( n532 ) | ( n541 )  ;
assign n3491 =  ( n3490 ) ? ( bv_1_0_n2 ) : ( n3181 ) ;
assign n3492 =  ( n3478 ) ? ( n3489 ) : ( n3491 ) ;
assign n3493 = ~ ( n3492 ) ;
assign n3494 =  ( n3477 ) | ( n3493 )  ;
assign n3495 = ~ ( n3494 ) ;
assign n3496 =  ( n3473 ) | ( n3495 )  ;
assign n3497 = ~ ( n3496 ) ;
assign n3498 = ~ ( n3413 ) ;
assign n3499 = ~ ( n3429 ) ;
assign n3500 =  ( n3498 ) | ( n3499 )  ;
assign n3501 = ~ ( n3500 ) ;
assign n3502 = ~ ( n3446 ) ;
assign n3503 = ~ ( n3463 ) ;
assign n3504 =  ( n3502 ) | ( n3503 )  ;
assign n3505 = ~ ( n3504 ) ;
assign n3506 =  ( n3501 ) | ( n3505 )  ;
assign n3507 = ~ ( n3506 ) ;
assign n3508 =  ( n3497 ) | ( n3507 )  ;
assign n3509 =  ( n3106 ) ^ ( n3122 )  ;
assign n3510 =  ( n3509 ) ^ ( n3139 )  ;
assign n3511 =  ( n3510 ) ^ ( n3156 )  ;
assign n3512 =  ( n3511 ) ^ ( n3185 )  ;
assign n3513 = ~ ( n3512 ) ;
assign n3514 =  ( n3508 ) | ( n3513 )  ;
assign n3515 =  ( n3216 ) ^ ( n3232 )  ;
assign n3516 =  ( n3515 ) ^ ( n3251 )  ;
assign n3517 = ~ ( n3516 ) ;
assign n3518 =  ( n3514 ) | ( n3517 )  ;
assign n3519 = ~ ( n3518 ) ;
assign n3520 =  ( n3496 ) ^ ( n3506 )  ;
assign n3521 = ~ ( n3520 ) ;
assign n3522 =  ( n3106 ) ^ ( n3122 )  ;
assign n3523 =  ( n3522 ) ^ ( n3139 )  ;
assign n3524 =  ( n3523 ) ^ ( n3156 )  ;
assign n3525 =  ( n3524 ) ^ ( n3185 )  ;
assign n3526 =  ( n3525 ) ^ ( n3216 )  ;
assign n3527 =  ( n3526 ) ^ ( n3232 )  ;
assign n3528 =  ( n3527 ) ^ ( n3251 )  ;
assign n3529 = ~ ( n3528 ) ;
assign n3530 =  ( n3521 ) | ( n3529 )  ;
assign n3531 = ~ ( n3530 ) ;
assign n3532 =  ( n3519 ) | ( n3531 )  ;
assign n3533 =  ( n3496 ) ^ ( n3506 )  ;
assign n3534 =  ( n3533 ) ^ ( n3106 )  ;
assign n3535 =  ( n3534 ) ^ ( n3122 )  ;
assign n3536 =  ( n3535 ) ^ ( n3139 )  ;
assign n3537 =  ( n3536 ) ^ ( n3156 )  ;
assign n3538 =  ( n3537 ) ^ ( n3185 )  ;
assign n3539 =  ( n3538 ) ^ ( n3216 )  ;
assign n3540 =  ( n3539 ) ^ ( n3232 )  ;
assign n3541 =  ( n3540 ) ^ ( n3251 )  ;
assign n3542 = ~ ( n3541 ) ;
assign n3543 = ki[15:15] ;
assign n3544 = ~ ( n3543 ) ;
assign n3545 =  ( n3542 ) | ( n3544 )  ;
assign n3546 =  ( n3545 ) | ( n3246 )  ;
assign n3547 = ~ ( n3546 ) ;
assign n3548 =  ( n3532 ) | ( n3547 )  ;
assign n3549 = ~ ( n3548 ) ;
assign n3550 = ~ ( n3496 ) ;
assign n3551 = ~ ( n3506 ) ;
assign n3552 =  ( n3550 ) | ( n3551 )  ;
assign n3553 = ~ ( n3552 ) ;
assign n3554 =  ( n3106 ) ^ ( n3122 )  ;
assign n3555 =  ( n3554 ) ^ ( n3139 )  ;
assign n3556 =  ( n3555 ) ^ ( n3156 )  ;
assign n3557 =  ( n3556 ) ^ ( n3185 )  ;
assign n3558 = ~ ( n3557 ) ;
assign n3559 =  ( n3216 ) ^ ( n3232 )  ;
assign n3560 =  ( n3559 ) ^ ( n3251 )  ;
assign n3561 = ~ ( n3560 ) ;
assign n3562 =  ( n3558 ) | ( n3561 )  ;
assign n3563 = ~ ( n3562 ) ;
assign n3564 =  ( n3553 ) | ( n3563 )  ;
assign n3565 = ~ ( n3564 ) ;
assign n3566 =  ( n3549 ) | ( n3565 )  ;
assign n3567 = ~ ( n3566 ) ;
assign n3568 =  ( n3519 ) | ( n3531 )  ;
assign n3569 =  ( n3568 ) | ( n3547 )  ;
assign n3570 =  ( n3569 ) ^ ( n3564 )  ;
assign n3571 = ~ ( n3570 ) ;
assign n3572 =  ( n3189 ) ^ ( n3199 )  ;
assign n3573 =  ( n3572 ) ^ ( n3255 )  ;
assign n3574 =  ( n3573 ) ^ ( n2763 )  ;
assign n3575 =  ( n3574 ) ^ ( n2779 )  ;
assign n3576 =  ( n3575 ) ^ ( n2796 )  ;
assign n3577 =  ( n3576 ) ^ ( n2813 )  ;
assign n3578 =  ( n3577 ) ^ ( n2842 )  ;
assign n3579 =  ( n3578 ) ^ ( n2873 )  ;
assign n3580 =  ( n3579 ) ^ ( n2889 )  ;
assign n3581 =  ( n3580 ) ^ ( n2915 )  ;
assign n3582 = ~ ( n3581 ) ;
assign n3583 =  ( n3571 ) | ( n3582 )  ;
assign n3584 = ~ ( n3583 ) ;
assign n3585 =  ( n3567 ) | ( n3584 )  ;
assign n3586 = ~ ( n3585 ) ;
assign n3587 =  ( n3264 ) | ( n3274 )  ;
assign n3588 =  ( n3587 ) | ( n3288 )  ;
assign n3589 =  ( n3588 ) ^ ( n3303 )  ;
assign n3590 =  ( n3589 ) ^ ( n2846 )  ;
assign n3591 =  ( n3590 ) ^ ( n2856 )  ;
assign n3592 =  ( n3591 ) ^ ( n2919 )  ;
assign n3593 = ~ ( n2468 ) ;
assign n3594 =  ( n3592 ) ^ ( n3593 )  ;
assign n3595 =  ( n3594 ) ^ ( n2483 )  ;
assign n3596 =  ( n3595 ) ^ ( n2500 )  ;
assign n3597 =  ( n3596 ) ^ ( n2517 )  ;
assign n3598 =  ( n3597 ) ^ ( n2548 )  ;
assign n3599 =  ( n3598 ) ^ ( n2578 )  ;
assign n3600 =  ( n3599 ) ^ ( n2594 )  ;
assign n3601 =  ( n3600 ) ^ ( n2620 )  ;
assign n3602 = ~ ( n3601 ) ;
assign n3603 =  ( n3586 ) | ( n3602 )  ;
assign n3604 = ~ ( n3603 ) ;
assign n3605 = ~ ( n3583 ) ;
assign n3606 =  ( n3567 ) | ( n3605 )  ;
assign n3607 =  ( n3264 ) | ( n3274 )  ;
assign n3608 =  ( n3607 ) | ( n3288 )  ;
assign n3609 =  ( n3606 ) ^ ( n3608 )  ;
assign n3610 =  ( n3609 ) ^ ( n3303 )  ;
assign n3611 =  ( n3610 ) ^ ( n2846 )  ;
assign n3612 =  ( n3611 ) ^ ( n2856 )  ;
assign n3613 =  ( n3612 ) ^ ( n2919 )  ;
assign n3614 = ~ ( n2468 ) ;
assign n3615 =  ( n3613 ) ^ ( n3614 )  ;
assign n3616 =  ( n3615 ) ^ ( n2483 )  ;
assign n3617 =  ( n3616 ) ^ ( n2500 )  ;
assign n3618 =  ( n3617 ) ^ ( n2517 )  ;
assign n3619 =  ( n3618 ) ^ ( n2548 )  ;
assign n3620 =  ( n3619 ) ^ ( n2578 )  ;
assign n3621 =  ( n3620 ) ^ ( n2594 )  ;
assign n3622 =  ( n3621 ) ^ ( n2620 )  ;
assign n3623 =  ( n3604 ) | ( n3622 )  ;
assign n3624 = ~ ( n3623 ) ;
assign n3625 =  ( n3393 ) | ( n3624 )  ;
assign n3626 = ~ ( n3323 ) ;
assign n3627 =  ( n3306 ) | ( n3626 )  ;
assign n3628 =  ( bv_1_1_n5 ) ^ ( n3627 )  ;
assign n3629 = ~ ( n2928 ) ;
assign n3630 = ~ ( n2939 ) ;
assign n3631 =  ( n3629 ) | ( n3630 )  ;
assign n3632 = ~ ( n2954 ) ;
assign n3633 =  ( n3631 ) | ( n3632 )  ;
assign n3634 =  ( n3628 ) ^ ( n3633 )  ;
assign n3635 =  ( n3634 ) ^ ( n2971 )  ;
assign n3636 =  ( n3635 ) ^ ( n2552 )  ;
assign n3637 =  ( n3636 ) ^ ( n2561 )  ;
assign n3638 =  ( n3637 ) ^ ( n2624 )  ;
assign n3639 =  ( n3638 ) ^ ( n2144 )  ;
assign n3640 =  ( n3639 ) ^ ( n2160 )  ;
assign n3641 =  ( n3640 ) ^ ( n2177 )  ;
assign n3642 =  ( n3641 ) ^ ( n2194 )  ;
assign n3643 =  ( n3642 ) ^ ( n2223 )  ;
assign n3644 =  ( n3643 ) ^ ( n2263 )  ;
assign n3645 =  ( n3644 ) ^ ( n2309 )  ;
assign n3646 = ~ ( n3645 ) ;
assign n3647 =  ( n3625 ) | ( n3646 )  ;
assign n3648 = ~ ( n3647 ) ;
assign n3649 =  ( n3367 ) | ( n3648 )  ;
assign n3650 = ~ ( n3392 ) ;
assign n3651 =  ( bv_1_1_n5 ) ^ ( n3623 )  ;
assign n3652 = ~ ( n3323 ) ;
assign n3653 =  ( n3306 ) | ( n3652 )  ;
assign n3654 =  ( n3651 ) ^ ( n3653 )  ;
assign n3655 = ~ ( n2928 ) ;
assign n3656 = ~ ( n2939 ) ;
assign n3657 =  ( n3655 ) | ( n3656 )  ;
assign n3658 = ~ ( n2954 ) ;
assign n3659 =  ( n3657 ) | ( n3658 )  ;
assign n3660 =  ( n3654 ) ^ ( n3659 )  ;
assign n3661 =  ( n3660 ) ^ ( n2971 )  ;
assign n3662 =  ( n3661 ) ^ ( n2552 )  ;
assign n3663 =  ( n3662 ) ^ ( n2561 )  ;
assign n3664 =  ( n3663 ) ^ ( n2624 )  ;
assign n3665 =  ( n3664 ) ^ ( n2144 )  ;
assign n3666 =  ( n3665 ) ^ ( n2160 )  ;
assign n3667 =  ( n3666 ) ^ ( n2177 )  ;
assign n3668 =  ( n3667 ) ^ ( n2194 )  ;
assign n3669 =  ( n3668 ) ^ ( n2223 )  ;
assign n3670 =  ( n3669 ) ^ ( n2263 )  ;
assign n3671 =  ( n3670 ) ^ ( n2309 )  ;
assign n3672 = ~ ( n3671 ) ;
assign n3673 =  ( n3650 ) | ( n3672 )  ;
assign n3674 = ki[0:0] ;
assign n3675 =  ( n3674 ) == ( bv_1_1_n5 )  ;
assign n3676 = ki[1:1] ;
assign n3677 =  ( n3676 ) == ( bv_1_0_n2 )  ;
assign n3678 =  ( n3675 ) | ( n3677 )  ;
assign n3679 = ki[1:1] ;
assign n3680 =  ( n3679 ) == ( bv_1_1_n5 )  ;
assign n3681 = ki[0:0] ;
assign n3682 =  ( n3681 ) == ( bv_1_1_n5 )  ;
assign n3683 =  ( n3680 ) | ( n3682 )  ;
assign n3684 = ki[1:1] ;
assign n3685 =  ( n3684 ) == ( bv_1_1_n5 )  ;
assign n3686 = i_wb_data[11:11] ;
assign n3687 = ~ ( n3686 ) ;
assign n3688 = sp[11:11] ;
assign n3689 =  ( n3687 ) ^ ( n3688 )  ;
assign n3690 =  ( n3689 ) ^ ( n423 )  ;
assign n3691 =  ( n3685 ) ? ( n648 ) : ( n3690 ) ;
assign n3692 =  ( n3683 ) ? ( n3691 ) : ( bv_1_0_n2 ) ;
assign n3693 =  ( n3678 ) ? ( n3412 ) : ( n3692 ) ;
assign n3694 = ~ ( n3693 ) ;
assign n3695 =  ( n2120 ) | ( n2129 )  ;
assign n3696 =  ( n1838 ) | ( n1847 )  ;
assign n3697 = ki[3:3] ;
assign n3698 =  ( n3697 ) == ( bv_1_0_n2 )  ;
assign n3699 =  ( n3698 ) | ( n1856 )  ;
assign n3700 = i_wb_data[9:9] ;
assign n3701 = ~ ( n3700 ) ;
assign n3702 = sp[9:9] ;
assign n3703 =  ( n3701 ) ^ ( n3702 )  ;
assign n3704 =  ( n3703 ) ^ ( n734 )  ;
assign n3705 =  ( n3699 ) ? ( n3704 ) : ( n985 ) ;
assign n3706 =  ( n3696 ) ? ( bv_1_0_n2 ) : ( n3705 ) ;
assign n3707 =  ( n1838 ) | ( n1847 )  ;
assign n3708 =  ( n3707 ) ? ( bv_1_0_n2 ) : ( n3425 ) ;
assign n3709 =  ( n3695 ) ? ( n3706 ) : ( n3708 ) ;
assign n3710 = ~ ( n3709 ) ;
assign n3711 =  ( n3694 ) | ( n3710 )  ;
assign n3712 =  ( n1456 ) | ( n1465 )  ;
assign n3713 =  ( n1475 ) | ( n1484 )  ;
assign n3714 = ki[5:5] ;
assign n3715 =  ( n3714 ) == ( bv_1_0_n2 )  ;
assign n3716 =  ( n3715 ) | ( n1493 )  ;
assign n3717 = i_wb_data[7:7] ;
assign n3718 = ~ ( n3717 ) ;
assign n3719 = sp[7:7] ;
assign n3720 =  ( n3718 ) ^ ( n3719 )  ;
assign n3721 =  ( n3720 ) ^ ( n330 )  ;
assign n3722 =  ( n3716 ) ? ( n3721 ) : ( n1035 ) ;
assign n3723 =  ( n3713 ) ? ( bv_1_0_n2 ) : ( n3722 ) ;
assign n3724 =  ( n1475 ) | ( n1484 )  ;
assign n3725 =  ( n3724 ) ? ( bv_1_0_n2 ) : ( n3442 ) ;
assign n3726 =  ( n3712 ) ? ( n3723 ) : ( n3725 ) ;
assign n3727 = ~ ( n3726 ) ;
assign n3728 =  ( n3711 ) | ( n3727 )  ;
assign n3729 =  ( n1257 ) | ( n1266 )  ;
assign n3730 =  ( n873 ) | ( n882 )  ;
assign n3731 = ki[7:7] ;
assign n3732 =  ( n3731 ) == ( bv_1_0_n2 )  ;
assign n3733 =  ( n3732 ) | ( n891 )  ;
assign n3734 = i_wb_data[5:5] ;
assign n3735 = ~ ( n3734 ) ;
assign n3736 = sp[5:5] ;
assign n3737 =  ( n3735 ) ^ ( n3736 )  ;
assign n3738 =  ( n3737 ) ^ ( n241 )  ;
assign n3739 =  ( n3733 ) ? ( n3738 ) : ( n2013 ) ;
assign n3740 =  ( n3730 ) ? ( bv_1_0_n2 ) : ( n3739 ) ;
assign n3741 =  ( n873 ) | ( n882 )  ;
assign n3742 =  ( n3741 ) ? ( bv_1_0_n2 ) : ( n3459 ) ;
assign n3743 =  ( n3729 ) ? ( n3740 ) : ( n3742 ) ;
assign n3744 = ~ ( n3743 ) ;
assign n3745 =  ( n3728 ) | ( n3744 )  ;
assign n3746 = ~ ( n3745 ) ;
assign n3747 =  ( n3693 ) ^ ( n3709 )  ;
assign n3748 = ~ ( n3747 ) ;
assign n3749 =  ( n3726 ) ^ ( n3743 )  ;
assign n3750 = ~ ( n3749 ) ;
assign n3751 =  ( n3748 ) | ( n3750 )  ;
assign n3752 = ~ ( n3751 ) ;
assign n3753 =  ( n3746 ) | ( n3752 )  ;
assign n3754 =  ( n3693 ) ^ ( n3709 )  ;
assign n3755 =  ( n3754 ) ^ ( n3726 )  ;
assign n3756 =  ( n3755 ) ^ ( n3743 )  ;
assign n3757 = ~ ( n3756 ) ;
assign n3758 =  ( n908 ) | ( n917 )  ;
assign n3759 =  ( n532 ) | ( n541 )  ;
assign n3760 = ki[9:9] ;
assign n3761 =  ( n3760 ) == ( bv_1_0_n2 )  ;
assign n3762 =  ( n3761 ) | ( n550 )  ;
assign n3763 = i_wb_data[3:3] ;
assign n3764 = ~ ( n3763 ) ;
assign n3765 = sp[3:3] ;
assign n3766 =  ( n3764 ) ^ ( n3765 )  ;
assign n3767 =  ( n3766 ) ^ ( n326 )  ;
assign n3768 =  ( n3762 ) ? ( n3767 ) : ( n2306 ) ;
assign n3769 =  ( n3759 ) ? ( bv_1_0_n2 ) : ( n3768 ) ;
assign n3770 =  ( n532 ) | ( n541 )  ;
assign n3771 =  ( n3770 ) ? ( bv_1_0_n2 ) : ( n3488 ) ;
assign n3772 =  ( n3758 ) ? ( n3769 ) : ( n3771 ) ;
assign n3773 = ~ ( n3772 ) ;
assign n3774 =  ( n3757 ) | ( n3773 )  ;
assign n3775 = ~ ( n3774 ) ;
assign n3776 =  ( n3753 ) | ( n3775 )  ;
assign n3777 = ~ ( n3776 ) ;
assign n3778 = ~ ( n3693 ) ;
assign n3779 = ~ ( n3709 ) ;
assign n3780 =  ( n3778 ) | ( n3779 )  ;
assign n3781 = ~ ( n3780 ) ;
assign n3782 = ~ ( n3726 ) ;
assign n3783 = ~ ( n3743 ) ;
assign n3784 =  ( n3782 ) | ( n3783 )  ;
assign n3785 = ~ ( n3784 ) ;
assign n3786 =  ( n3781 ) | ( n3785 )  ;
assign n3787 = ~ ( n3786 ) ;
assign n3788 =  ( n3777 ) | ( n3787 )  ;
assign n3789 =  ( n567 ) | ( n576 )  ;
assign n3790 =  ( n586 ) | ( n595 )  ;
assign n3791 = ki[11:11] ;
assign n3792 =  ( n3791 ) == ( bv_1_0_n2 )  ;
assign n3793 =  ( n3792 ) | ( n604 )  ;
assign n3794 = i_wb_data[1:1] ;
assign n3795 = ~ ( n3794 ) ;
assign n3796 = sp[1:1] ;
assign n3797 =  ( n3795 ) ^ ( n3796 )  ;
assign n3798 =  ( n3797 ) ^ ( n237 )  ;
assign n3799 =  ( n3793 ) ? ( n3798 ) : ( n2615 ) ;
assign n3800 =  ( n3790 ) ? ( bv_1_0_n2 ) : ( n3799 ) ;
assign n3801 =  ( n586 ) | ( n595 )  ;
assign n3802 = ki[11:11] ;
assign n3803 =  ( n3802 ) == ( bv_1_0_n2 )  ;
assign n3804 =  ( n3803 ) | ( n604 )  ;
assign n3805 = i_wb_data[2:2] ;
assign n3806 = ~ ( n3805 ) ;
assign n3807 = sp[2:2] ;
assign n3808 =  ( n3806 ) ^ ( n3807 )  ;
assign n3809 =  ( n3808 ) ^ ( n2282 )  ;
assign n3810 =  ( n3804 ) ? ( n3809 ) : ( n2289 ) ;
assign n3811 =  ( n3801 ) ? ( bv_1_0_n2 ) : ( n3810 ) ;
assign n3812 =  ( n3789 ) ? ( n3800 ) : ( n3811 ) ;
assign n3813 = ~ ( n3812 ) ;
assign n3814 =  ( n11 ) | ( n20 )  ;
assign n3815 = ki[13:13] ;
assign n3816 = ~ ( n3815 ) ;
assign n3817 = ki[12:12] ;
assign n3818 = ~ ( n3817 ) ;
assign n3819 = ki[11:11] ;
assign n3820 = ~ ( n3819 ) ;
assign n3821 =  ( n3818 ) | ( n3820 )  ;
assign n3822 = ~ ( n3821 ) ;
assign n3823 =  ( n3816 ) | ( n3822 )  ;
assign n3824 = ~ ( n3823 ) ;
assign n3825 =  ( n30 ) | ( n39 )  ;
assign n3826 = ki[13:13] ;
assign n3827 =  ( n3826 ) == ( bv_1_0_n2 )  ;
assign n3828 =  ( n3827 ) | ( n48 )  ;
assign n3829 = i_wb_data[0:0] ;
assign n3830 = ~ ( n3829 ) ;
assign n3831 =  ( bv_1_1_n5 ) ^ ( n3830 )  ;
assign n3832 = sp[0:0] ;
assign n3833 =  ( n3831 ) ^ ( n3832 )  ;
assign n3834 =  ( n3828 ) ? ( n3833 ) : ( n2910 ) ;
assign n3835 =  ( n3825 ) ? ( bv_1_0_n2 ) : ( n3834 ) ;
assign n3836 =  ( n3814 ) ? ( n3824 ) : ( n3835 ) ;
assign n3837 = ~ ( n3836 ) ;
assign n3838 =  ( n3813 ) | ( n3837 )  ;
assign n3839 = ~ ( n3838 ) ;
assign n3840 =  ( n3812 ) ^ ( n3836 )  ;
assign n3841 = ~ ( n3840 ) ;
assign n3842 = ki[13:13] ;
assign n3843 = ~ ( n3842 ) ;
assign n3844 =  ( n3841 ) | ( n3843 )  ;
assign n3845 =  ( n3844 ) | ( n3822 )  ;
assign n3846 = ~ ( n3845 ) ;
assign n3847 =  ( n3839 ) | ( n3846 )  ;
assign n3848 = ~ ( n3847 ) ;
assign n3849 =  ( n3788 ) | ( n3848 )  ;
assign n3850 =  ( n3413 ) ^ ( n3429 )  ;
assign n3851 =  ( n3850 ) ^ ( n3446 )  ;
assign n3852 =  ( n3851 ) ^ ( n3463 )  ;
assign n3853 =  ( n3852 ) ^ ( n3492 )  ;
assign n3854 = ~ ( n3853 ) ;
assign n3855 =  ( n3849 ) | ( n3854 )  ;
assign n3856 = ~ ( n3855 ) ;
assign n3857 =  ( n3776 ) ^ ( n3786 )  ;
assign n3858 = ~ ( n3857 ) ;
assign n3859 =  ( n3847 ) ^ ( n3413 )  ;
assign n3860 =  ( n3859 ) ^ ( n3429 )  ;
assign n3861 =  ( n3860 ) ^ ( n3446 )  ;
assign n3862 =  ( n3861 ) ^ ( n3463 )  ;
assign n3863 =  ( n3862 ) ^ ( n3492 )  ;
assign n3864 = ~ ( n3863 ) ;
assign n3865 =  ( n3858 ) | ( n3864 )  ;
assign n3866 = ~ ( n3865 ) ;
assign n3867 =  ( n3856 ) | ( n3866 )  ;
assign n3868 =  ( n3776 ) ^ ( n3786 )  ;
assign n3869 =  ( n3868 ) ^ ( n3847 )  ;
assign n3870 =  ( n3869 ) ^ ( n3413 )  ;
assign n3871 =  ( n3870 ) ^ ( n3429 )  ;
assign n3872 =  ( n3871 ) ^ ( n3446 )  ;
assign n3873 =  ( n3872 ) ^ ( n3463 )  ;
assign n3874 =  ( n3873 ) ^ ( n3492 )  ;
assign n3875 = ~ ( n3874 ) ;
assign n3876 =  ( n567 ) | ( n576 )  ;
assign n3877 =  ( n586 ) | ( n595 )  ;
assign n3878 =  ( n3877 ) ? ( bv_1_0_n2 ) : ( n3810 ) ;
assign n3879 =  ( n586 ) | ( n595 )  ;
assign n3880 =  ( n3879 ) ? ( bv_1_0_n2 ) : ( n3212 ) ;
assign n3881 =  ( n3876 ) ? ( n3878 ) : ( n3880 ) ;
assign n3882 = ~ ( n3881 ) ;
assign n3883 =  ( n3875 ) | ( n3882 )  ;
assign n3884 = ~ ( n3883 ) ;
assign n3885 =  ( n3867 ) | ( n3884 )  ;
assign n3886 = ~ ( n3885 ) ;
assign n3887 = ~ ( n3776 ) ;
assign n3888 = ~ ( n3786 ) ;
assign n3889 =  ( n3887 ) | ( n3888 )  ;
assign n3890 = ~ ( n3889 ) ;
assign n3891 = ~ ( n3847 ) ;
assign n3892 =  ( n3413 ) ^ ( n3429 )  ;
assign n3893 =  ( n3892 ) ^ ( n3446 )  ;
assign n3894 =  ( n3893 ) ^ ( n3463 )  ;
assign n3895 =  ( n3894 ) ^ ( n3492 )  ;
assign n3896 = ~ ( n3895 ) ;
assign n3897 =  ( n3891 ) | ( n3896 )  ;
assign n3898 = ~ ( n3897 ) ;
assign n3899 =  ( n3890 ) | ( n3898 )  ;
assign n3900 = ~ ( n3899 ) ;
assign n3901 =  ( n3886 ) | ( n3900 )  ;
assign n3902 = ~ ( n3901 ) ;
assign n3903 =  ( n3856 ) | ( n3866 )  ;
assign n3904 =  ( n3903 ) | ( n3884 )  ;
assign n3905 =  ( n3904 ) ^ ( n3899 )  ;
assign n3906 = ~ ( n3905 ) ;
assign n3907 =  ( n3496 ) ^ ( n3506 )  ;
assign n3908 =  ( n3907 ) ^ ( n3106 )  ;
assign n3909 =  ( n3908 ) ^ ( n3122 )  ;
assign n3910 =  ( n3909 ) ^ ( n3139 )  ;
assign n3911 =  ( n3910 ) ^ ( n3156 )  ;
assign n3912 =  ( n3911 ) ^ ( n3185 )  ;
assign n3913 =  ( n3912 ) ^ ( n3216 )  ;
assign n3914 =  ( n3913 ) ^ ( n3232 )  ;
assign n3915 =  ( n3914 ) ^ ( n3251 )  ;
assign n3916 =  ( n3915 ) ^ ( n3248 )  ;
assign n3917 = ~ ( n3916 ) ;
assign n3918 =  ( n3906 ) | ( n3917 )  ;
assign n3919 = ~ ( n3918 ) ;
assign n3920 =  ( n3902 ) | ( n3919 )  ;
assign n3921 = ~ ( n3920 ) ;
assign n3922 =  ( n3519 ) | ( n3531 )  ;
assign n3923 =  ( n3922 ) | ( n3547 )  ;
assign n3924 =  ( n3923 ) ^ ( n3564 )  ;
assign n3925 =  ( n3924 ) ^ ( n3189 )  ;
assign n3926 =  ( n3925 ) ^ ( n3199 )  ;
assign n3927 =  ( n3926 ) ^ ( n3255 )  ;
assign n3928 =  ( n3927 ) ^ ( n2763 )  ;
assign n3929 =  ( n3928 ) ^ ( n2779 )  ;
assign n3930 =  ( n3929 ) ^ ( n2796 )  ;
assign n3931 =  ( n3930 ) ^ ( n2813 )  ;
assign n3932 =  ( n3931 ) ^ ( n2842 )  ;
assign n3933 =  ( n3932 ) ^ ( n2873 )  ;
assign n3934 =  ( n3933 ) ^ ( n2889 )  ;
assign n3935 =  ( n3934 ) ^ ( n2915 )  ;
assign n3936 = ~ ( n3935 ) ;
assign n3937 =  ( n3921 ) | ( n3936 )  ;
assign n3938 = ~ ( n3583 ) ;
assign n3939 =  ( n3567 ) | ( n3938 )  ;
assign n3940 =  ( bv_1_1_n5 ) ^ ( n3939 )  ;
assign n3941 =  ( n3264 ) | ( n3274 )  ;
assign n3942 =  ( n3941 ) | ( n3288 )  ;
assign n3943 =  ( n3940 ) ^ ( n3942 )  ;
assign n3944 =  ( n3943 ) ^ ( n3303 )  ;
assign n3945 =  ( n3944 ) ^ ( n2846 )  ;
assign n3946 =  ( n3945 ) ^ ( n2856 )  ;
assign n3947 =  ( n3946 ) ^ ( n2919 )  ;
assign n3948 = ~ ( n2468 ) ;
assign n3949 =  ( n3947 ) ^ ( n3948 )  ;
assign n3950 =  ( n3949 ) ^ ( n2483 )  ;
assign n3951 =  ( n3950 ) ^ ( n2500 )  ;
assign n3952 =  ( n3951 ) ^ ( n2517 )  ;
assign n3953 =  ( n3952 ) ^ ( n2548 )  ;
assign n3954 =  ( n3953 ) ^ ( n2578 )  ;
assign n3955 =  ( n3954 ) ^ ( n2594 )  ;
assign n3956 =  ( n3955 ) ^ ( n2620 )  ;
assign n3957 = ~ ( n3956 ) ;
assign n3958 =  ( n3937 ) | ( n3957 )  ;
assign n3959 = ~ ( n3958 ) ;
assign n3960 = ~ ( n3918 ) ;
assign n3961 =  ( n3902 ) | ( n3960 )  ;
assign n3962 = ~ ( n3961 ) ;
assign n3963 =  ( n3962 ) | ( n3936 )  ;
assign n3964 = ~ ( n3963 ) ;
assign n3965 =  ( bv_1_1_n5 ) ^ ( n3964 )  ;
assign n3966 = ~ ( n3583 ) ;
assign n3967 =  ( n3567 ) | ( n3966 )  ;
assign n3968 =  ( n3965 ) ^ ( n3967 )  ;
assign n3969 =  ( n3264 ) | ( n3274 )  ;
assign n3970 =  ( n3969 ) | ( n3288 )  ;
assign n3971 =  ( n3968 ) ^ ( n3970 )  ;
assign n3972 =  ( n3971 ) ^ ( n3303 )  ;
assign n3973 =  ( n3972 ) ^ ( n2846 )  ;
assign n3974 =  ( n3973 ) ^ ( n2856 )  ;
assign n3975 =  ( n3974 ) ^ ( n2919 )  ;
assign n3976 = ~ ( n2468 ) ;
assign n3977 =  ( n3975 ) ^ ( n3976 )  ;
assign n3978 =  ( n3977 ) ^ ( n2483 )  ;
assign n3979 =  ( n3978 ) ^ ( n2500 )  ;
assign n3980 =  ( n3979 ) ^ ( n2517 )  ;
assign n3981 =  ( n3980 ) ^ ( n2548 )  ;
assign n3982 =  ( n3981 ) ^ ( n2578 )  ;
assign n3983 =  ( n3982 ) ^ ( n2594 )  ;
assign n3984 =  ( n3983 ) ^ ( n2620 )  ;
assign n3985 = ~ ( n3984 ) ;
assign n3986 = ki[0:0] ;
assign n3987 =  ( n3986 ) == ( bv_1_1_n5 )  ;
assign n3988 = ki[1:1] ;
assign n3989 =  ( n3988 ) == ( bv_1_0_n2 )  ;
assign n3990 =  ( n3987 ) | ( n3989 )  ;
assign n3991 = ki[1:1] ;
assign n3992 =  ( n3991 ) == ( bv_1_1_n5 )  ;
assign n3993 = ki[0:0] ;
assign n3994 =  ( n3993 ) == ( bv_1_1_n5 )  ;
assign n3995 =  ( n3992 ) | ( n3994 )  ;
assign n3996 = ki[1:1] ;
assign n3997 =  ( n3996 ) == ( bv_1_1_n5 )  ;
assign n3998 = i_wb_data[10:10] ;
assign n3999 = ~ ( n3998 ) ;
assign n4000 = sp[10:10] ;
assign n4001 =  ( n3999 ) ^ ( n4000 )  ;
assign n4002 =  ( n4001 ) ^ ( n738 )  ;
assign n4003 =  ( n3997 ) ? ( n745 ) : ( n4002 ) ;
assign n4004 =  ( n3995 ) ? ( n4003 ) : ( bv_1_0_n2 ) ;
assign n4005 =  ( n3990 ) ? ( n3692 ) : ( n4004 ) ;
assign n4006 = ~ ( n4005 ) ;
assign n4007 =  ( n2120 ) | ( n2129 )  ;
assign n4008 =  ( n1838 ) | ( n1847 )  ;
assign n4009 = ki[3:3] ;
assign n4010 =  ( n4009 ) == ( bv_1_0_n2 )  ;
assign n4011 =  ( n4010 ) | ( n1856 )  ;
assign n4012 = i_wb_data[8:8] ;
assign n4013 = ~ ( n4012 ) ;
assign n4014 = sp[8:8] ;
assign n4015 =  ( n4013 ) ^ ( n4014 )  ;
assign n4016 =  ( n4015 ) ^ ( n1054 )  ;
assign n4017 =  ( n4011 ) ? ( n4016 ) : ( n1061 ) ;
assign n4018 =  ( n4008 ) ? ( bv_1_0_n2 ) : ( n4017 ) ;
assign n4019 =  ( n1838 ) | ( n1847 )  ;
assign n4020 =  ( n4019 ) ? ( bv_1_0_n2 ) : ( n3705 ) ;
assign n4021 =  ( n4007 ) ? ( n4018 ) : ( n4020 ) ;
assign n4022 = ~ ( n4021 ) ;
assign n4023 =  ( n4006 ) | ( n4022 )  ;
assign n4024 =  ( n1456 ) | ( n1465 )  ;
assign n4025 =  ( n1475 ) | ( n1484 )  ;
assign n4026 = ki[5:5] ;
assign n4027 =  ( n4026 ) == ( bv_1_0_n2 )  ;
assign n4028 =  ( n4027 ) | ( n1493 )  ;
assign n4029 = i_wb_data[6:6] ;
assign n4030 = ~ ( n4029 ) ;
assign n4031 = sp[6:6] ;
assign n4032 =  ( n4030 ) ^ ( n4031 )  ;
assign n4033 =  ( n4032 ) ^ ( n1363 )  ;
assign n4034 =  ( n4028 ) ? ( n4033 ) : ( n1370 ) ;
assign n4035 =  ( n4025 ) ? ( bv_1_0_n2 ) : ( n4034 ) ;
assign n4036 =  ( n1475 ) | ( n1484 )  ;
assign n4037 =  ( n4036 ) ? ( bv_1_0_n2 ) : ( n3722 ) ;
assign n4038 =  ( n4024 ) ? ( n4035 ) : ( n4037 ) ;
assign n4039 = ~ ( n4038 ) ;
assign n4040 =  ( n4023 ) | ( n4039 )  ;
assign n4041 =  ( n1257 ) | ( n1266 )  ;
assign n4042 =  ( n873 ) | ( n882 )  ;
assign n4043 = ki[7:7] ;
assign n4044 =  ( n4043 ) == ( bv_1_0_n2 )  ;
assign n4045 =  ( n4044 ) | ( n891 )  ;
assign n4046 = i_wb_data[4:4] ;
assign n4047 = ~ ( n4046 ) ;
assign n4048 = sp[4:4] ;
assign n4049 =  ( n4047 ) ^ ( n4048 )  ;
assign n4050 =  ( n4049 ) ^ ( n1989 )  ;
assign n4051 =  ( n4045 ) ? ( n4050 ) : ( n1996 ) ;
assign n4052 =  ( n4042 ) ? ( bv_1_0_n2 ) : ( n4051 ) ;
assign n4053 =  ( n873 ) | ( n882 )  ;
assign n4054 =  ( n4053 ) ? ( bv_1_0_n2 ) : ( n3739 ) ;
assign n4055 =  ( n4041 ) ? ( n4052 ) : ( n4054 ) ;
assign n4056 = ~ ( n4055 ) ;
assign n4057 =  ( n4040 ) | ( n4056 )  ;
assign n4058 = ~ ( n4057 ) ;
assign n4059 =  ( n4005 ) ^ ( n4021 )  ;
assign n4060 = ~ ( n4059 ) ;
assign n4061 =  ( n4038 ) ^ ( n4055 )  ;
assign n4062 = ~ ( n4061 ) ;
assign n4063 =  ( n4060 ) | ( n4062 )  ;
assign n4064 = ~ ( n4063 ) ;
assign n4065 =  ( n4058 ) | ( n4064 )  ;
assign n4066 =  ( n4005 ) ^ ( n4021 )  ;
assign n4067 =  ( n4066 ) ^ ( n4038 )  ;
assign n4068 =  ( n4067 ) ^ ( n4055 )  ;
assign n4069 = ~ ( n4068 ) ;
assign n4070 =  ( n908 ) | ( n917 )  ;
assign n4071 =  ( n532 ) | ( n541 )  ;
assign n4072 = ki[9:9] ;
assign n4073 =  ( n4072 ) == ( bv_1_0_n2 )  ;
assign n4074 =  ( n4073 ) | ( n550 )  ;
assign n4075 = i_wb_data[2:2] ;
assign n4076 = ~ ( n4075 ) ;
assign n4077 = sp[2:2] ;
assign n4078 =  ( n4076 ) ^ ( n4077 )  ;
assign n4079 =  ( n4078 ) ^ ( n2282 )  ;
assign n4080 =  ( n4074 ) ? ( n4079 ) : ( n2289 ) ;
assign n4081 =  ( n4071 ) ? ( bv_1_0_n2 ) : ( n4080 ) ;
assign n4082 =  ( n532 ) | ( n541 )  ;
assign n4083 =  ( n4082 ) ? ( bv_1_0_n2 ) : ( n3768 ) ;
assign n4084 =  ( n4070 ) ? ( n4081 ) : ( n4083 ) ;
assign n4085 = ~ ( n4084 ) ;
assign n4086 =  ( n4069 ) | ( n4085 )  ;
assign n4087 = ~ ( n4086 ) ;
assign n4088 =  ( n4065 ) | ( n4087 )  ;
assign n4089 = ~ ( n4088 ) ;
assign n4090 = ~ ( n4005 ) ;
assign n4091 = ~ ( n4021 ) ;
assign n4092 =  ( n4090 ) | ( n4091 )  ;
assign n4093 = ~ ( n4092 ) ;
assign n4094 = ~ ( n4038 ) ;
assign n4095 = ~ ( n4055 ) ;
assign n4096 =  ( n4094 ) | ( n4095 )  ;
assign n4097 = ~ ( n4096 ) ;
assign n4098 =  ( n4093 ) | ( n4097 )  ;
assign n4099 = ~ ( n4098 ) ;
assign n4100 =  ( n4089 ) | ( n4099 )  ;
assign n4101 = ~ ( n4100 ) ;
assign n4102 =  ( n4088 ) ^ ( n4098 )  ;
assign n4103 = ~ ( n4102 ) ;
assign n4104 =  ( n3693 ) ^ ( n3709 )  ;
assign n4105 =  ( n4104 ) ^ ( n3726 )  ;
assign n4106 =  ( n4105 ) ^ ( n3743 )  ;
assign n4107 =  ( n4106 ) ^ ( n3772 )  ;
assign n4108 = ~ ( n4107 ) ;
assign n4109 =  ( n4103 ) | ( n4108 )  ;
assign n4110 = ~ ( n4109 ) ;
assign n4111 =  ( n4101 ) | ( n4110 )  ;
assign n4112 = ~ ( n4111 ) ;
assign n4113 =  ( n3776 ) ^ ( n3786 )  ;
assign n4114 =  ( n4113 ) ^ ( n3847 )  ;
assign n4115 =  ( n4114 ) ^ ( n3413 )  ;
assign n4116 =  ( n4115 ) ^ ( n3429 )  ;
assign n4117 =  ( n4116 ) ^ ( n3446 )  ;
assign n4118 =  ( n4117 ) ^ ( n3463 )  ;
assign n4119 =  ( n4118 ) ^ ( n3492 )  ;
assign n4120 =  ( n4119 ) ^ ( n3881 )  ;
assign n4121 = ~ ( n4120 ) ;
assign n4122 =  ( n4112 ) | ( n4121 )  ;
assign n4123 = ~ ( n4122 ) ;
assign n4124 =  ( n4111 ) ^ ( n3776 )  ;
assign n4125 =  ( n4124 ) ^ ( n3786 )  ;
assign n4126 =  ( n4125 ) ^ ( n3847 )  ;
assign n4127 =  ( n4126 ) ^ ( n3413 )  ;
assign n4128 =  ( n4127 ) ^ ( n3429 )  ;
assign n4129 =  ( n4128 ) ^ ( n3446 )  ;
assign n4130 =  ( n4129 ) ^ ( n3463 )  ;
assign n4131 =  ( n4130 ) ^ ( n3492 )  ;
assign n4132 =  ( n4131 ) ^ ( n3881 )  ;
assign n4133 = ~ ( n4132 ) ;
assign n4134 =  ( n11 ) | ( n20 )  ;
assign n4135 =  ( n30 ) | ( n39 )  ;
assign n4136 =  ( n4135 ) ? ( bv_1_0_n2 ) : ( n3834 ) ;
assign n4137 =  ( n30 ) | ( n39 )  ;
assign n4138 =  ( n4137 ) ? ( bv_1_0_n2 ) : ( n3228 ) ;
assign n4139 =  ( n4134 ) ? ( n4136 ) : ( n4138 ) ;
assign n4140 = ~ ( n4139 ) ;
assign n4141 =  ( n4133 ) | ( n4140 )  ;
assign n4142 = ~ ( n4141 ) ;
assign n4143 =  ( n4123 ) | ( n4142 )  ;
assign n4144 = ~ ( n4143 ) ;
assign n4145 =  ( n3985 ) | ( n4144 )  ;
assign n4146 =  ( n3856 ) | ( n3866 )  ;
assign n4147 =  ( n4146 ) | ( n3884 )  ;
assign n4148 =  ( n4147 ) ^ ( n3899 )  ;
assign n4149 =  ( n4148 ) ^ ( n3496 )  ;
assign n4150 =  ( n4149 ) ^ ( n3506 )  ;
assign n4151 =  ( n4150 ) ^ ( n3106 )  ;
assign n4152 =  ( n4151 ) ^ ( n3122 )  ;
assign n4153 =  ( n4152 ) ^ ( n3139 )  ;
assign n4154 =  ( n4153 ) ^ ( n3156 )  ;
assign n4155 =  ( n4154 ) ^ ( n3185 )  ;
assign n4156 =  ( n4155 ) ^ ( n3216 )  ;
assign n4157 =  ( n4156 ) ^ ( n3232 )  ;
assign n4158 =  ( n4157 ) ^ ( n3251 )  ;
assign n4159 =  ( n4158 ) ^ ( n3248 )  ;
assign n4160 = ~ ( n4159 ) ;
assign n4161 =  ( n4145 ) | ( n4160 )  ;
assign n4162 = ~ ( n3918 ) ;
assign n4163 =  ( n3902 ) | ( n4162 )  ;
assign n4164 =  ( n3519 ) | ( n3531 )  ;
assign n4165 =  ( n4164 ) | ( n3547 )  ;
assign n4166 =  ( n4163 ) ^ ( n4165 )  ;
assign n4167 =  ( n4166 ) ^ ( n3564 )  ;
assign n4168 =  ( n4167 ) ^ ( n3189 )  ;
assign n4169 =  ( n4168 ) ^ ( n3199 )  ;
assign n4170 =  ( n4169 ) ^ ( n3255 )  ;
assign n4171 =  ( n4170 ) ^ ( n2763 )  ;
assign n4172 =  ( n4171 ) ^ ( n2779 )  ;
assign n4173 =  ( n4172 ) ^ ( n2796 )  ;
assign n4174 =  ( n4173 ) ^ ( n2813 )  ;
assign n4175 =  ( n4174 ) ^ ( n2842 )  ;
assign n4176 =  ( n4175 ) ^ ( n2873 )  ;
assign n4177 =  ( n4176 ) ^ ( n2889 )  ;
assign n4178 =  ( n4177 ) ^ ( n2915 )  ;
assign n4179 = ~ ( n4178 ) ;
assign n4180 =  ( n4161 ) | ( n4179 )  ;
assign n4181 = ~ ( n4180 ) ;
assign n4182 =  ( n3959 ) | ( n4181 )  ;
assign n4183 = ~ ( n4182 ) ;
assign n4184 =  ( n3673 ) | ( n4183 )  ;
assign n4185 = ~ ( n4184 ) ;
assign n4186 =  ( n3649 ) | ( n4185 )  ;
assign n4187 = ~ ( n4186 ) ;
assign n4188 =  ( n3086 ) | ( n4187 )  ;
assign n4189 = ~ ( n4188 ) ;
assign n4190 =  ( n3066 ) | ( n4189 )  ;
assign n4191 = ~ ( n4190 ) ;
assign n4192 =  ( n1829 ) | ( n4191 )  ;
assign n4193 = ~ ( n4192 ) ;
assign n4194 =  ( n1794 ) | ( n4193 )  ;
assign n4195 = ~ ( n518 ) ;
assign n4196 =  ( bv_1_1_n5 ) ^ ( n488 )  ;
assign n4197 =  ( n4196 ) ^ ( n504 )  ;
assign n4198 = ~ ( n4197 ) ;
assign n4199 =  ( n4195 ) | ( n4198 )  ;
assign n4200 = ~ ( n856 ) ;
assign n4201 =  ( n4199 ) | ( n4200 )  ;
assign n4202 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n4203 =  ( n4202 ) ^ ( n823 )  ;
assign n4204 =  ( n4203 ) ^ ( n344 )  ;
assign n4205 =  ( n4204 ) ^ ( n454 )  ;
assign n4206 = ~ ( n4205 ) ;
assign n4207 =  ( n4201 ) | ( n4206 )  ;
assign n4208 = ~ ( n1239 ) ;
assign n4209 =  ( n4207 ) | ( n4208 )  ;
assign n4210 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n4211 =  ( n4210 ) ^ ( n1199 )  ;
assign n4212 =  ( n4211 ) ^ ( n666 )  ;
assign n4213 =  ( n4212 ) ^ ( n682 )  ;
assign n4214 =  ( n4213 ) ^ ( n697 )  ;
assign n4215 =  ( n4214 ) ^ ( n759 )  ;
assign n4216 = ~ ( n4215 ) ;
assign n4217 =  ( n4209 ) | ( n4216 )  ;
assign n4218 = ~ ( n1446 ) ;
assign n4219 =  ( n4217 ) | ( n4218 )  ;
assign n4220 =  ( n4219 ) | ( n1828 )  ;
assign n4221 = ~ ( n2110 ) ;
assign n4222 =  ( n4220 ) | ( n4221 )  ;
assign n4223 =  ( n4222 ) | ( n2453 )  ;
assign n4224 = ~ ( n2742 ) ;
assign n4225 =  ( n4223 ) | ( n4224 )  ;
assign n4226 =  ( n4225 ) | ( n3085 )  ;
assign n4227 = ~ ( n3392 ) ;
assign n4228 =  ( n4226 ) | ( n4227 )  ;
assign n4229 =  ( n4228 ) | ( n3672 )  ;
assign n4230 =  ( n4229 ) | ( n3985 )  ;
assign n4231 =  ( n4123 ) | ( n4142 )  ;
assign n4232 = ~ ( n4231 ) ;
assign n4233 =  ( n4232 ) | ( n4160 )  ;
assign n4234 = ~ ( n4233 ) ;
assign n4235 = ~ ( n3918 ) ;
assign n4236 =  ( n3902 ) | ( n4235 )  ;
assign n4237 =  ( n4234 ) ^ ( n4236 )  ;
assign n4238 =  ( n3519 ) | ( n3531 )  ;
assign n4239 =  ( n4238 ) | ( n3547 )  ;
assign n4240 =  ( n4237 ) ^ ( n4239 )  ;
assign n4241 =  ( n4240 ) ^ ( n3564 )  ;
assign n4242 =  ( n4241 ) ^ ( n3189 )  ;
assign n4243 =  ( n4242 ) ^ ( n3199 )  ;
assign n4244 =  ( n4243 ) ^ ( n3255 )  ;
assign n4245 =  ( n4244 ) ^ ( n2763 )  ;
assign n4246 =  ( n4245 ) ^ ( n2779 )  ;
assign n4247 =  ( n4246 ) ^ ( n2796 )  ;
assign n4248 =  ( n4247 ) ^ ( n2813 )  ;
assign n4249 =  ( n4248 ) ^ ( n2842 )  ;
assign n4250 =  ( n4249 ) ^ ( n2873 )  ;
assign n4251 =  ( n4250 ) ^ ( n2889 )  ;
assign n4252 =  ( n4251 ) ^ ( n2915 )  ;
assign n4253 = ~ ( n4252 ) ;
assign n4254 =  ( n4230 ) | ( n4253 )  ;
assign n4255 = ki[0:0] ;
assign n4256 =  ( n4255 ) == ( bv_1_1_n5 )  ;
assign n4257 = ki[1:1] ;
assign n4258 =  ( n4257 ) == ( bv_1_0_n2 )  ;
assign n4259 =  ( n4256 ) | ( n4258 )  ;
assign n4260 = ki[1:1] ;
assign n4261 =  ( n4260 ) == ( bv_1_1_n5 )  ;
assign n4262 = ki[0:0] ;
assign n4263 =  ( n4262 ) == ( bv_1_1_n5 )  ;
assign n4264 =  ( n4261 ) | ( n4263 )  ;
assign n4265 = ki[1:1] ;
assign n4266 =  ( n4265 ) == ( bv_1_1_n5 )  ;
assign n4267 = i_wb_data[9:9] ;
assign n4268 = ~ ( n4267 ) ;
assign n4269 = sp[9:9] ;
assign n4270 =  ( n4268 ) ^ ( n4269 )  ;
assign n4271 =  ( n4270 ) ^ ( n734 )  ;
assign n4272 =  ( n4266 ) ? ( n985 ) : ( n4271 ) ;
assign n4273 =  ( n4264 ) ? ( n4272 ) : ( bv_1_0_n2 ) ;
assign n4274 =  ( n4259 ) ? ( n4004 ) : ( n4273 ) ;
assign n4275 = ~ ( n4274 ) ;
assign n4276 =  ( n2120 ) | ( n2129 )  ;
assign n4277 =  ( n1838 ) | ( n1847 )  ;
assign n4278 = ki[3:3] ;
assign n4279 =  ( n4278 ) == ( bv_1_0_n2 )  ;
assign n4280 =  ( n4279 ) | ( n1856 )  ;
assign n4281 = i_wb_data[7:7] ;
assign n4282 = ~ ( n4281 ) ;
assign n4283 = sp[7:7] ;
assign n4284 =  ( n4282 ) ^ ( n4283 )  ;
assign n4285 =  ( n4284 ) ^ ( n330 )  ;
assign n4286 =  ( n4280 ) ? ( n4285 ) : ( n1035 ) ;
assign n4287 =  ( n4277 ) ? ( bv_1_0_n2 ) : ( n4286 ) ;
assign n4288 =  ( n1838 ) | ( n1847 )  ;
assign n4289 =  ( n4288 ) ? ( bv_1_0_n2 ) : ( n4017 ) ;
assign n4290 =  ( n4276 ) ? ( n4287 ) : ( n4289 ) ;
assign n4291 = ~ ( n4290 ) ;
assign n4292 =  ( n4275 ) | ( n4291 )  ;
assign n4293 =  ( n1456 ) | ( n1465 )  ;
assign n4294 =  ( n1475 ) | ( n1484 )  ;
assign n4295 = ki[5:5] ;
assign n4296 =  ( n4295 ) == ( bv_1_0_n2 )  ;
assign n4297 =  ( n4296 ) | ( n1493 )  ;
assign n4298 = i_wb_data[5:5] ;
assign n4299 = ~ ( n4298 ) ;
assign n4300 = sp[5:5] ;
assign n4301 =  ( n4299 ) ^ ( n4300 )  ;
assign n4302 =  ( n4301 ) ^ ( n241 )  ;
assign n4303 =  ( n4297 ) ? ( n4302 ) : ( n2013 ) ;
assign n4304 =  ( n4294 ) ? ( bv_1_0_n2 ) : ( n4303 ) ;
assign n4305 =  ( n1475 ) | ( n1484 )  ;
assign n4306 =  ( n4305 ) ? ( bv_1_0_n2 ) : ( n4034 ) ;
assign n4307 =  ( n4293 ) ? ( n4304 ) : ( n4306 ) ;
assign n4308 = ~ ( n4307 ) ;
assign n4309 =  ( n4292 ) | ( n4308 )  ;
assign n4310 =  ( n1257 ) | ( n1266 )  ;
assign n4311 =  ( n873 ) | ( n882 )  ;
assign n4312 = ki[7:7] ;
assign n4313 =  ( n4312 ) == ( bv_1_0_n2 )  ;
assign n4314 =  ( n4313 ) | ( n891 )  ;
assign n4315 = i_wb_data[3:3] ;
assign n4316 = ~ ( n4315 ) ;
assign n4317 = sp[3:3] ;
assign n4318 =  ( n4316 ) ^ ( n4317 )  ;
assign n4319 =  ( n4318 ) ^ ( n326 )  ;
assign n4320 =  ( n4314 ) ? ( n4319 ) : ( n2306 ) ;
assign n4321 =  ( n4311 ) ? ( bv_1_0_n2 ) : ( n4320 ) ;
assign n4322 =  ( n873 ) | ( n882 )  ;
assign n4323 =  ( n4322 ) ? ( bv_1_0_n2 ) : ( n4051 ) ;
assign n4324 =  ( n4310 ) ? ( n4321 ) : ( n4323 ) ;
assign n4325 = ~ ( n4324 ) ;
assign n4326 =  ( n4309 ) | ( n4325 )  ;
assign n4327 = ~ ( n4326 ) ;
assign n4328 =  ( n4274 ) ^ ( n4290 )  ;
assign n4329 = ~ ( n4328 ) ;
assign n4330 =  ( n4307 ) ^ ( n4324 )  ;
assign n4331 = ~ ( n4330 ) ;
assign n4332 =  ( n4329 ) | ( n4331 )  ;
assign n4333 = ~ ( n4332 ) ;
assign n4334 =  ( n4327 ) | ( n4333 )  ;
assign n4335 =  ( n4274 ) ^ ( n4290 )  ;
assign n4336 =  ( n4335 ) ^ ( n4307 )  ;
assign n4337 =  ( n4336 ) ^ ( n4324 )  ;
assign n4338 = ~ ( n4337 ) ;
assign n4339 =  ( n908 ) | ( n917 )  ;
assign n4340 =  ( n532 ) | ( n541 )  ;
assign n4341 = ki[9:9] ;
assign n4342 =  ( n4341 ) == ( bv_1_0_n2 )  ;
assign n4343 =  ( n4342 ) | ( n550 )  ;
assign n4344 = i_wb_data[1:1] ;
assign n4345 = ~ ( n4344 ) ;
assign n4346 = sp[1:1] ;
assign n4347 =  ( n4345 ) ^ ( n4346 )  ;
assign n4348 =  ( n4347 ) ^ ( n237 )  ;
assign n4349 =  ( n4343 ) ? ( n4348 ) : ( n2615 ) ;
assign n4350 =  ( n4340 ) ? ( bv_1_0_n2 ) : ( n4349 ) ;
assign n4351 =  ( n532 ) | ( n541 )  ;
assign n4352 =  ( n4351 ) ? ( bv_1_0_n2 ) : ( n4080 ) ;
assign n4353 =  ( n4339 ) ? ( n4350 ) : ( n4352 ) ;
assign n4354 = ~ ( n4353 ) ;
assign n4355 =  ( n4338 ) | ( n4354 )  ;
assign n4356 = ~ ( n4355 ) ;
assign n4357 =  ( n4334 ) | ( n4356 )  ;
assign n4358 = ~ ( n4357 ) ;
assign n4359 = ~ ( n4274 ) ;
assign n4360 = ~ ( n4290 ) ;
assign n4361 =  ( n4359 ) | ( n4360 )  ;
assign n4362 = ~ ( n4361 ) ;
assign n4363 = ~ ( n4307 ) ;
assign n4364 = ~ ( n4324 ) ;
assign n4365 =  ( n4363 ) | ( n4364 )  ;
assign n4366 = ~ ( n4365 ) ;
assign n4367 =  ( n4362 ) | ( n4366 )  ;
assign n4368 = ~ ( n4367 ) ;
assign n4369 =  ( n4358 ) | ( n4368 )  ;
assign n4370 = ~ ( n4369 ) ;
assign n4371 =  ( n4357 ) ^ ( n4367 )  ;
assign n4372 = ~ ( n4371 ) ;
assign n4373 =  ( n4005 ) ^ ( n4021 )  ;
assign n4374 =  ( n4373 ) ^ ( n4038 )  ;
assign n4375 =  ( n4374 ) ^ ( n4055 )  ;
assign n4376 =  ( n4375 ) ^ ( n4084 )  ;
assign n4377 = ~ ( n4376 ) ;
assign n4378 =  ( n4372 ) | ( n4377 )  ;
assign n4379 = ~ ( n4378 ) ;
assign n4380 =  ( n4370 ) | ( n4379 )  ;
assign n4381 = ~ ( n4380 ) ;
assign n4382 =  ( n4088 ) ^ ( n4098 )  ;
assign n4383 =  ( n4382 ) ^ ( n3693 )  ;
assign n4384 =  ( n4383 ) ^ ( n3709 )  ;
assign n4385 =  ( n4384 ) ^ ( n3726 )  ;
assign n4386 =  ( n4385 ) ^ ( n3743 )  ;
assign n4387 =  ( n4386 ) ^ ( n3772 )  ;
assign n4388 = ~ ( n4387 ) ;
assign n4389 =  ( n4381 ) | ( n4388 )  ;
assign n4390 = ~ ( n4389 ) ;
assign n4391 =  ( n4380 ) ^ ( n4088 )  ;
assign n4392 =  ( n4391 ) ^ ( n4098 )  ;
assign n4393 =  ( n4392 ) ^ ( n3693 )  ;
assign n4394 =  ( n4393 ) ^ ( n3709 )  ;
assign n4395 =  ( n4394 ) ^ ( n3726 )  ;
assign n4396 =  ( n4395 ) ^ ( n3743 )  ;
assign n4397 =  ( n4396 ) ^ ( n3772 )  ;
assign n4398 = ~ ( n4397 ) ;
assign n4399 =  ( n3812 ) ^ ( n3836 )  ;
assign n4400 =  ( n4399 ) ^ ( n3824 )  ;
assign n4401 = ~ ( n4400 ) ;
assign n4402 =  ( n4398 ) | ( n4401 )  ;
assign n4403 = ~ ( n4402 ) ;
assign n4404 =  ( n4390 ) | ( n4403 )  ;
assign n4405 = ~ ( n4404 ) ;
assign n4406 =  ( n4111 ) ^ ( n3776 )  ;
assign n4407 =  ( n4406 ) ^ ( n3786 )  ;
assign n4408 =  ( n4407 ) ^ ( n3847 )  ;
assign n4409 =  ( n4408 ) ^ ( n3413 )  ;
assign n4410 =  ( n4409 ) ^ ( n3429 )  ;
assign n4411 =  ( n4410 ) ^ ( n3446 )  ;
assign n4412 =  ( n4411 ) ^ ( n3463 )  ;
assign n4413 =  ( n4412 ) ^ ( n3492 )  ;
assign n4414 =  ( n4413 ) ^ ( n3881 )  ;
assign n4415 =  ( n4414 ) ^ ( n4139 )  ;
assign n4416 = ~ ( n4415 ) ;
assign n4417 =  ( n4405 ) | ( n4416 )  ;
assign n4418 =  ( n4123 ) | ( n4142 )  ;
assign n4419 =  ( n3856 ) | ( n3866 )  ;
assign n4420 =  ( n4419 ) | ( n3884 )  ;
assign n4421 =  ( n4418 ) ^ ( n4420 )  ;
assign n4422 =  ( n4421 ) ^ ( n3899 )  ;
assign n4423 =  ( n4422 ) ^ ( n3496 )  ;
assign n4424 =  ( n4423 ) ^ ( n3506 )  ;
assign n4425 =  ( n4424 ) ^ ( n3106 )  ;
assign n4426 =  ( n4425 ) ^ ( n3122 )  ;
assign n4427 =  ( n4426 ) ^ ( n3139 )  ;
assign n4428 =  ( n4427 ) ^ ( n3156 )  ;
assign n4429 =  ( n4428 ) ^ ( n3185 )  ;
assign n4430 =  ( n4429 ) ^ ( n3216 )  ;
assign n4431 =  ( n4430 ) ^ ( n3232 )  ;
assign n4432 =  ( n4431 ) ^ ( n3251 )  ;
assign n4433 =  ( n4432 ) ^ ( n3248 )  ;
assign n4434 = ~ ( n4433 ) ;
assign n4435 =  ( n4417 ) | ( n4434 )  ;
assign n4436 = ~ ( n4435 ) ;
assign n4437 =  ( n4390 ) | ( n4403 )  ;
assign n4438 = ~ ( n4437 ) ;
assign n4439 =  ( n4438 ) | ( n4416 )  ;
assign n4440 = ~ ( n4439 ) ;
assign n4441 =  ( n4123 ) | ( n4142 )  ;
assign n4442 =  ( n4440 ) ^ ( n4441 )  ;
assign n4443 =  ( n3856 ) | ( n3866 )  ;
assign n4444 =  ( n4443 ) | ( n3884 )  ;
assign n4445 =  ( n4442 ) ^ ( n4444 )  ;
assign n4446 =  ( n4445 ) ^ ( n3899 )  ;
assign n4447 =  ( n4446 ) ^ ( n3496 )  ;
assign n4448 =  ( n4447 ) ^ ( n3506 )  ;
assign n4449 =  ( n4448 ) ^ ( n3106 )  ;
assign n4450 =  ( n4449 ) ^ ( n3122 )  ;
assign n4451 =  ( n4450 ) ^ ( n3139 )  ;
assign n4452 =  ( n4451 ) ^ ( n3156 )  ;
assign n4453 =  ( n4452 ) ^ ( n3185 )  ;
assign n4454 =  ( n4453 ) ^ ( n3216 )  ;
assign n4455 =  ( n4454 ) ^ ( n3232 )  ;
assign n4456 =  ( n4455 ) ^ ( n3251 )  ;
assign n4457 =  ( n4456 ) ^ ( n3248 )  ;
assign n4458 = ~ ( n4457 ) ;
assign n4459 = ki[0:0] ;
assign n4460 =  ( n4459 ) == ( bv_1_1_n5 )  ;
assign n4461 = ki[1:1] ;
assign n4462 =  ( n4461 ) == ( bv_1_0_n2 )  ;
assign n4463 =  ( n4460 ) | ( n4462 )  ;
assign n4464 = ki[1:1] ;
assign n4465 =  ( n4464 ) == ( bv_1_1_n5 )  ;
assign n4466 = ki[0:0] ;
assign n4467 =  ( n4466 ) == ( bv_1_1_n5 )  ;
assign n4468 =  ( n4465 ) | ( n4467 )  ;
assign n4469 = ki[1:1] ;
assign n4470 =  ( n4469 ) == ( bv_1_1_n5 )  ;
assign n4471 = i_wb_data[8:8] ;
assign n4472 = ~ ( n4471 ) ;
assign n4473 = sp[8:8] ;
assign n4474 =  ( n4472 ) ^ ( n4473 )  ;
assign n4475 =  ( n4474 ) ^ ( n1054 )  ;
assign n4476 =  ( n4470 ) ? ( n1061 ) : ( n4475 ) ;
assign n4477 =  ( n4468 ) ? ( n4476 ) : ( bv_1_0_n2 ) ;
assign n4478 =  ( n4463 ) ? ( n4273 ) : ( n4477 ) ;
assign n4479 = ~ ( n4478 ) ;
assign n4480 =  ( n2120 ) | ( n2129 )  ;
assign n4481 =  ( n1838 ) | ( n1847 )  ;
assign n4482 = ki[3:3] ;
assign n4483 =  ( n4482 ) == ( bv_1_0_n2 )  ;
assign n4484 =  ( n4483 ) | ( n1856 )  ;
assign n4485 = i_wb_data[6:6] ;
assign n4486 = ~ ( n4485 ) ;
assign n4487 = sp[6:6] ;
assign n4488 =  ( n4486 ) ^ ( n4487 )  ;
assign n4489 =  ( n4488 ) ^ ( n1363 )  ;
assign n4490 =  ( n4484 ) ? ( n4489 ) : ( n1370 ) ;
assign n4491 =  ( n4481 ) ? ( bv_1_0_n2 ) : ( n4490 ) ;
assign n4492 =  ( n1838 ) | ( n1847 )  ;
assign n4493 =  ( n4492 ) ? ( bv_1_0_n2 ) : ( n4286 ) ;
assign n4494 =  ( n4480 ) ? ( n4491 ) : ( n4493 ) ;
assign n4495 = ~ ( n4494 ) ;
assign n4496 =  ( n4479 ) | ( n4495 )  ;
assign n4497 =  ( n1456 ) | ( n1465 )  ;
assign n4498 =  ( n1475 ) | ( n1484 )  ;
assign n4499 = ki[5:5] ;
assign n4500 =  ( n4499 ) == ( bv_1_0_n2 )  ;
assign n4501 =  ( n4500 ) | ( n1493 )  ;
assign n4502 = i_wb_data[4:4] ;
assign n4503 = ~ ( n4502 ) ;
assign n4504 = sp[4:4] ;
assign n4505 =  ( n4503 ) ^ ( n4504 )  ;
assign n4506 =  ( n4505 ) ^ ( n1989 )  ;
assign n4507 =  ( n4501 ) ? ( n4506 ) : ( n1996 ) ;
assign n4508 =  ( n4498 ) ? ( bv_1_0_n2 ) : ( n4507 ) ;
assign n4509 =  ( n1475 ) | ( n1484 )  ;
assign n4510 =  ( n4509 ) ? ( bv_1_0_n2 ) : ( n4303 ) ;
assign n4511 =  ( n4497 ) ? ( n4508 ) : ( n4510 ) ;
assign n4512 = ~ ( n4511 ) ;
assign n4513 =  ( n4496 ) | ( n4512 )  ;
assign n4514 =  ( n1257 ) | ( n1266 )  ;
assign n4515 =  ( n873 ) | ( n882 )  ;
assign n4516 = ki[7:7] ;
assign n4517 =  ( n4516 ) == ( bv_1_0_n2 )  ;
assign n4518 =  ( n4517 ) | ( n891 )  ;
assign n4519 = i_wb_data[2:2] ;
assign n4520 = ~ ( n4519 ) ;
assign n4521 = sp[2:2] ;
assign n4522 =  ( n4520 ) ^ ( n4521 )  ;
assign n4523 =  ( n4522 ) ^ ( n2282 )  ;
assign n4524 =  ( n4518 ) ? ( n4523 ) : ( n2289 ) ;
assign n4525 =  ( n4515 ) ? ( bv_1_0_n2 ) : ( n4524 ) ;
assign n4526 =  ( n873 ) | ( n882 )  ;
assign n4527 =  ( n4526 ) ? ( bv_1_0_n2 ) : ( n4320 ) ;
assign n4528 =  ( n4514 ) ? ( n4525 ) : ( n4527 ) ;
assign n4529 = ~ ( n4528 ) ;
assign n4530 =  ( n4513 ) | ( n4529 )  ;
assign n4531 = ~ ( n4530 ) ;
assign n4532 =  ( n4478 ) ^ ( n4494 )  ;
assign n4533 = ~ ( n4532 ) ;
assign n4534 =  ( n4511 ) ^ ( n4528 )  ;
assign n4535 = ~ ( n4534 ) ;
assign n4536 =  ( n4533 ) | ( n4535 )  ;
assign n4537 = ~ ( n4536 ) ;
assign n4538 =  ( n4531 ) | ( n4537 )  ;
assign n4539 =  ( n4478 ) ^ ( n4494 )  ;
assign n4540 =  ( n4539 ) ^ ( n4511 )  ;
assign n4541 =  ( n4540 ) ^ ( n4528 )  ;
assign n4542 = ~ ( n4541 ) ;
assign n4543 =  ( n908 ) | ( n917 )  ;
assign n4544 =  ( n532 ) | ( n541 )  ;
assign n4545 = ki[9:9] ;
assign n4546 =  ( n4545 ) == ( bv_1_0_n2 )  ;
assign n4547 =  ( n4546 ) | ( n550 )  ;
assign n4548 = i_wb_data[0:0] ;
assign n4549 = ~ ( n4548 ) ;
assign n4550 =  ( bv_1_1_n5 ) ^ ( n4549 )  ;
assign n4551 = sp[0:0] ;
assign n4552 =  ( n4550 ) ^ ( n4551 )  ;
assign n4553 =  ( n4547 ) ? ( n4552 ) : ( n2910 ) ;
assign n4554 =  ( n4544 ) ? ( bv_1_0_n2 ) : ( n4553 ) ;
assign n4555 =  ( n532 ) | ( n541 )  ;
assign n4556 =  ( n4555 ) ? ( bv_1_0_n2 ) : ( n4349 ) ;
assign n4557 =  ( n4543 ) ? ( n4554 ) : ( n4556 ) ;
assign n4558 = ~ ( n4557 ) ;
assign n4559 =  ( n4542 ) | ( n4558 )  ;
assign n4560 = ~ ( n4559 ) ;
assign n4561 =  ( n4538 ) | ( n4560 )  ;
assign n4562 = ~ ( n4561 ) ;
assign n4563 = ~ ( n4478 ) ;
assign n4564 = ~ ( n4494 ) ;
assign n4565 =  ( n4563 ) | ( n4564 )  ;
assign n4566 = ~ ( n4565 ) ;
assign n4567 = ~ ( n4511 ) ;
assign n4568 = ~ ( n4528 ) ;
assign n4569 =  ( n4567 ) | ( n4568 )  ;
assign n4570 = ~ ( n4569 ) ;
assign n4571 =  ( n4566 ) | ( n4570 )  ;
assign n4572 = ~ ( n4571 ) ;
assign n4573 =  ( n4562 ) | ( n4572 )  ;
assign n4574 =  ( n4274 ) ^ ( n4290 )  ;
assign n4575 =  ( n4574 ) ^ ( n4307 )  ;
assign n4576 =  ( n4575 ) ^ ( n4324 )  ;
assign n4577 =  ( n4576 ) ^ ( n4353 )  ;
assign n4578 = ~ ( n4577 ) ;
assign n4579 =  ( n4573 ) | ( n4578 )  ;
assign n4580 =  ( n567 ) | ( n576 )  ;
assign n4581 = ki[11:11] ;
assign n4582 = ~ ( n4581 ) ;
assign n4583 = ki[10:10] ;
assign n4584 = ~ ( n4583 ) ;
assign n4585 = ki[9:9] ;
assign n4586 = ~ ( n4585 ) ;
assign n4587 =  ( n4584 ) | ( n4586 )  ;
assign n4588 = ~ ( n4587 ) ;
assign n4589 =  ( n4582 ) | ( n4588 )  ;
assign n4590 = ~ ( n4589 ) ;
assign n4591 =  ( n586 ) | ( n595 )  ;
assign n4592 = ki[11:11] ;
assign n4593 =  ( n4592 ) == ( bv_1_0_n2 )  ;
assign n4594 =  ( n4593 ) | ( n604 )  ;
assign n4595 = i_wb_data[0:0] ;
assign n4596 = ~ ( n4595 ) ;
assign n4597 =  ( bv_1_1_n5 ) ^ ( n4596 )  ;
assign n4598 = sp[0:0] ;
assign n4599 =  ( n4597 ) ^ ( n4598 )  ;
assign n4600 =  ( n4594 ) ? ( n4599 ) : ( n2910 ) ;
assign n4601 =  ( n4591 ) ? ( bv_1_0_n2 ) : ( n4600 ) ;
assign n4602 =  ( n4580 ) ? ( n4590 ) : ( n4601 ) ;
assign n4603 = ~ ( n4602 ) ;
assign n4604 =  ( n4579 ) | ( n4603 )  ;
assign n4605 = ~ ( n4604 ) ;
assign n4606 =  ( n4561 ) ^ ( n4571 )  ;
assign n4607 = ~ ( n4606 ) ;
assign n4608 =  ( n4274 ) ^ ( n4290 )  ;
assign n4609 =  ( n4608 ) ^ ( n4307 )  ;
assign n4610 =  ( n4609 ) ^ ( n4324 )  ;
assign n4611 =  ( n4610 ) ^ ( n4353 )  ;
assign n4612 =  ( n4611 ) ^ ( n4602 )  ;
assign n4613 = ~ ( n4612 ) ;
assign n4614 =  ( n4607 ) | ( n4613 )  ;
assign n4615 = ~ ( n4614 ) ;
assign n4616 =  ( n4605 ) | ( n4615 )  ;
assign n4617 =  ( n4561 ) ^ ( n4571 )  ;
assign n4618 =  ( n4617 ) ^ ( n4274 )  ;
assign n4619 =  ( n4618 ) ^ ( n4290 )  ;
assign n4620 =  ( n4619 ) ^ ( n4307 )  ;
assign n4621 =  ( n4620 ) ^ ( n4324 )  ;
assign n4622 =  ( n4621 ) ^ ( n4353 )  ;
assign n4623 =  ( n4622 ) ^ ( n4602 )  ;
assign n4624 = ~ ( n4623 ) ;
assign n4625 = ki[11:11] ;
assign n4626 = ~ ( n4625 ) ;
assign n4627 =  ( n4624 ) | ( n4626 )  ;
assign n4628 =  ( n4627 ) | ( n4588 )  ;
assign n4629 = ~ ( n4628 ) ;
assign n4630 =  ( n4616 ) | ( n4629 )  ;
assign n4631 = ~ ( n4630 ) ;
assign n4632 = ~ ( n4561 ) ;
assign n4633 = ~ ( n4571 ) ;
assign n4634 =  ( n4632 ) | ( n4633 )  ;
assign n4635 = ~ ( n4634 ) ;
assign n4636 =  ( n4274 ) ^ ( n4290 )  ;
assign n4637 =  ( n4636 ) ^ ( n4307 )  ;
assign n4638 =  ( n4637 ) ^ ( n4324 )  ;
assign n4639 =  ( n4638 ) ^ ( n4353 )  ;
assign n4640 = ~ ( n4639 ) ;
assign n4641 = ~ ( n4602 ) ;
assign n4642 =  ( n4640 ) | ( n4641 )  ;
assign n4643 = ~ ( n4642 ) ;
assign n4644 =  ( n4635 ) | ( n4643 )  ;
assign n4645 = ~ ( n4644 ) ;
assign n4646 =  ( n4631 ) | ( n4645 )  ;
assign n4647 = ~ ( n4646 ) ;
assign n4648 =  ( n4605 ) | ( n4615 )  ;
assign n4649 =  ( n4648 ) | ( n4629 )  ;
assign n4650 =  ( n4649 ) ^ ( n4644 )  ;
assign n4651 = ~ ( n4650 ) ;
assign n4652 =  ( n4357 ) ^ ( n4367 )  ;
assign n4653 =  ( n4652 ) ^ ( n4005 )  ;
assign n4654 =  ( n4653 ) ^ ( n4021 )  ;
assign n4655 =  ( n4654 ) ^ ( n4038 )  ;
assign n4656 =  ( n4655 ) ^ ( n4055 )  ;
assign n4657 =  ( n4656 ) ^ ( n4084 )  ;
assign n4658 = ~ ( n4657 ) ;
assign n4659 =  ( n4651 ) | ( n4658 )  ;
assign n4660 = ~ ( n4659 ) ;
assign n4661 =  ( n4647 ) | ( n4660 )  ;
assign n4662 = ~ ( n4661 ) ;
assign n4663 =  ( n4458 ) | ( n4662 )  ;
assign n4664 =  ( n4380 ) ^ ( n4088 )  ;
assign n4665 =  ( n4664 ) ^ ( n4098 )  ;
assign n4666 =  ( n4665 ) ^ ( n3693 )  ;
assign n4667 =  ( n4666 ) ^ ( n3709 )  ;
assign n4668 =  ( n4667 ) ^ ( n3726 )  ;
assign n4669 =  ( n4668 ) ^ ( n3743 )  ;
assign n4670 =  ( n4669 ) ^ ( n3772 )  ;
assign n4671 =  ( n4670 ) ^ ( n3812 )  ;
assign n4672 =  ( n4671 ) ^ ( n3836 )  ;
assign n4673 =  ( n4672 ) ^ ( n3824 )  ;
assign n4674 = ~ ( n4673 ) ;
assign n4675 =  ( n4663 ) | ( n4674 )  ;
assign n4676 =  ( n4390 ) | ( n4403 )  ;
assign n4677 =  ( n4676 ) ^ ( n4111 )  ;
assign n4678 =  ( n4677 ) ^ ( n3776 )  ;
assign n4679 =  ( n4678 ) ^ ( n3786 )  ;
assign n4680 =  ( n4679 ) ^ ( n3847 )  ;
assign n4681 =  ( n4680 ) ^ ( n3413 )  ;
assign n4682 =  ( n4681 ) ^ ( n3429 )  ;
assign n4683 =  ( n4682 ) ^ ( n3446 )  ;
assign n4684 =  ( n4683 ) ^ ( n3463 )  ;
assign n4685 =  ( n4684 ) ^ ( n3492 )  ;
assign n4686 =  ( n4685 ) ^ ( n3881 )  ;
assign n4687 =  ( n4686 ) ^ ( n4139 )  ;
assign n4688 = ~ ( n4687 ) ;
assign n4689 =  ( n4675 ) | ( n4688 )  ;
assign n4690 = ~ ( n4689 ) ;
assign n4691 =  ( n4436 ) | ( n4690 )  ;
assign n4692 = ~ ( n4659 ) ;
assign n4693 =  ( n4647 ) | ( n4692 )  ;
assign n4694 = ~ ( n4693 ) ;
assign n4695 =  ( n4694 ) | ( n4674 )  ;
assign n4696 = ~ ( n4695 ) ;
assign n4697 =  ( n4390 ) | ( n4403 )  ;
assign n4698 =  ( n4696 ) ^ ( n4697 )  ;
assign n4699 =  ( n4698 ) ^ ( n4111 )  ;
assign n4700 =  ( n4699 ) ^ ( n3776 )  ;
assign n4701 =  ( n4700 ) ^ ( n3786 )  ;
assign n4702 =  ( n4701 ) ^ ( n3847 )  ;
assign n4703 =  ( n4702 ) ^ ( n3413 )  ;
assign n4704 =  ( n4703 ) ^ ( n3429 )  ;
assign n4705 =  ( n4704 ) ^ ( n3446 )  ;
assign n4706 =  ( n4705 ) ^ ( n3463 )  ;
assign n4707 =  ( n4706 ) ^ ( n3492 )  ;
assign n4708 =  ( n4707 ) ^ ( n3881 )  ;
assign n4709 =  ( n4708 ) ^ ( n4139 )  ;
assign n4710 = ~ ( n4709 ) ;
assign n4711 =  ( n4458 ) | ( n4710 )  ;
assign n4712 =  ( n4605 ) | ( n4615 )  ;
assign n4713 =  ( n4712 ) | ( n4629 )  ;
assign n4714 =  ( n4713 ) ^ ( n4644 )  ;
assign n4715 =  ( n4714 ) ^ ( n4357 )  ;
assign n4716 =  ( n4715 ) ^ ( n4367 )  ;
assign n4717 =  ( n4716 ) ^ ( n4005 )  ;
assign n4718 =  ( n4717 ) ^ ( n4021 )  ;
assign n4719 =  ( n4718 ) ^ ( n4038 )  ;
assign n4720 =  ( n4719 ) ^ ( n4055 )  ;
assign n4721 =  ( n4720 ) ^ ( n4084 )  ;
assign n4722 = ~ ( n4721 ) ;
assign n4723 =  ( n567 ) | ( n576 )  ;
assign n4724 =  ( n586 ) | ( n595 )  ;
assign n4725 =  ( n4724 ) ? ( bv_1_0_n2 ) : ( n4600 ) ;
assign n4726 =  ( n586 ) | ( n595 )  ;
assign n4727 =  ( n4726 ) ? ( bv_1_0_n2 ) : ( n3799 ) ;
assign n4728 =  ( n4723 ) ? ( n4725 ) : ( n4727 ) ;
assign n4729 = ~ ( n4728 ) ;
assign n4730 =  ( n4722 ) | ( n4729 )  ;
assign n4731 = ~ ( n4659 ) ;
assign n4732 =  ( n4647 ) | ( n4731 )  ;
assign n4733 =  ( n4732 ) ^ ( n4380 )  ;
assign n4734 =  ( n4733 ) ^ ( n4088 )  ;
assign n4735 =  ( n4734 ) ^ ( n4098 )  ;
assign n4736 =  ( n4735 ) ^ ( n3693 )  ;
assign n4737 =  ( n4736 ) ^ ( n3709 )  ;
assign n4738 =  ( n4737 ) ^ ( n3726 )  ;
assign n4739 =  ( n4738 ) ^ ( n3743 )  ;
assign n4740 =  ( n4739 ) ^ ( n3772 )  ;
assign n4741 =  ( n4740 ) ^ ( n3812 )  ;
assign n4742 =  ( n4741 ) ^ ( n3836 )  ;
assign n4743 =  ( n4742 ) ^ ( n3824 )  ;
assign n4744 = ~ ( n4743 ) ;
assign n4745 =  ( n4730 ) | ( n4744 )  ;
assign n4746 = ~ ( n4745 ) ;
assign n4747 = ~ ( n4728 ) ;
assign n4748 =  ( n4722 ) | ( n4747 )  ;
assign n4749 = ~ ( n4748 ) ;
assign n4750 = ~ ( n4659 ) ;
assign n4751 =  ( n4647 ) | ( n4750 )  ;
assign n4752 =  ( n4749 ) ^ ( n4751 )  ;
assign n4753 =  ( n4752 ) ^ ( n4380 )  ;
assign n4754 =  ( n4753 ) ^ ( n4088 )  ;
assign n4755 =  ( n4754 ) ^ ( n4098 )  ;
assign n4756 =  ( n4755 ) ^ ( n3693 )  ;
assign n4757 =  ( n4756 ) ^ ( n3709 )  ;
assign n4758 =  ( n4757 ) ^ ( n3726 )  ;
assign n4759 =  ( n4758 ) ^ ( n3743 )  ;
assign n4760 =  ( n4759 ) ^ ( n3772 )  ;
assign n4761 =  ( n4760 ) ^ ( n3812 )  ;
assign n4762 =  ( n4761 ) ^ ( n3836 )  ;
assign n4763 =  ( n4762 ) ^ ( n3824 )  ;
assign n4764 = ~ ( n4763 ) ;
assign n4765 = ki[0:0] ;
assign n4766 =  ( n4765 ) == ( bv_1_1_n5 )  ;
assign n4767 = ki[1:1] ;
assign n4768 =  ( n4767 ) == ( bv_1_0_n2 )  ;
assign n4769 =  ( n4766 ) | ( n4768 )  ;
assign n4770 = ki[1:1] ;
assign n4771 =  ( n4770 ) == ( bv_1_1_n5 )  ;
assign n4772 = ki[0:0] ;
assign n4773 =  ( n4772 ) == ( bv_1_1_n5 )  ;
assign n4774 =  ( n4771 ) | ( n4773 )  ;
assign n4775 = ki[1:1] ;
assign n4776 =  ( n4775 ) == ( bv_1_1_n5 )  ;
assign n4777 = i_wb_data[7:7] ;
assign n4778 = ~ ( n4777 ) ;
assign n4779 = sp[7:7] ;
assign n4780 =  ( n4778 ) ^ ( n4779 )  ;
assign n4781 =  ( n4780 ) ^ ( n330 )  ;
assign n4782 =  ( n4776 ) ? ( n1035 ) : ( n4781 ) ;
assign n4783 =  ( n4774 ) ? ( n4782 ) : ( bv_1_0_n2 ) ;
assign n4784 =  ( n4769 ) ? ( n4477 ) : ( n4783 ) ;
assign n4785 = ~ ( n4784 ) ;
assign n4786 =  ( n2120 ) | ( n2129 )  ;
assign n4787 =  ( n1838 ) | ( n1847 )  ;
assign n4788 = ki[3:3] ;
assign n4789 =  ( n4788 ) == ( bv_1_0_n2 )  ;
assign n4790 =  ( n4789 ) | ( n1856 )  ;
assign n4791 = i_wb_data[5:5] ;
assign n4792 = ~ ( n4791 ) ;
assign n4793 = sp[5:5] ;
assign n4794 =  ( n4792 ) ^ ( n4793 )  ;
assign n4795 =  ( n4794 ) ^ ( n241 )  ;
assign n4796 =  ( n4790 ) ? ( n4795 ) : ( n2013 ) ;
assign n4797 =  ( n4787 ) ? ( bv_1_0_n2 ) : ( n4796 ) ;
assign n4798 =  ( n1838 ) | ( n1847 )  ;
assign n4799 =  ( n4798 ) ? ( bv_1_0_n2 ) : ( n4490 ) ;
assign n4800 =  ( n4786 ) ? ( n4797 ) : ( n4799 ) ;
assign n4801 = ~ ( n4800 ) ;
assign n4802 =  ( n4785 ) | ( n4801 )  ;
assign n4803 =  ( n1456 ) | ( n1465 )  ;
assign n4804 =  ( n1475 ) | ( n1484 )  ;
assign n4805 = ki[5:5] ;
assign n4806 =  ( n4805 ) == ( bv_1_0_n2 )  ;
assign n4807 =  ( n4806 ) | ( n1493 )  ;
assign n4808 = i_wb_data[3:3] ;
assign n4809 = ~ ( n4808 ) ;
assign n4810 = sp[3:3] ;
assign n4811 =  ( n4809 ) ^ ( n4810 )  ;
assign n4812 =  ( n4811 ) ^ ( n326 )  ;
assign n4813 =  ( n4807 ) ? ( n4812 ) : ( n2306 ) ;
assign n4814 =  ( n4804 ) ? ( bv_1_0_n2 ) : ( n4813 ) ;
assign n4815 =  ( n1475 ) | ( n1484 )  ;
assign n4816 =  ( n4815 ) ? ( bv_1_0_n2 ) : ( n4507 ) ;
assign n4817 =  ( n4803 ) ? ( n4814 ) : ( n4816 ) ;
assign n4818 = ~ ( n4817 ) ;
assign n4819 =  ( n4802 ) | ( n4818 )  ;
assign n4820 =  ( n1257 ) | ( n1266 )  ;
assign n4821 =  ( n873 ) | ( n882 )  ;
assign n4822 = ki[7:7] ;
assign n4823 =  ( n4822 ) == ( bv_1_0_n2 )  ;
assign n4824 =  ( n4823 ) | ( n891 )  ;
assign n4825 = i_wb_data[1:1] ;
assign n4826 = ~ ( n4825 ) ;
assign n4827 = sp[1:1] ;
assign n4828 =  ( n4826 ) ^ ( n4827 )  ;
assign n4829 =  ( n4828 ) ^ ( n237 )  ;
assign n4830 =  ( n4824 ) ? ( n4829 ) : ( n2615 ) ;
assign n4831 =  ( n4821 ) ? ( bv_1_0_n2 ) : ( n4830 ) ;
assign n4832 =  ( n873 ) | ( n882 )  ;
assign n4833 =  ( n4832 ) ? ( bv_1_0_n2 ) : ( n4524 ) ;
assign n4834 =  ( n4820 ) ? ( n4831 ) : ( n4833 ) ;
assign n4835 = ~ ( n4834 ) ;
assign n4836 =  ( n4819 ) | ( n4835 )  ;
assign n4837 = ~ ( n4836 ) ;
assign n4838 =  ( n4784 ) ^ ( n4800 )  ;
assign n4839 = ~ ( n4838 ) ;
assign n4840 =  ( n4817 ) ^ ( n4834 )  ;
assign n4841 = ~ ( n4840 ) ;
assign n4842 =  ( n4839 ) | ( n4841 )  ;
assign n4843 = ~ ( n4842 ) ;
assign n4844 =  ( n4837 ) | ( n4843 )  ;
assign n4845 =  ( n4784 ) ^ ( n4800 )  ;
assign n4846 =  ( n4845 ) ^ ( n4817 )  ;
assign n4847 =  ( n4846 ) ^ ( n4834 )  ;
assign n4848 = ~ ( n4847 ) ;
assign n4849 =  ( n908 ) | ( n917 )  ;
assign n4850 = ki[9:9] ;
assign n4851 = ~ ( n4850 ) ;
assign n4852 = ki[8:8] ;
assign n4853 = ~ ( n4852 ) ;
assign n4854 = ki[7:7] ;
assign n4855 = ~ ( n4854 ) ;
assign n4856 =  ( n4853 ) | ( n4855 )  ;
assign n4857 = ~ ( n4856 ) ;
assign n4858 =  ( n4851 ) | ( n4857 )  ;
assign n4859 = ~ ( n4858 ) ;
assign n4860 =  ( n532 ) | ( n541 )  ;
assign n4861 =  ( n4860 ) ? ( bv_1_0_n2 ) : ( n4553 ) ;
assign n4862 =  ( n4849 ) ? ( n4859 ) : ( n4861 ) ;
assign n4863 = ~ ( n4862 ) ;
assign n4864 =  ( n4848 ) | ( n4863 )  ;
assign n4865 = ~ ( n4864 ) ;
assign n4866 =  ( n4844 ) | ( n4865 )  ;
assign n4867 = ~ ( n4866 ) ;
assign n4868 = ~ ( n4784 ) ;
assign n4869 = ~ ( n4800 ) ;
assign n4870 =  ( n4868 ) | ( n4869 )  ;
assign n4871 = ~ ( n4870 ) ;
assign n4872 = ~ ( n4817 ) ;
assign n4873 = ~ ( n4834 ) ;
assign n4874 =  ( n4872 ) | ( n4873 )  ;
assign n4875 = ~ ( n4874 ) ;
assign n4876 =  ( n4871 ) | ( n4875 )  ;
assign n4877 = ~ ( n4876 ) ;
assign n4878 =  ( n4867 ) | ( n4877 )  ;
assign n4879 = ~ ( n4878 ) ;
assign n4880 =  ( n4866 ) ^ ( n4876 )  ;
assign n4881 = ~ ( n4880 ) ;
assign n4882 =  ( n4478 ) ^ ( n4494 )  ;
assign n4883 =  ( n4882 ) ^ ( n4511 )  ;
assign n4884 =  ( n4883 ) ^ ( n4528 )  ;
assign n4885 =  ( n4884 ) ^ ( n4557 )  ;
assign n4886 = ~ ( n4885 ) ;
assign n4887 =  ( n4881 ) | ( n4886 )  ;
assign n4888 = ~ ( n4887 ) ;
assign n4889 =  ( n4879 ) | ( n4888 )  ;
assign n4890 = ~ ( n4889 ) ;
assign n4891 =  ( n4764 ) | ( n4890 )  ;
assign n4892 =  ( n4561 ) ^ ( n4571 )  ;
assign n4893 =  ( n4892 ) ^ ( n4274 )  ;
assign n4894 =  ( n4893 ) ^ ( n4290 )  ;
assign n4895 =  ( n4894 ) ^ ( n4307 )  ;
assign n4896 =  ( n4895 ) ^ ( n4324 )  ;
assign n4897 =  ( n4896 ) ^ ( n4353 )  ;
assign n4898 =  ( n4897 ) ^ ( n4602 )  ;
assign n4899 =  ( n4898 ) ^ ( n4590 )  ;
assign n4900 = ~ ( n4899 ) ;
assign n4901 =  ( n4891 ) | ( n4900 )  ;
assign n4902 =  ( n4605 ) | ( n4615 )  ;
assign n4903 =  ( n4902 ) | ( n4629 )  ;
assign n4904 =  ( n4903 ) ^ ( n4644 )  ;
assign n4905 =  ( n4904 ) ^ ( n4357 )  ;
assign n4906 =  ( n4905 ) ^ ( n4367 )  ;
assign n4907 =  ( n4906 ) ^ ( n4005 )  ;
assign n4908 =  ( n4907 ) ^ ( n4021 )  ;
assign n4909 =  ( n4908 ) ^ ( n4038 )  ;
assign n4910 =  ( n4909 ) ^ ( n4055 )  ;
assign n4911 =  ( n4910 ) ^ ( n4084 )  ;
assign n4912 =  ( n4911 ) ^ ( n4728 )  ;
assign n4913 = ~ ( n4912 ) ;
assign n4914 =  ( n4901 ) | ( n4913 )  ;
assign n4915 = ~ ( n4914 ) ;
assign n4916 =  ( n4746 ) | ( n4915 )  ;
assign n4917 = ~ ( n4916 ) ;
assign n4918 =  ( n4711 ) | ( n4917 )  ;
assign n4919 = ~ ( n4918 ) ;
assign n4920 =  ( n4691 ) | ( n4919 )  ;
assign n4921 =  ( n4458 ) | ( n4710 )  ;
assign n4922 = ~ ( n4763 ) ;
assign n4923 =  ( n4921 ) | ( n4922 )  ;
assign n4924 = ~ ( n4889 ) ;
assign n4925 =  ( n4924 ) | ( n4900 )  ;
assign n4926 = ~ ( n4925 ) ;
assign n4927 =  ( n4605 ) | ( n4615 )  ;
assign n4928 =  ( n4927 ) | ( n4629 )  ;
assign n4929 =  ( n4926 ) ^ ( n4928 )  ;
assign n4930 =  ( n4929 ) ^ ( n4644 )  ;
assign n4931 =  ( n4930 ) ^ ( n4357 )  ;
assign n4932 =  ( n4931 ) ^ ( n4367 )  ;
assign n4933 =  ( n4932 ) ^ ( n4005 )  ;
assign n4934 =  ( n4933 ) ^ ( n4021 )  ;
assign n4935 =  ( n4934 ) ^ ( n4038 )  ;
assign n4936 =  ( n4935 ) ^ ( n4055 )  ;
assign n4937 =  ( n4936 ) ^ ( n4084 )  ;
assign n4938 =  ( n4937 ) ^ ( n4728 )  ;
assign n4939 = ~ ( n4938 ) ;
assign n4940 =  ( n4923 ) | ( n4939 )  ;
assign n4941 = ki[0:0] ;
assign n4942 =  ( n4941 ) == ( bv_1_1_n5 )  ;
assign n4943 = ki[1:1] ;
assign n4944 =  ( n4943 ) == ( bv_1_0_n2 )  ;
assign n4945 =  ( n4942 ) | ( n4944 )  ;
assign n4946 = ki[1:1] ;
assign n4947 =  ( n4946 ) == ( bv_1_1_n5 )  ;
assign n4948 = ki[0:0] ;
assign n4949 =  ( n4948 ) == ( bv_1_1_n5 )  ;
assign n4950 =  ( n4947 ) | ( n4949 )  ;
assign n4951 = ki[1:1] ;
assign n4952 =  ( n4951 ) == ( bv_1_1_n5 )  ;
assign n4953 = i_wb_data[6:6] ;
assign n4954 = ~ ( n4953 ) ;
assign n4955 = sp[6:6] ;
assign n4956 =  ( n4954 ) ^ ( n4955 )  ;
assign n4957 =  ( n4956 ) ^ ( n1363 )  ;
assign n4958 =  ( n4952 ) ? ( n1370 ) : ( n4957 ) ;
assign n4959 =  ( n4950 ) ? ( n4958 ) : ( bv_1_0_n2 ) ;
assign n4960 =  ( n4945 ) ? ( n4783 ) : ( n4959 ) ;
assign n4961 = ~ ( n4960 ) ;
assign n4962 =  ( n2120 ) | ( n2129 )  ;
assign n4963 =  ( n1838 ) | ( n1847 )  ;
assign n4964 = ki[3:3] ;
assign n4965 =  ( n4964 ) == ( bv_1_0_n2 )  ;
assign n4966 =  ( n4965 ) | ( n1856 )  ;
assign n4967 = i_wb_data[4:4] ;
assign n4968 = ~ ( n4967 ) ;
assign n4969 = sp[4:4] ;
assign n4970 =  ( n4968 ) ^ ( n4969 )  ;
assign n4971 =  ( n4970 ) ^ ( n1989 )  ;
assign n4972 =  ( n4966 ) ? ( n4971 ) : ( n1996 ) ;
assign n4973 =  ( n4963 ) ? ( bv_1_0_n2 ) : ( n4972 ) ;
assign n4974 =  ( n1838 ) | ( n1847 )  ;
assign n4975 =  ( n4974 ) ? ( bv_1_0_n2 ) : ( n4796 ) ;
assign n4976 =  ( n4962 ) ? ( n4973 ) : ( n4975 ) ;
assign n4977 = ~ ( n4976 ) ;
assign n4978 =  ( n4961 ) | ( n4977 )  ;
assign n4979 = ~ ( n4978 ) ;
assign n4980 =  ( n4960 ) ^ ( n4976 )  ;
assign n4981 = ~ ( n4980 ) ;
assign n4982 =  ( n1456 ) | ( n1465 )  ;
assign n4983 =  ( n1475 ) | ( n1484 )  ;
assign n4984 = ki[5:5] ;
assign n4985 =  ( n4984 ) == ( bv_1_0_n2 )  ;
assign n4986 =  ( n4985 ) | ( n1493 )  ;
assign n4987 = i_wb_data[2:2] ;
assign n4988 = ~ ( n4987 ) ;
assign n4989 = sp[2:2] ;
assign n4990 =  ( n4988 ) ^ ( n4989 )  ;
assign n4991 =  ( n4990 ) ^ ( n2282 )  ;
assign n4992 =  ( n4986 ) ? ( n4991 ) : ( n2289 ) ;
assign n4993 =  ( n4983 ) ? ( bv_1_0_n2 ) : ( n4992 ) ;
assign n4994 =  ( n1475 ) | ( n1484 )  ;
assign n4995 =  ( n4994 ) ? ( bv_1_0_n2 ) : ( n4813 ) ;
assign n4996 =  ( n4982 ) ? ( n4993 ) : ( n4995 ) ;
assign n4997 = ~ ( n4996 ) ;
assign n4998 =  ( n4981 ) | ( n4997 )  ;
assign n4999 = ~ ( n4998 ) ;
assign n5000 =  ( n4979 ) | ( n4999 )  ;
assign n5001 = ~ ( n5000 ) ;
assign n5002 =  ( n4784 ) ^ ( n4800 )  ;
assign n5003 =  ( n5002 ) ^ ( n4817 )  ;
assign n5004 =  ( n5003 ) ^ ( n4834 )  ;
assign n5005 =  ( n5004 ) ^ ( n4862 )  ;
assign n5006 = ~ ( n5005 ) ;
assign n5007 =  ( n5001 ) | ( n5006 )  ;
assign n5008 = ~ ( n5007 ) ;
assign n5009 =  ( n5000 ) ^ ( n4784 )  ;
assign n5010 =  ( n5009 ) ^ ( n4800 )  ;
assign n5011 =  ( n5010 ) ^ ( n4817 )  ;
assign n5012 =  ( n5011 ) ^ ( n4834 )  ;
assign n5013 =  ( n5012 ) ^ ( n4862 )  ;
assign n5014 = ~ ( n5013 ) ;
assign n5015 = ki[9:9] ;
assign n5016 = ~ ( n5015 ) ;
assign n5017 =  ( n5014 ) | ( n5016 )  ;
assign n5018 =  ( n5017 ) | ( n4857 )  ;
assign n5019 = ~ ( n5018 ) ;
assign n5020 =  ( n5008 ) | ( n5019 )  ;
assign n5021 = ~ ( n5020 ) ;
assign n5022 =  ( n4866 ) ^ ( n4876 )  ;
assign n5023 =  ( n5022 ) ^ ( n4478 )  ;
assign n5024 =  ( n5023 ) ^ ( n4494 )  ;
assign n5025 =  ( n5024 ) ^ ( n4511 )  ;
assign n5026 =  ( n5025 ) ^ ( n4528 )  ;
assign n5027 =  ( n5026 ) ^ ( n4557 )  ;
assign n5028 = ~ ( n5027 ) ;
assign n5029 =  ( n5021 ) | ( n5028 )  ;
assign n5030 =  ( n4889 ) ^ ( n4561 )  ;
assign n5031 =  ( n5030 ) ^ ( n4571 )  ;
assign n5032 =  ( n5031 ) ^ ( n4274 )  ;
assign n5033 =  ( n5032 ) ^ ( n4290 )  ;
assign n5034 =  ( n5033 ) ^ ( n4307 )  ;
assign n5035 =  ( n5034 ) ^ ( n4324 )  ;
assign n5036 =  ( n5035 ) ^ ( n4353 )  ;
assign n5037 =  ( n5036 ) ^ ( n4602 )  ;
assign n5038 =  ( n5037 ) ^ ( n4590 )  ;
assign n5039 = ~ ( n5038 ) ;
assign n5040 =  ( n5029 ) | ( n5039 )  ;
assign n5041 = ~ ( n5040 ) ;
assign n5042 =  ( n5008 ) | ( n5019 )  ;
assign n5043 = ~ ( n5042 ) ;
assign n5044 =  ( n4866 ) ^ ( n4876 )  ;
assign n5045 =  ( n5044 ) ^ ( n4478 )  ;
assign n5046 =  ( n5045 ) ^ ( n4494 )  ;
assign n5047 =  ( n5046 ) ^ ( n4511 )  ;
assign n5048 =  ( n5047 ) ^ ( n4528 )  ;
assign n5049 =  ( n5048 ) ^ ( n4557 )  ;
assign n5050 = ~ ( n5049 ) ;
assign n5051 =  ( n5043 ) | ( n5050 )  ;
assign n5052 = ~ ( n5051 ) ;
assign n5053 =  ( n5052 ) ^ ( n4889 )  ;
assign n5054 =  ( n5053 ) ^ ( n4561 )  ;
assign n5055 =  ( n5054 ) ^ ( n4571 )  ;
assign n5056 =  ( n5055 ) ^ ( n4274 )  ;
assign n5057 =  ( n5056 ) ^ ( n4290 )  ;
assign n5058 =  ( n5057 ) ^ ( n4307 )  ;
assign n5059 =  ( n5058 ) ^ ( n4324 )  ;
assign n5060 =  ( n5059 ) ^ ( n4353 )  ;
assign n5061 =  ( n5060 ) ^ ( n4602 )  ;
assign n5062 =  ( n5061 ) ^ ( n4590 )  ;
assign n5063 = ~ ( n5062 ) ;
assign n5064 = ki[0:0] ;
assign n5065 =  ( n5064 ) == ( bv_1_1_n5 )  ;
assign n5066 = ki[1:1] ;
assign n5067 =  ( n5066 ) == ( bv_1_0_n2 )  ;
assign n5068 =  ( n5065 ) | ( n5067 )  ;
assign n5069 = ki[1:1] ;
assign n5070 =  ( n5069 ) == ( bv_1_1_n5 )  ;
assign n5071 = ki[0:0] ;
assign n5072 =  ( n5071 ) == ( bv_1_1_n5 )  ;
assign n5073 =  ( n5070 ) | ( n5072 )  ;
assign n5074 = ki[1:1] ;
assign n5075 =  ( n5074 ) == ( bv_1_1_n5 )  ;
assign n5076 = i_wb_data[5:5] ;
assign n5077 = ~ ( n5076 ) ;
assign n5078 = sp[5:5] ;
assign n5079 =  ( n5077 ) ^ ( n5078 )  ;
assign n5080 =  ( n5079 ) ^ ( n241 )  ;
assign n5081 =  ( n5075 ) ? ( n2013 ) : ( n5080 ) ;
assign n5082 =  ( n5073 ) ? ( n5081 ) : ( bv_1_0_n2 ) ;
assign n5083 =  ( n5068 ) ? ( n4959 ) : ( n5082 ) ;
assign n5084 = ~ ( n5083 ) ;
assign n5085 =  ( n2120 ) | ( n2129 )  ;
assign n5086 =  ( n1838 ) | ( n1847 )  ;
assign n5087 = ki[3:3] ;
assign n5088 =  ( n5087 ) == ( bv_1_0_n2 )  ;
assign n5089 =  ( n5088 ) | ( n1856 )  ;
assign n5090 = i_wb_data[3:3] ;
assign n5091 = ~ ( n5090 ) ;
assign n5092 = sp[3:3] ;
assign n5093 =  ( n5091 ) ^ ( n5092 )  ;
assign n5094 =  ( n5093 ) ^ ( n326 )  ;
assign n5095 =  ( n5089 ) ? ( n5094 ) : ( n2306 ) ;
assign n5096 =  ( n5086 ) ? ( bv_1_0_n2 ) : ( n5095 ) ;
assign n5097 =  ( n1838 ) | ( n1847 )  ;
assign n5098 =  ( n5097 ) ? ( bv_1_0_n2 ) : ( n4972 ) ;
assign n5099 =  ( n5085 ) ? ( n5096 ) : ( n5098 ) ;
assign n5100 = ~ ( n5099 ) ;
assign n5101 =  ( n5084 ) | ( n5100 )  ;
assign n5102 =  ( n1456 ) | ( n1465 )  ;
assign n5103 =  ( n1475 ) | ( n1484 )  ;
assign n5104 = ki[5:5] ;
assign n5105 =  ( n5104 ) == ( bv_1_0_n2 )  ;
assign n5106 =  ( n5105 ) | ( n1493 )  ;
assign n5107 = i_wb_data[1:1] ;
assign n5108 = ~ ( n5107 ) ;
assign n5109 = sp[1:1] ;
assign n5110 =  ( n5108 ) ^ ( n5109 )  ;
assign n5111 =  ( n5110 ) ^ ( n237 )  ;
assign n5112 =  ( n5106 ) ? ( n5111 ) : ( n2615 ) ;
assign n5113 =  ( n5103 ) ? ( bv_1_0_n2 ) : ( n5112 ) ;
assign n5114 =  ( n1475 ) | ( n1484 )  ;
assign n5115 =  ( n5114 ) ? ( bv_1_0_n2 ) : ( n4992 ) ;
assign n5116 =  ( n5102 ) ? ( n5113 ) : ( n5115 ) ;
assign n5117 = ~ ( n5116 ) ;
assign n5118 =  ( n5101 ) | ( n5117 )  ;
assign n5119 =  ( n1257 ) | ( n1266 )  ;
assign n5120 = ki[7:7] ;
assign n5121 = ~ ( n5120 ) ;
assign n5122 = ki[6:6] ;
assign n5123 = ~ ( n5122 ) ;
assign n5124 = ki[5:5] ;
assign n5125 = ~ ( n5124 ) ;
assign n5126 =  ( n5123 ) | ( n5125 )  ;
assign n5127 = ~ ( n5126 ) ;
assign n5128 =  ( n5121 ) | ( n5127 )  ;
assign n5129 = ~ ( n5128 ) ;
assign n5130 =  ( n873 ) | ( n882 )  ;
assign n5131 = ki[7:7] ;
assign n5132 =  ( n5131 ) == ( bv_1_0_n2 )  ;
assign n5133 =  ( n5132 ) | ( n891 )  ;
assign n5134 = i_wb_data[0:0] ;
assign n5135 = ~ ( n5134 ) ;
assign n5136 =  ( bv_1_1_n5 ) ^ ( n5135 )  ;
assign n5137 = sp[0:0] ;
assign n5138 =  ( n5136 ) ^ ( n5137 )  ;
assign n5139 =  ( n5133 ) ? ( n5138 ) : ( n2910 ) ;
assign n5140 =  ( n5130 ) ? ( bv_1_0_n2 ) : ( n5139 ) ;
assign n5141 =  ( n5119 ) ? ( n5129 ) : ( n5140 ) ;
assign n5142 = ~ ( n5141 ) ;
assign n5143 =  ( n5118 ) | ( n5142 )  ;
assign n5144 = ~ ( n5143 ) ;
assign n5145 =  ( n5083 ) ^ ( n5099 )  ;
assign n5146 = ~ ( n5145 ) ;
assign n5147 =  ( n5116 ) ^ ( n5141 )  ;
assign n5148 = ~ ( n5147 ) ;
assign n5149 =  ( n5146 ) | ( n5148 )  ;
assign n5150 = ~ ( n5149 ) ;
assign n5151 =  ( n5144 ) | ( n5150 )  ;
assign n5152 =  ( n5083 ) ^ ( n5099 )  ;
assign n5153 =  ( n5152 ) ^ ( n5116 )  ;
assign n5154 =  ( n5153 ) ^ ( n5141 )  ;
assign n5155 = ~ ( n5154 ) ;
assign n5156 = ki[7:7] ;
assign n5157 = ~ ( n5156 ) ;
assign n5158 =  ( n5155 ) | ( n5157 )  ;
assign n5159 =  ( n5158 ) | ( n5127 )  ;
assign n5160 = ~ ( n5159 ) ;
assign n5161 =  ( n5151 ) | ( n5160 )  ;
assign n5162 = ~ ( n5161 ) ;
assign n5163 = ~ ( n5083 ) ;
assign n5164 = ~ ( n5099 ) ;
assign n5165 =  ( n5163 ) | ( n5164 )  ;
assign n5166 = ~ ( n5165 ) ;
assign n5167 = ~ ( n5116 ) ;
assign n5168 = ~ ( n5141 ) ;
assign n5169 =  ( n5167 ) | ( n5168 )  ;
assign n5170 = ~ ( n5169 ) ;
assign n5171 =  ( n5166 ) | ( n5170 )  ;
assign n5172 = ~ ( n5171 ) ;
assign n5173 =  ( n5162 ) | ( n5172 )  ;
assign n5174 = ~ ( n5173 ) ;
assign n5175 =  ( n5161 ) ^ ( n5171 )  ;
assign n5176 = ~ ( n5175 ) ;
assign n5177 =  ( n4960 ) ^ ( n4976 )  ;
assign n5178 =  ( n5177 ) ^ ( n4996 )  ;
assign n5179 = ~ ( n5178 ) ;
assign n5180 =  ( n5176 ) | ( n5179 )  ;
assign n5181 = ~ ( n5180 ) ;
assign n5182 =  ( n5174 ) | ( n5181 )  ;
assign n5183 = ~ ( n5182 ) ;
assign n5184 =  ( n5063 ) | ( n5183 )  ;
assign n5185 =  ( n5000 ) ^ ( n4784 )  ;
assign n5186 =  ( n5185 ) ^ ( n4800 )  ;
assign n5187 =  ( n5186 ) ^ ( n4817 )  ;
assign n5188 =  ( n5187 ) ^ ( n4834 )  ;
assign n5189 =  ( n5188 ) ^ ( n4862 )  ;
assign n5190 =  ( n5189 ) ^ ( n4859 )  ;
assign n5191 = ~ ( n5190 ) ;
assign n5192 =  ( n5184 ) | ( n5191 )  ;
assign n5193 =  ( n5008 ) | ( n5019 )  ;
assign n5194 =  ( n5193 ) ^ ( n4866 )  ;
assign n5195 =  ( n5194 ) ^ ( n4876 )  ;
assign n5196 =  ( n5195 ) ^ ( n4478 )  ;
assign n5197 =  ( n5196 ) ^ ( n4494 )  ;
assign n5198 =  ( n5197 ) ^ ( n4511 )  ;
assign n5199 =  ( n5198 ) ^ ( n4528 )  ;
assign n5200 =  ( n5199 ) ^ ( n4557 )  ;
assign n5201 = ~ ( n5200 ) ;
assign n5202 =  ( n5192 ) | ( n5201 )  ;
assign n5203 = ~ ( n5202 ) ;
assign n5204 =  ( n5041 ) | ( n5203 )  ;
assign n5205 = ~ ( n5182 ) ;
assign n5206 =  ( n5000 ) ^ ( n4784 )  ;
assign n5207 =  ( n5206 ) ^ ( n4800 )  ;
assign n5208 =  ( n5207 ) ^ ( n4817 )  ;
assign n5209 =  ( n5208 ) ^ ( n4834 )  ;
assign n5210 =  ( n5209 ) ^ ( n4862 )  ;
assign n5211 =  ( n5210 ) ^ ( n4859 )  ;
assign n5212 = ~ ( n5211 ) ;
assign n5213 =  ( n5205 ) | ( n5212 )  ;
assign n5214 = ~ ( n5213 ) ;
assign n5215 =  ( n5008 ) | ( n5019 )  ;
assign n5216 =  ( n5214 ) ^ ( n5215 )  ;
assign n5217 =  ( n5216 ) ^ ( n4866 )  ;
assign n5218 =  ( n5217 ) ^ ( n4876 )  ;
assign n5219 =  ( n5218 ) ^ ( n4478 )  ;
assign n5220 =  ( n5219 ) ^ ( n4494 )  ;
assign n5221 =  ( n5220 ) ^ ( n4511 )  ;
assign n5222 =  ( n5221 ) ^ ( n4528 )  ;
assign n5223 =  ( n5222 ) ^ ( n4557 )  ;
assign n5224 = ~ ( n5223 ) ;
assign n5225 =  ( n5063 ) | ( n5224 )  ;
assign n5226 =  ( n5161 ) ^ ( n5171 )  ;
assign n5227 =  ( n5226 ) ^ ( n4960 )  ;
assign n5228 =  ( n5227 ) ^ ( n4976 )  ;
assign n5229 =  ( n5228 ) ^ ( n4996 )  ;
assign n5230 = ~ ( n5229 ) ;
assign n5231 =  ( n1257 ) | ( n1266 )  ;
assign n5232 =  ( n873 ) | ( n882 )  ;
assign n5233 =  ( n5232 ) ? ( bv_1_0_n2 ) : ( n5139 ) ;
assign n5234 =  ( n873 ) | ( n882 )  ;
assign n5235 =  ( n5234 ) ? ( bv_1_0_n2 ) : ( n4830 ) ;
assign n5236 =  ( n5231 ) ? ( n5233 ) : ( n5235 ) ;
assign n5237 = ~ ( n5236 ) ;
assign n5238 =  ( n5230 ) | ( n5237 )  ;
assign n5239 =  ( n5182 ) ^ ( n5000 )  ;
assign n5240 =  ( n5239 ) ^ ( n4784 )  ;
assign n5241 =  ( n5240 ) ^ ( n4800 )  ;
assign n5242 =  ( n5241 ) ^ ( n4817 )  ;
assign n5243 =  ( n5242 ) ^ ( n4834 )  ;
assign n5244 =  ( n5243 ) ^ ( n4862 )  ;
assign n5245 =  ( n5244 ) ^ ( n4859 )  ;
assign n5246 = ~ ( n5245 ) ;
assign n5247 =  ( n5238 ) | ( n5246 )  ;
assign n5248 = ~ ( n5247 ) ;
assign n5249 =  ( n5161 ) ^ ( n5171 )  ;
assign n5250 =  ( n5249 ) ^ ( n4960 )  ;
assign n5251 =  ( n5250 ) ^ ( n4976 )  ;
assign n5252 =  ( n5251 ) ^ ( n4996 )  ;
assign n5253 = ~ ( n5252 ) ;
assign n5254 = ~ ( n5236 ) ;
assign n5255 =  ( n5253 ) | ( n5254 )  ;
assign n5256 = ~ ( n5255 ) ;
assign n5257 =  ( n5256 ) ^ ( n5182 )  ;
assign n5258 =  ( n5257 ) ^ ( n5000 )  ;
assign n5259 =  ( n5258 ) ^ ( n4784 )  ;
assign n5260 =  ( n5259 ) ^ ( n4800 )  ;
assign n5261 =  ( n5260 ) ^ ( n4817 )  ;
assign n5262 =  ( n5261 ) ^ ( n4834 )  ;
assign n5263 =  ( n5262 ) ^ ( n4862 )  ;
assign n5264 =  ( n5263 ) ^ ( n4859 )  ;
assign n5265 = ~ ( n5264 ) ;
assign n5266 = ki[0:0] ;
assign n5267 =  ( n5266 ) == ( bv_1_1_n5 )  ;
assign n5268 = ki[1:1] ;
assign n5269 =  ( n5268 ) == ( bv_1_0_n2 )  ;
assign n5270 =  ( n5267 ) | ( n5269 )  ;
assign n5271 = ki[1:1] ;
assign n5272 =  ( n5271 ) == ( bv_1_1_n5 )  ;
assign n5273 = ki[0:0] ;
assign n5274 =  ( n5273 ) == ( bv_1_1_n5 )  ;
assign n5275 =  ( n5272 ) | ( n5274 )  ;
assign n5276 = ki[1:1] ;
assign n5277 =  ( n5276 ) == ( bv_1_1_n5 )  ;
assign n5278 = i_wb_data[4:4] ;
assign n5279 = ~ ( n5278 ) ;
assign n5280 = sp[4:4] ;
assign n5281 =  ( n5279 ) ^ ( n5280 )  ;
assign n5282 =  ( n5281 ) ^ ( n1989 )  ;
assign n5283 =  ( n5277 ) ? ( n1996 ) : ( n5282 ) ;
assign n5284 =  ( n5275 ) ? ( n5283 ) : ( bv_1_0_n2 ) ;
assign n5285 =  ( n5270 ) ? ( n5082 ) : ( n5284 ) ;
assign n5286 = ~ ( n5285 ) ;
assign n5287 =  ( n2120 ) | ( n2129 )  ;
assign n5288 =  ( n1838 ) | ( n1847 )  ;
assign n5289 = ki[3:3] ;
assign n5290 =  ( n5289 ) == ( bv_1_0_n2 )  ;
assign n5291 =  ( n5290 ) | ( n1856 )  ;
assign n5292 = i_wb_data[2:2] ;
assign n5293 = ~ ( n5292 ) ;
assign n5294 = sp[2:2] ;
assign n5295 =  ( n5293 ) ^ ( n5294 )  ;
assign n5296 =  ( n5295 ) ^ ( n2282 )  ;
assign n5297 =  ( n5291 ) ? ( n5296 ) : ( n2289 ) ;
assign n5298 =  ( n5288 ) ? ( bv_1_0_n2 ) : ( n5297 ) ;
assign n5299 =  ( n1838 ) | ( n1847 )  ;
assign n5300 =  ( n5299 ) ? ( bv_1_0_n2 ) : ( n5095 ) ;
assign n5301 =  ( n5287 ) ? ( n5298 ) : ( n5300 ) ;
assign n5302 = ~ ( n5301 ) ;
assign n5303 =  ( n5286 ) | ( n5302 )  ;
assign n5304 = ~ ( n5303 ) ;
assign n5305 =  ( n5285 ) ^ ( n5301 )  ;
assign n5306 = ~ ( n5305 ) ;
assign n5307 =  ( n1456 ) | ( n1465 )  ;
assign n5308 =  ( n1475 ) | ( n1484 )  ;
assign n5309 = ki[5:5] ;
assign n5310 =  ( n5309 ) == ( bv_1_0_n2 )  ;
assign n5311 =  ( n5310 ) | ( n1493 )  ;
assign n5312 = i_wb_data[0:0] ;
assign n5313 = ~ ( n5312 ) ;
assign n5314 =  ( bv_1_1_n5 ) ^ ( n5313 )  ;
assign n5315 = sp[0:0] ;
assign n5316 =  ( n5314 ) ^ ( n5315 )  ;
assign n5317 =  ( n5311 ) ? ( n5316 ) : ( n2910 ) ;
assign n5318 =  ( n5308 ) ? ( bv_1_0_n2 ) : ( n5317 ) ;
assign n5319 =  ( n1475 ) | ( n1484 )  ;
assign n5320 =  ( n5319 ) ? ( bv_1_0_n2 ) : ( n5112 ) ;
assign n5321 =  ( n5307 ) ? ( n5318 ) : ( n5320 ) ;
assign n5322 = ~ ( n5321 ) ;
assign n5323 =  ( n5306 ) | ( n5322 )  ;
assign n5324 = ~ ( n5323 ) ;
assign n5325 =  ( n5304 ) | ( n5324 )  ;
assign n5326 = ~ ( n5325 ) ;
assign n5327 =  ( n5265 ) | ( n5326 )  ;
assign n5328 =  ( n5083 ) ^ ( n5099 )  ;
assign n5329 =  ( n5328 ) ^ ( n5116 )  ;
assign n5330 =  ( n5329 ) ^ ( n5141 )  ;
assign n5331 =  ( n5330 ) ^ ( n5129 )  ;
assign n5332 = ~ ( n5331 ) ;
assign n5333 =  ( n5327 ) | ( n5332 )  ;
assign n5334 =  ( n5161 ) ^ ( n5171 )  ;
assign n5335 =  ( n5334 ) ^ ( n4960 )  ;
assign n5336 =  ( n5335 ) ^ ( n4976 )  ;
assign n5337 =  ( n5336 ) ^ ( n4996 )  ;
assign n5338 =  ( n5337 ) ^ ( n5236 )  ;
assign n5339 = ~ ( n5338 ) ;
assign n5340 =  ( n5333 ) | ( n5339 )  ;
assign n5341 = ~ ( n5340 ) ;
assign n5342 =  ( n5248 ) | ( n5341 )  ;
assign n5343 = ~ ( n5342 ) ;
assign n5344 =  ( n5225 ) | ( n5343 )  ;
assign n5345 = ~ ( n5344 ) ;
assign n5346 =  ( n5204 ) | ( n5345 )  ;
assign n5347 = ~ ( n5346 ) ;
assign n5348 =  ( n4940 ) | ( n5347 )  ;
assign n5349 = ~ ( n5348 ) ;
assign n5350 =  ( n4920 ) | ( n5349 )  ;
assign n5351 =  ( n4458 ) | ( n4710 )  ;
assign n5352 = ~ ( n4763 ) ;
assign n5353 =  ( n5351 ) | ( n5352 )  ;
assign n5354 = ~ ( n4938 ) ;
assign n5355 =  ( n5353 ) | ( n5354 )  ;
assign n5356 =  ( n5355 ) | ( n5063 )  ;
assign n5357 =  ( n5356 ) | ( n5224 )  ;
assign n5358 =  ( n5357 ) | ( n5265 )  ;
assign n5359 = ~ ( n5325 ) ;
assign n5360 =  ( n5083 ) ^ ( n5099 )  ;
assign n5361 =  ( n5360 ) ^ ( n5116 )  ;
assign n5362 =  ( n5361 ) ^ ( n5141 )  ;
assign n5363 =  ( n5362 ) ^ ( n5129 )  ;
assign n5364 = ~ ( n5363 ) ;
assign n5365 =  ( n5359 ) | ( n5364 )  ;
assign n5366 = ~ ( n5365 ) ;
assign n5367 =  ( n5366 ) ^ ( n5161 )  ;
assign n5368 =  ( n5367 ) ^ ( n5171 )  ;
assign n5369 =  ( n5368 ) ^ ( n4960 )  ;
assign n5370 =  ( n5369 ) ^ ( n4976 )  ;
assign n5371 =  ( n5370 ) ^ ( n4996 )  ;
assign n5372 =  ( n5371 ) ^ ( n5236 )  ;
assign n5373 = ~ ( n5372 ) ;
assign n5374 =  ( n5358 ) | ( n5373 )  ;
assign n5375 = ki[0:0] ;
assign n5376 =  ( n5375 ) == ( bv_1_1_n5 )  ;
assign n5377 = ki[1:1] ;
assign n5378 =  ( n5377 ) == ( bv_1_0_n2 )  ;
assign n5379 =  ( n5376 ) | ( n5378 )  ;
assign n5380 = ki[1:1] ;
assign n5381 =  ( n5380 ) == ( bv_1_1_n5 )  ;
assign n5382 = ki[0:0] ;
assign n5383 =  ( n5382 ) == ( bv_1_1_n5 )  ;
assign n5384 =  ( n5381 ) | ( n5383 )  ;
assign n5385 = ki[1:1] ;
assign n5386 =  ( n5385 ) == ( bv_1_1_n5 )  ;
assign n5387 = i_wb_data[3:3] ;
assign n5388 = ~ ( n5387 ) ;
assign n5389 = sp[3:3] ;
assign n5390 =  ( n5388 ) ^ ( n5389 )  ;
assign n5391 =  ( n5390 ) ^ ( n326 )  ;
assign n5392 =  ( n5386 ) ? ( n2306 ) : ( n5391 ) ;
assign n5393 =  ( n5384 ) ? ( n5392 ) : ( bv_1_0_n2 ) ;
assign n5394 =  ( n5379 ) ? ( n5284 ) : ( n5393 ) ;
assign n5395 = ~ ( n5394 ) ;
assign n5396 =  ( n2120 ) | ( n2129 )  ;
assign n5397 =  ( n1838 ) | ( n1847 )  ;
assign n5398 = ki[3:3] ;
assign n5399 =  ( n5398 ) == ( bv_1_0_n2 )  ;
assign n5400 =  ( n5399 ) | ( n1856 )  ;
assign n5401 = i_wb_data[1:1] ;
assign n5402 = ~ ( n5401 ) ;
assign n5403 = sp[1:1] ;
assign n5404 =  ( n5402 ) ^ ( n5403 )  ;
assign n5405 =  ( n5404 ) ^ ( n237 )  ;
assign n5406 =  ( n5400 ) ? ( n5405 ) : ( n2615 ) ;
assign n5407 =  ( n5397 ) ? ( bv_1_0_n2 ) : ( n5406 ) ;
assign n5408 =  ( n1838 ) | ( n1847 )  ;
assign n5409 =  ( n5408 ) ? ( bv_1_0_n2 ) : ( n5297 ) ;
assign n5410 =  ( n5396 ) ? ( n5407 ) : ( n5409 ) ;
assign n5411 = ~ ( n5410 ) ;
assign n5412 =  ( n5395 ) | ( n5411 )  ;
assign n5413 = ~ ( n5412 ) ;
assign n5414 =  ( n5394 ) ^ ( n5410 )  ;
assign n5415 = ~ ( n5414 ) ;
assign n5416 =  ( n1456 ) | ( n1465 )  ;
assign n5417 = ki[5:5] ;
assign n5418 = ~ ( n5417 ) ;
assign n5419 = ki[4:4] ;
assign n5420 = ~ ( n5419 ) ;
assign n5421 = ki[3:3] ;
assign n5422 = ~ ( n5421 ) ;
assign n5423 =  ( n5420 ) | ( n5422 )  ;
assign n5424 = ~ ( n5423 ) ;
assign n5425 =  ( n5418 ) | ( n5424 )  ;
assign n5426 = ~ ( n5425 ) ;
assign n5427 =  ( n1475 ) | ( n1484 )  ;
assign n5428 =  ( n5427 ) ? ( bv_1_0_n2 ) : ( n5317 ) ;
assign n5429 =  ( n5416 ) ? ( n5426 ) : ( n5428 ) ;
assign n5430 = ~ ( n5429 ) ;
assign n5431 =  ( n5415 ) | ( n5430 )  ;
assign n5432 = ~ ( n5431 ) ;
assign n5433 =  ( n5413 ) | ( n5432 )  ;
assign n5434 = ~ ( n5433 ) ;
assign n5435 =  ( n5285 ) ^ ( n5301 )  ;
assign n5436 =  ( n5435 ) ^ ( n5321 )  ;
assign n5437 = ~ ( n5436 ) ;
assign n5438 =  ( n5434 ) | ( n5437 )  ;
assign n5439 =  ( n5325 ) ^ ( n5083 )  ;
assign n5440 =  ( n5439 ) ^ ( n5099 )  ;
assign n5441 =  ( n5440 ) ^ ( n5116 )  ;
assign n5442 =  ( n5441 ) ^ ( n5141 )  ;
assign n5443 =  ( n5442 ) ^ ( n5129 )  ;
assign n5444 = ~ ( n5443 ) ;
assign n5445 =  ( n5438 ) | ( n5444 )  ;
assign n5446 = ~ ( n5445 ) ;
assign n5447 = ~ ( n5433 ) ;
assign n5448 =  ( n5285 ) ^ ( n5301 )  ;
assign n5449 =  ( n5448 ) ^ ( n5321 )  ;
assign n5450 = ~ ( n5449 ) ;
assign n5451 =  ( n5447 ) | ( n5450 )  ;
assign n5452 = ~ ( n5451 ) ;
assign n5453 =  ( n5452 ) ^ ( n5325 )  ;
assign n5454 =  ( n5453 ) ^ ( n5083 )  ;
assign n5455 =  ( n5454 ) ^ ( n5099 )  ;
assign n5456 =  ( n5455 ) ^ ( n5116 )  ;
assign n5457 =  ( n5456 ) ^ ( n5141 )  ;
assign n5458 =  ( n5457 ) ^ ( n5129 )  ;
assign n5459 = ~ ( n5458 ) ;
assign n5460 =  ( n5394 ) ^ ( n5410 )  ;
assign n5461 =  ( n5460 ) ^ ( n5429 )  ;
assign n5462 = ~ ( n5461 ) ;
assign n5463 =  ( n5459 ) | ( n5462 )  ;
assign n5464 = ki[5:5] ;
assign n5465 = ~ ( n5464 ) ;
assign n5466 =  ( n5463 ) | ( n5465 )  ;
assign n5467 =  ( n5466 ) | ( n5424 )  ;
assign n5468 =  ( n5433 ) ^ ( n5285 )  ;
assign n5469 =  ( n5468 ) ^ ( n5301 )  ;
assign n5470 =  ( n5469 ) ^ ( n5321 )  ;
assign n5471 = ~ ( n5470 ) ;
assign n5472 =  ( n5467 ) | ( n5471 )  ;
assign n5473 = ~ ( n5472 ) ;
assign n5474 =  ( n5446 ) | ( n5473 )  ;
assign n5475 =  ( n5452 ) ^ ( n5325 )  ;
assign n5476 =  ( n5475 ) ^ ( n5083 )  ;
assign n5477 =  ( n5476 ) ^ ( n5099 )  ;
assign n5478 =  ( n5477 ) ^ ( n5116 )  ;
assign n5479 =  ( n5478 ) ^ ( n5141 )  ;
assign n5480 =  ( n5479 ) ^ ( n5129 )  ;
assign n5481 = ~ ( n5480 ) ;
assign n5482 =  ( n5394 ) ^ ( n5410 )  ;
assign n5483 =  ( n5482 ) ^ ( n5429 )  ;
assign n5484 = ~ ( n5483 ) ;
assign n5485 = ki[5:5] ;
assign n5486 = ~ ( n5485 ) ;
assign n5487 =  ( n5484 ) | ( n5486 )  ;
assign n5488 =  ( n5487 ) | ( n5424 )  ;
assign n5489 = ~ ( n5488 ) ;
assign n5490 =  ( n5489 ) ^ ( n5433 )  ;
assign n5491 =  ( n5490 ) ^ ( n5285 )  ;
assign n5492 =  ( n5491 ) ^ ( n5301 )  ;
assign n5493 =  ( n5492 ) ^ ( n5321 )  ;
assign n5494 = ~ ( n5493 ) ;
assign n5495 =  ( n5481 ) | ( n5494 )  ;
assign n5496 = ki[0:0] ;
assign n5497 =  ( n5496 ) == ( bv_1_1_n5 )  ;
assign n5498 = ki[1:1] ;
assign n5499 =  ( n5498 ) == ( bv_1_0_n2 )  ;
assign n5500 =  ( n5497 ) | ( n5499 )  ;
assign n5501 = ki[1:1] ;
assign n5502 =  ( n5501 ) == ( bv_1_1_n5 )  ;
assign n5503 = ki[0:0] ;
assign n5504 =  ( n5503 ) == ( bv_1_1_n5 )  ;
assign n5505 =  ( n5502 ) | ( n5504 )  ;
assign n5506 = ki[1:1] ;
assign n5507 =  ( n5506 ) == ( bv_1_1_n5 )  ;
assign n5508 = i_wb_data[2:2] ;
assign n5509 = ~ ( n5508 ) ;
assign n5510 = sp[2:2] ;
assign n5511 =  ( n5509 ) ^ ( n5510 )  ;
assign n5512 =  ( n5511 ) ^ ( n2282 )  ;
assign n5513 =  ( n5507 ) ? ( n2289 ) : ( n5512 ) ;
assign n5514 =  ( n5505 ) ? ( n5513 ) : ( bv_1_0_n2 ) ;
assign n5515 =  ( n5500 ) ? ( n5393 ) : ( n5514 ) ;
assign n5516 = ~ ( n5515 ) ;
assign n5517 =  ( n2120 ) | ( n2129 )  ;
assign n5518 =  ( n1838 ) | ( n1847 )  ;
assign n5519 = ki[3:3] ;
assign n5520 =  ( n5519 ) == ( bv_1_0_n2 )  ;
assign n5521 =  ( n5520 ) | ( n1856 )  ;
assign n5522 = i_wb_data[0:0] ;
assign n5523 = ~ ( n5522 ) ;
assign n5524 =  ( bv_1_1_n5 ) ^ ( n5523 )  ;
assign n5525 = sp[0:0] ;
assign n5526 =  ( n5524 ) ^ ( n5525 )  ;
assign n5527 =  ( n5521 ) ? ( n5526 ) : ( n2910 ) ;
assign n5528 =  ( n5518 ) ? ( bv_1_0_n2 ) : ( n5527 ) ;
assign n5529 =  ( n1838 ) | ( n1847 )  ;
assign n5530 =  ( n5529 ) ? ( bv_1_0_n2 ) : ( n5406 ) ;
assign n5531 =  ( n5517 ) ? ( n5528 ) : ( n5530 ) ;
assign n5532 = ~ ( n5531 ) ;
assign n5533 =  ( n5516 ) | ( n5532 )  ;
assign n5534 =  ( n5394 ) ^ ( n5410 )  ;
assign n5535 =  ( n5534 ) ^ ( n5429 )  ;
assign n5536 =  ( n5535 ) ^ ( n5426 )  ;
assign n5537 = ~ ( n5536 ) ;
assign n5538 =  ( n5533 ) | ( n5537 )  ;
assign n5539 = ~ ( n5538 ) ;
assign n5540 = ~ ( n5515 ) ;
assign n5541 = ~ ( n5531 ) ;
assign n5542 =  ( n5540 ) | ( n5541 )  ;
assign n5543 = ~ ( n5542 ) ;
assign n5544 =  ( n5543 ) ^ ( n5394 )  ;
assign n5545 =  ( n5544 ) ^ ( n5410 )  ;
assign n5546 =  ( n5545 ) ^ ( n5429 )  ;
assign n5547 =  ( n5546 ) ^ ( n5426 )  ;
assign n5548 = ~ ( n5547 ) ;
assign n5549 = ki[0:0] ;
assign n5550 =  ( n5549 ) == ( bv_1_1_n5 )  ;
assign n5551 = ki[1:1] ;
assign n5552 =  ( n5551 ) == ( bv_1_0_n2 )  ;
assign n5553 =  ( n5550 ) | ( n5552 )  ;
assign n5554 = ki[1:1] ;
assign n5555 =  ( n5554 ) == ( bv_1_1_n5 )  ;
assign n5556 = ki[0:0] ;
assign n5557 =  ( n5556 ) == ( bv_1_1_n5 )  ;
assign n5558 =  ( n5555 ) | ( n5557 )  ;
assign n5559 = ki[1:1] ;
assign n5560 =  ( n5559 ) == ( bv_1_1_n5 )  ;
assign n5561 = i_wb_data[1:1] ;
assign n5562 = ~ ( n5561 ) ;
assign n5563 = sp[1:1] ;
assign n5564 =  ( n5562 ) ^ ( n5563 )  ;
assign n5565 =  ( n5564 ) ^ ( n237 )  ;
assign n5566 =  ( n5560 ) ? ( n2615 ) : ( n5565 ) ;
assign n5567 =  ( n5558 ) ? ( n5566 ) : ( bv_1_0_n2 ) ;
assign n5568 =  ( n5553 ) ? ( n5514 ) : ( n5567 ) ;
assign n5569 = ~ ( n5568 ) ;
assign n5570 =  ( n2120 ) | ( n2129 )  ;
assign n5571 = ki[3:3] ;
assign n5572 = ~ ( n5571 ) ;
assign n5573 = ki[2:2] ;
assign n5574 = ~ ( n5573 ) ;
assign n5575 = ki[1:1] ;
assign n5576 = ~ ( n5575 ) ;
assign n5577 =  ( n5574 ) | ( n5576 )  ;
assign n5578 = ~ ( n5577 ) ;
assign n5579 =  ( n5572 ) | ( n5578 )  ;
assign n5580 = ~ ( n5579 ) ;
assign n5581 =  ( n1838 ) | ( n1847 )  ;
assign n5582 =  ( n5581 ) ? ( bv_1_0_n2 ) : ( n5527 ) ;
assign n5583 =  ( n5570 ) ? ( n5580 ) : ( n5582 ) ;
assign n5584 = ~ ( n5583 ) ;
assign n5585 =  ( n5569 ) | ( n5584 )  ;
assign n5586 = ~ ( n5585 ) ;
assign n5587 =  ( n5568 ) ^ ( n5583 )  ;
assign n5588 = ~ ( n5587 ) ;
assign n5589 = ki[3:3] ;
assign n5590 = ~ ( n5589 ) ;
assign n5591 =  ( n5588 ) | ( n5590 )  ;
assign n5592 =  ( n5591 ) | ( n5578 )  ;
assign n5593 = ~ ( n5592 ) ;
assign n5594 =  ( n5586 ) | ( n5593 )  ;
assign n5595 = ~ ( n5594 ) ;
assign n5596 =  ( n5548 ) | ( n5595 )  ;
assign n5597 =  ( n5515 ) ^ ( n5531 )  ;
assign n5598 = ~ ( n5597 ) ;
assign n5599 =  ( n5596 ) | ( n5598 )  ;
assign n5600 = ~ ( n5599 ) ;
assign n5601 =  ( n5539 ) | ( n5600 )  ;
assign n5602 = ~ ( n5601 ) ;
assign n5603 =  ( n5495 ) | ( n5602 )  ;
assign n5604 = ~ ( n5603 ) ;
assign n5605 =  ( n5474 ) | ( n5604 )  ;
assign n5606 =  ( n5452 ) ^ ( n5325 )  ;
assign n5607 =  ( n5606 ) ^ ( n5083 )  ;
assign n5608 =  ( n5607 ) ^ ( n5099 )  ;
assign n5609 =  ( n5608 ) ^ ( n5116 )  ;
assign n5610 =  ( n5609 ) ^ ( n5141 )  ;
assign n5611 =  ( n5610 ) ^ ( n5129 )  ;
assign n5612 = ~ ( n5611 ) ;
assign n5613 =  ( n5489 ) ^ ( n5433 )  ;
assign n5614 =  ( n5613 ) ^ ( n5285 )  ;
assign n5615 =  ( n5614 ) ^ ( n5301 )  ;
assign n5616 =  ( n5615 ) ^ ( n5321 )  ;
assign n5617 = ~ ( n5616 ) ;
assign n5618 =  ( n5612 ) | ( n5617 )  ;
assign n5619 = ~ ( n5547 ) ;
assign n5620 =  ( n5618 ) | ( n5619 )  ;
assign n5621 =  ( n5594 ) ^ ( n5515 )  ;
assign n5622 =  ( n5621 ) ^ ( n5531 )  ;
assign n5623 = ~ ( n5622 ) ;
assign n5624 =  ( n5620 ) | ( n5623 )  ;
assign n5625 =  ( n5568 ) ^ ( n5583 )  ;
assign n5626 =  ( n5625 ) ^ ( n5580 )  ;
assign n5627 = ~ ( n5626 ) ;
assign n5628 =  ( n5624 ) | ( n5627 )  ;
assign n5629 = ki[0:0] ;
assign n5630 =  ( n5629 ) == ( bv_1_1_n5 )  ;
assign n5631 = ki[1:1] ;
assign n5632 =  ( n5631 ) == ( bv_1_0_n2 )  ;
assign n5633 =  ( n5630 ) | ( n5632 )  ;
assign n5634 = ki[1:1] ;
assign n5635 =  ( n5634 ) == ( bv_1_1_n5 )  ;
assign n5636 = ki[0:0] ;
assign n5637 =  ( n5636 ) == ( bv_1_1_n5 )  ;
assign n5638 =  ( n5635 ) | ( n5637 )  ;
assign n5639 = ki[1:1] ;
assign n5640 =  ( n5639 ) == ( bv_1_1_n5 )  ;
assign n5641 = i_wb_data[0:0] ;
assign n5642 = ~ ( n5641 ) ;
assign n5643 =  ( bv_1_1_n5 ) ^ ( n5642 )  ;
assign n5644 = sp[0:0] ;
assign n5645 =  ( n5643 ) ^ ( n5644 )  ;
assign n5646 =  ( n5640 ) ? ( n2910 ) : ( n5645 ) ;
assign n5647 =  ( n5638 ) ? ( n5646 ) : ( bv_1_0_n2 ) ;
assign n5648 =  ( n5633 ) ? ( n5567 ) : ( n5647 ) ;
assign n5649 = ~ ( n5648 ) ;
assign n5650 =  ( n5628 ) | ( n5649 )  ;
assign n5651 = ki[0:0] ;
assign n5652 =  ( n5651 ) == ( bv_1_1_n5 )  ;
assign n5653 = ki[1:1] ;
assign n5654 =  ( n5653 ) == ( bv_1_0_n2 )  ;
assign n5655 =  ( n5652 ) | ( n5654 )  ;
assign n5656 = ki[1:1] ;
assign n5657 =  ( n5655 ) ? ( n5647 ) : ( n5656 ) ;
assign n5658 = ~ ( n5657 ) ;
assign n5659 =  ( n5650 ) | ( n5658 )  ;
assign n5660 = ki[1:1] ;
assign n5661 = ~ ( n5660 ) ;
assign n5662 =  ( n5659 ) | ( n5661 )  ;
assign n5663 = ~ ( n5662 ) ;
assign n5664 =  ( n5605 ) | ( n5663 )  ;
assign n5665 = ~ ( n5664 ) ;
assign n5666 =  ( n5374 ) | ( n5665 )  ;
assign n5667 = ~ ( n5666 ) ;
assign n5668 =  ( n5350 ) | ( n5667 )  ;
assign n5669 = ~ ( n5668 ) ;
assign n5670 =  ( n4254 ) | ( n5669 )  ;
assign n5671 = ~ ( n5670 ) ;
assign n5672 =  ( n4194 ) | ( n5671 )  ;
assign n5673 = ~ ( n5672 ) ;
assign n5674 = kd[13:13] ;
assign n5675 =  ( n5674 ) == ( bv_1_0_n2 )  ;
assign n5676 = kd[12:12] ;
assign n5677 =  ( n5676 ) == ( bv_1_0_n2 )  ;
assign n5678 =  ( n5675 ) | ( n5677 )  ;
assign n5679 = kd[11:11] ;
assign n5680 =  ( n5679 ) == ( bv_1_0_n2 )  ;
assign n5681 =  ( n5678 ) | ( n5680 )  ;
assign n5682 = ~ ( n5681 )  ;
assign n5683 = kd[13:13] ;
assign n5684 =  ( n5683 ) == ( bv_1_1_n5 )  ;
assign n5685 = kd[12:12] ;
assign n5686 =  ( n5685 ) == ( bv_1_1_n5 )  ;
assign n5687 =  ( n5684 ) | ( n5686 )  ;
assign n5688 = kd[11:11] ;
assign n5689 =  ( n5688 ) == ( bv_1_1_n5 )  ;
assign n5690 =  ( n5687 ) | ( n5689 )  ;
assign n5691 = ~ ( n5690 )  ;
assign n5692 =  ( n5682 ) | ( n5691 )  ;
assign n5693 = kd[13:13] ;
assign n5694 =  ( n5693 ) == ( bv_1_0_n2 )  ;
assign n5695 = kd[12:12] ;
assign n5696 =  ( n5695 ) == ( bv_1_0_n2 )  ;
assign n5697 = kd[11:11] ;
assign n5698 =  ( n5697 ) == ( bv_1_0_n2 )  ;
assign n5699 =  ( n5696 ) | ( n5698 )  ;
assign n5700 = ~ ( n5699 )  ;
assign n5701 =  ( n5694 ) | ( n5700 )  ;
assign n5702 =  ( n5701 ) ? ( bv_1_0_n2 ) : ( bv_1_1_n5 ) ;
assign n5703 =  ( n5692 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5704 = ~ ( n5703 ) ;
assign n5705 = kd[15:15] ;
assign n5706 =  ( n5705 ) == ( bv_1_0_n2 )  ;
assign n5707 = kd[14:14] ;
assign n5708 =  ( n5707 ) == ( bv_1_0_n2 )  ;
assign n5709 =  ( n5706 ) | ( n5708 )  ;
assign n5710 = kd[13:13] ;
assign n5711 =  ( n5710 ) == ( bv_1_0_n2 )  ;
assign n5712 =  ( n5709 ) | ( n5711 )  ;
assign n5713 = ~ ( n5712 )  ;
assign n5714 = kd[14:14] ;
assign n5715 =  ( n5714 ) == ( bv_1_1_n5 )  ;
assign n5716 = kd[13:13] ;
assign n5717 =  ( n5716 ) == ( bv_1_1_n5 )  ;
assign n5718 =  ( n5715 ) | ( n5717 )  ;
assign n5719 = kd[15:15] ;
assign n5720 =  ( n5719 ) == ( bv_1_1_n5 )  ;
assign n5721 =  ( n5718 ) | ( n5720 )  ;
assign n5722 = ~ ( n5721 )  ;
assign n5723 =  ( n5713 ) | ( n5722 )  ;
assign n5724 = kd[15:15] ;
assign n5725 =  ( n5724 ) == ( bv_1_0_n2 )  ;
assign n5726 = kd[14:14] ;
assign n5727 =  ( n5726 ) == ( bv_1_0_n2 )  ;
assign n5728 = kd[13:13] ;
assign n5729 =  ( n5728 ) == ( bv_1_0_n2 )  ;
assign n5730 =  ( n5727 ) | ( n5729 )  ;
assign n5731 = ~ ( n5730 )  ;
assign n5732 =  ( n5725 ) | ( n5731 )  ;
assign n5733 =  ( n5732 ) ? ( bv_1_0_n2 ) : ( bv_1_1_n5 ) ;
assign n5734 =  ( n5723 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5735 = ~ ( n5734 ) ;
assign n5736 =  ( n5704 ) | ( n5735 )  ;
assign n5737 = ~ ( n5736 ) ;
assign n5738 =  ( n5682 ) | ( n5691 )  ;
assign n5739 =  ( n5738 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5740 =  ( n5713 ) | ( n5722 )  ;
assign n5741 =  ( n5740 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5742 =  ( n5739 ) ^ ( n5741 )  ;
assign n5743 =  ( n5737 ) | ( n5742 )  ;
assign n5744 = ~ ( n5743 ) ;
assign n5745 =  ( n5682 ) | ( n5691 )  ;
assign n5746 =  ( n5745 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5747 =  ( n5744 ) | ( n5746 )  ;
assign n5748 = ~ ( n5747 ) ;
assign n5749 = ~ ( n5736 ) ;
assign n5750 =  ( n5749 ) | ( n5742 )  ;
assign n5751 =  ( n5682 ) | ( n5691 )  ;
assign n5752 =  ( n5751 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5753 = ~ ( n5752 ) ;
assign n5754 =  ( n5750 ) ^ ( n5753 )  ;
assign n5755 = ~ ( n5754 ) ;
assign n5756 =  ( n5713 ) | ( n5722 )  ;
assign n5757 =  ( n5756 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5758 = ~ ( n5757 ) ;
assign n5759 =  ( n5755 ) | ( n5758 )  ;
assign n5760 = ~ ( n5759 ) ;
assign n5761 =  ( n5748 ) | ( n5760 )  ;
assign n5762 = ~ ( n5761 ) ;
assign n5763 =  ( n5713 ) | ( n5722 )  ;
assign n5764 =  ( n5763 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5765 = ~ ( n5764 ) ;
assign n5766 =  ( n5762 ) | ( n5765 )  ;
assign n5767 = ~ ( n5766 ) ;
assign n5768 = ~ ( n5747 ) ;
assign n5769 = ~ ( n5759 ) ;
assign n5770 =  ( n5768 ) | ( n5769 )  ;
assign n5771 =  ( n5713 ) | ( n5722 )  ;
assign n5772 =  ( n5771 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5773 =  ( n5770 ) ^ ( n5772 )  ;
assign n5774 =  ( n5767 ) | ( n5773 )  ;
assign n5775 = ~ ( n5774 ) ;
assign n5776 =  ( n5713 ) | ( n5722 )  ;
assign n5777 =  ( n5776 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5778 =  ( n5775 ) | ( n5777 )  ;
assign n5779 = ~ ( n5778 ) ;
assign n5780 =  ( n5713 ) | ( n5722 )  ;
assign n5781 =  ( n5780 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5782 = ~ ( n5781 ) ;
assign n5783 =  ( n5774 ) ^ ( n5782 )  ;
assign n5784 = ~ ( n5783 ) ;
assign n5785 = ~ ( n5747 ) ;
assign n5786 = ~ ( n5759 ) ;
assign n5787 =  ( n5785 ) | ( n5786 )  ;
assign n5788 =  ( bv_1_1_n5 ) ^ ( n5787 )  ;
assign n5789 =  ( n5713 ) | ( n5722 )  ;
assign n5790 =  ( n5789 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5791 =  ( n5788 ) ^ ( n5790 )  ;
assign n5792 = ~ ( n5791 ) ;
assign n5793 =  ( n5784 ) | ( n5792 )  ;
assign n5794 = kd[9:9] ;
assign n5795 =  ( n5794 ) == ( bv_1_0_n2 )  ;
assign n5796 = kd[8:8] ;
assign n5797 =  ( n5796 ) == ( bv_1_0_n2 )  ;
assign n5798 =  ( n5795 ) | ( n5797 )  ;
assign n5799 = kd[7:7] ;
assign n5800 =  ( n5799 ) == ( bv_1_0_n2 )  ;
assign n5801 =  ( n5798 ) | ( n5800 )  ;
assign n5802 = ~ ( n5801 )  ;
assign n5803 = kd[9:9] ;
assign n5804 =  ( n5803 ) == ( bv_1_1_n5 )  ;
assign n5805 = kd[8:8] ;
assign n5806 =  ( n5805 ) == ( bv_1_1_n5 )  ;
assign n5807 =  ( n5804 ) | ( n5806 )  ;
assign n5808 = kd[7:7] ;
assign n5809 =  ( n5808 ) == ( bv_1_1_n5 )  ;
assign n5810 =  ( n5807 ) | ( n5809 )  ;
assign n5811 = ~ ( n5810 )  ;
assign n5812 =  ( n5802 ) | ( n5811 )  ;
assign n5813 = kd[9:9] ;
assign n5814 =  ( n5813 ) == ( bv_1_0_n2 )  ;
assign n5815 = kd[8:8] ;
assign n5816 =  ( n5815 ) == ( bv_1_0_n2 )  ;
assign n5817 = kd[7:7] ;
assign n5818 =  ( n5817 ) == ( bv_1_0_n2 )  ;
assign n5819 =  ( n5816 ) | ( n5818 )  ;
assign n5820 = ~ ( n5819 )  ;
assign n5821 =  ( n5814 ) | ( n5820 )  ;
assign n5822 =  ( n5821 ) ? ( bv_1_0_n2 ) : ( bv_1_1_n5 ) ;
assign n5823 =  ( n5812 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n5824 = kd[11:11] ;
assign n5825 =  ( n5824 ) == ( bv_1_0_n2 )  ;
assign n5826 = kd[10:10] ;
assign n5827 =  ( n5826 ) == ( bv_1_0_n2 )  ;
assign n5828 =  ( n5825 ) | ( n5827 )  ;
assign n5829 = kd[9:9] ;
assign n5830 =  ( n5829 ) == ( bv_1_0_n2 )  ;
assign n5831 =  ( n5828 ) | ( n5830 )  ;
assign n5832 = ~ ( n5831 )  ;
assign n5833 = kd[11:11] ;
assign n5834 =  ( n5833 ) == ( bv_1_1_n5 )  ;
assign n5835 = kd[10:10] ;
assign n5836 =  ( n5835 ) == ( bv_1_1_n5 )  ;
assign n5837 =  ( n5834 ) | ( n5836 )  ;
assign n5838 = kd[9:9] ;
assign n5839 =  ( n5838 ) == ( bv_1_1_n5 )  ;
assign n5840 =  ( n5837 ) | ( n5839 )  ;
assign n5841 = ~ ( n5840 )  ;
assign n5842 =  ( n5832 ) | ( n5841 )  ;
assign n5843 = kd[11:11] ;
assign n5844 =  ( n5843 ) == ( bv_1_0_n2 )  ;
assign n5845 = kd[10:10] ;
assign n5846 =  ( n5845 ) == ( bv_1_0_n2 )  ;
assign n5847 = kd[9:9] ;
assign n5848 =  ( n5847 ) == ( bv_1_0_n2 )  ;
assign n5849 =  ( n5846 ) | ( n5848 )  ;
assign n5850 = ~ ( n5849 )  ;
assign n5851 =  ( n5844 ) | ( n5850 )  ;
assign n5852 =  ( n5851 ) ? ( bv_1_0_n2 ) : ( bv_1_1_n5 ) ;
assign n5853 =  ( n5842 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5854 = ~ ( n5853 ) ;
assign n5855 =  ( n5823 ) | ( n5854 )  ;
assign n5856 = ~ ( n5855 ) ;
assign n5857 =  ( n5802 ) | ( n5811 )  ;
assign n5858 =  ( n5857 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n5859 = ~ ( n5858 ) ;
assign n5860 =  ( n5832 ) | ( n5841 )  ;
assign n5861 =  ( n5860 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5862 =  ( n5859 ) ^ ( n5861 )  ;
assign n5863 = ~ ( n5862 ) ;
assign n5864 =  ( n5682 ) | ( n5691 )  ;
assign n5865 =  ( n5864 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5866 = ~ ( n5865 ) ;
assign n5867 =  ( n5863 ) | ( n5866 )  ;
assign n5868 = ~ ( n5867 ) ;
assign n5869 =  ( n5856 ) | ( n5868 )  ;
assign n5870 = ~ ( n5869 ) ;
assign n5871 =  ( n5832 ) | ( n5841 )  ;
assign n5872 =  ( n5871 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5873 =  ( n5682 ) | ( n5691 )  ;
assign n5874 =  ( n5873 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5875 =  ( n5872 ) ^ ( n5874 )  ;
assign n5876 =  ( n5713 ) | ( n5722 )  ;
assign n5877 =  ( n5876 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5878 =  ( n5875 ) ^ ( n5877 )  ;
assign n5879 = ~ ( n5878 ) ;
assign n5880 =  ( n5870 ) | ( n5879 )  ;
assign n5881 = ~ ( n5880 ) ;
assign n5882 = ~ ( n5855 ) ;
assign n5883 = ~ ( n5867 ) ;
assign n5884 =  ( n5882 ) | ( n5883 )  ;
assign n5885 =  ( n5832 ) | ( n5841 )  ;
assign n5886 =  ( n5885 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5887 =  ( n5884 ) ^ ( n5886 )  ;
assign n5888 =  ( n5682 ) | ( n5691 )  ;
assign n5889 =  ( n5888 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5890 =  ( n5887 ) ^ ( n5889 )  ;
assign n5891 =  ( n5713 ) | ( n5722 )  ;
assign n5892 =  ( n5891 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5893 =  ( n5890 ) ^ ( n5892 )  ;
assign n5894 =  ( n5881 ) | ( n5893 )  ;
assign n5895 = ~ ( n5894 ) ;
assign n5896 =  ( n5832 ) | ( n5841 )  ;
assign n5897 =  ( n5896 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5898 = ~ ( n5897 ) ;
assign n5899 =  ( n5682 ) | ( n5691 )  ;
assign n5900 =  ( n5899 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5901 = ~ ( n5900 ) ;
assign n5902 =  ( n5898 ) | ( n5901 )  ;
assign n5903 = ~ ( n5902 ) ;
assign n5904 =  ( n5832 ) | ( n5841 )  ;
assign n5905 =  ( n5904 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5906 =  ( n5682 ) | ( n5691 )  ;
assign n5907 =  ( n5906 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5908 =  ( n5905 ) ^ ( n5907 )  ;
assign n5909 = ~ ( n5908 ) ;
assign n5910 =  ( n5713 ) | ( n5722 )  ;
assign n5911 =  ( n5910 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5912 = ~ ( n5911 ) ;
assign n5913 =  ( n5909 ) | ( n5912 )  ;
assign n5914 = ~ ( n5913 ) ;
assign n5915 =  ( n5903 ) | ( n5914 )  ;
assign n5916 = ~ ( n5915 ) ;
assign n5917 =  ( n5895 ) | ( n5916 )  ;
assign n5918 = ~ ( n5917 ) ;
assign n5919 = ~ ( n5902 ) ;
assign n5920 = ~ ( n5913 ) ;
assign n5921 =  ( n5919 ) | ( n5920 )  ;
assign n5922 =  ( n5894 ) ^ ( n5921 )  ;
assign n5923 = ~ ( n5922 ) ;
assign n5924 =  ( n5832 ) | ( n5841 )  ;
assign n5925 =  ( n5924 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5926 = ~ ( n5925 ) ;
assign n5927 =  ( n5682 ) | ( n5691 )  ;
assign n5928 =  ( n5927 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5929 =  ( n5926 ) ^ ( n5928 )  ;
assign n5930 =  ( n5713 ) | ( n5722 )  ;
assign n5931 =  ( n5930 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5932 =  ( n5929 ) ^ ( n5931 )  ;
assign n5933 = ~ ( n5932 ) ;
assign n5934 =  ( n5923 ) | ( n5933 )  ;
assign n5935 = ~ ( n5934 ) ;
assign n5936 =  ( n5918 ) | ( n5935 )  ;
assign n5937 = ~ ( n5936 ) ;
assign n5938 =  ( n5832 ) | ( n5841 )  ;
assign n5939 =  ( n5938 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5940 =  ( n5682 ) | ( n5691 )  ;
assign n5941 =  ( n5940 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5942 = ~ ( n5941 ) ;
assign n5943 =  ( n5939 ) | ( n5942 )  ;
assign n5944 = ~ ( n5943 ) ;
assign n5945 =  ( n5832 ) | ( n5841 )  ;
assign n5946 =  ( n5945 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n5947 = ~ ( n5946 ) ;
assign n5948 =  ( n5682 ) | ( n5691 )  ;
assign n5949 =  ( n5948 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5950 =  ( n5947 ) ^ ( n5949 )  ;
assign n5951 = ~ ( n5950 ) ;
assign n5952 =  ( n5713 ) | ( n5722 )  ;
assign n5953 =  ( n5952 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5954 = ~ ( n5953 ) ;
assign n5955 =  ( n5951 ) | ( n5954 )  ;
assign n5956 = ~ ( n5955 ) ;
assign n5957 =  ( n5944 ) | ( n5956 )  ;
assign n5958 = ~ ( n5957 ) ;
assign n5959 =  ( n5937 ) | ( n5958 )  ;
assign n5960 = ~ ( n5959 ) ;
assign n5961 = ~ ( n5943 ) ;
assign n5962 = ~ ( n5955 ) ;
assign n5963 =  ( n5961 ) | ( n5962 )  ;
assign n5964 =  ( n5936 ) ^ ( n5963 )  ;
assign n5965 = ~ ( n5964 ) ;
assign n5966 =  ( n5682 ) | ( n5691 )  ;
assign n5967 =  ( n5966 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5968 =  ( bv_1_1_n5 ) ^ ( n5967 )  ;
assign n5969 =  ( n5713 ) | ( n5722 )  ;
assign n5970 =  ( n5969 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5971 =  ( n5968 ) ^ ( n5970 )  ;
assign n5972 = ~ ( n5971 ) ;
assign n5973 =  ( n5965 ) | ( n5972 )  ;
assign n5974 = ~ ( n5973 ) ;
assign n5975 =  ( n5960 ) | ( n5974 )  ;
assign n5976 = ~ ( n5975 ) ;
assign n5977 =  ( n5793 ) | ( n5976 )  ;
assign n5978 = ~ ( n5736 ) ;
assign n5979 =  ( n5978 ) | ( n5742 )  ;
assign n5980 =  ( n5682 ) | ( n5691 )  ;
assign n5981 =  ( n5980 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n5982 = ~ ( n5981 ) ;
assign n5983 =  ( n5979 ) ^ ( n5982 )  ;
assign n5984 =  ( n5713 ) | ( n5722 )  ;
assign n5985 =  ( n5984 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n5986 =  ( n5983 ) ^ ( n5985 )  ;
assign n5987 = ~ ( n5986 ) ;
assign n5988 =  ( n5977 ) | ( n5987 )  ;
assign n5989 = ~ ( n5988 ) ;
assign n5990 =  ( n5779 ) | ( n5989 )  ;
assign n5991 = ~ ( n5783 ) ;
assign n5992 =  ( n5991 ) | ( n5792 )  ;
assign n5993 = ~ ( n5959 ) ;
assign n5994 =  ( n5965 ) | ( n5972 )  ;
assign n5995 = ~ ( n5994 ) ;
assign n5996 =  ( n5993 ) | ( n5995 )  ;
assign n5997 = ~ ( n5736 ) ;
assign n5998 =  ( n5997 ) | ( n5742 )  ;
assign n5999 =  ( n5996 ) ^ ( n5998 )  ;
assign n6000 =  ( n5682 ) | ( n5691 )  ;
assign n6001 =  ( n6000 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6002 = ~ ( n6001 ) ;
assign n6003 =  ( n5999 ) ^ ( n6002 )  ;
assign n6004 =  ( n5713 ) | ( n5722 )  ;
assign n6005 =  ( n6004 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6006 =  ( n6003 ) ^ ( n6005 )  ;
assign n6007 = ~ ( n6006 ) ;
assign n6008 =  ( n5992 ) | ( n6007 )  ;
assign n6009 =  ( bv_1_1_n5 ) ^ ( n5936 )  ;
assign n6010 = ~ ( n5943 ) ;
assign n6011 = ~ ( n5955 ) ;
assign n6012 =  ( n6010 ) | ( n6011 )  ;
assign n6013 =  ( n6009 ) ^ ( n6012 )  ;
assign n6014 =  ( n5682 ) | ( n5691 )  ;
assign n6015 =  ( n6014 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6016 =  ( n6013 ) ^ ( n6015 )  ;
assign n6017 =  ( n5713 ) | ( n5722 )  ;
assign n6018 =  ( n6017 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6019 =  ( n6016 ) ^ ( n6018 )  ;
assign n6020 = ~ ( n6019 ) ;
assign n6021 =  ( n6008 ) | ( n6020 )  ;
assign n6022 = kd[7:7] ;
assign n6023 =  ( n6022 ) == ( bv_1_0_n2 )  ;
assign n6024 = kd[6:6] ;
assign n6025 =  ( n6024 ) == ( bv_1_0_n2 )  ;
assign n6026 =  ( n6023 ) | ( n6025 )  ;
assign n6027 = kd[5:5] ;
assign n6028 =  ( n6027 ) == ( bv_1_0_n2 )  ;
assign n6029 =  ( n6026 ) | ( n6028 )  ;
assign n6030 = ~ ( n6029 )  ;
assign n6031 = kd[7:7] ;
assign n6032 =  ( n6031 ) == ( bv_1_1_n5 )  ;
assign n6033 = kd[6:6] ;
assign n6034 =  ( n6033 ) == ( bv_1_1_n5 )  ;
assign n6035 =  ( n6032 ) | ( n6034 )  ;
assign n6036 = kd[5:5] ;
assign n6037 =  ( n6036 ) == ( bv_1_1_n5 )  ;
assign n6038 =  ( n6035 ) | ( n6037 )  ;
assign n6039 = ~ ( n6038 )  ;
assign n6040 =  ( n6030 ) | ( n6039 )  ;
assign n6041 = kd[7:7] ;
assign n6042 =  ( n6041 ) == ( bv_1_0_n2 )  ;
assign n6043 = kd[6:6] ;
assign n6044 =  ( n6043 ) == ( bv_1_0_n2 )  ;
assign n6045 = kd[5:5] ;
assign n6046 =  ( n6045 ) == ( bv_1_0_n2 )  ;
assign n6047 =  ( n6044 ) | ( n6046 )  ;
assign n6048 = ~ ( n6047 )  ;
assign n6049 =  ( n6042 ) | ( n6048 )  ;
assign n6050 =  ( n6049 ) ? ( bv_1_0_n2 ) : ( bv_1_1_n5 ) ;
assign n6051 =  ( n6040 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6052 =  ( n5802 ) | ( n5811 )  ;
assign n6053 =  ( n6052 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6054 = ~ ( n6053 ) ;
assign n6055 =  ( n6051 ) | ( n6054 )  ;
assign n6056 =  ( n5832 ) | ( n5841 )  ;
assign n6057 =  ( n6056 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6058 = ~ ( n6057 ) ;
assign n6059 =  ( n6055 ) | ( n6058 )  ;
assign n6060 =  ( n5682 ) | ( n5691 )  ;
assign n6061 =  ( n6060 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6062 = ~ ( n6061 ) ;
assign n6063 =  ( n6059 ) | ( n6062 )  ;
assign n6064 = ~ ( n6063 ) ;
assign n6065 =  ( n6030 ) | ( n6039 )  ;
assign n6066 =  ( n6065 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6067 = ~ ( n6066 ) ;
assign n6068 =  ( n5802 ) | ( n5811 )  ;
assign n6069 =  ( n6068 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6070 =  ( n6067 ) ^ ( n6069 )  ;
assign n6071 = ~ ( n6070 ) ;
assign n6072 =  ( n6071 ) | ( n5909 )  ;
assign n6073 = ~ ( n6072 ) ;
assign n6074 =  ( n6064 ) | ( n6073 )  ;
assign n6075 =  ( n6030 ) | ( n6039 )  ;
assign n6076 =  ( n6075 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6077 = ~ ( n6076 ) ;
assign n6078 =  ( n5802 ) | ( n5811 )  ;
assign n6079 =  ( n6078 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6080 =  ( n6077 ) ^ ( n6079 )  ;
assign n6081 =  ( n5832 ) | ( n5841 )  ;
assign n6082 =  ( n6081 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6083 =  ( n6080 ) ^ ( n6082 )  ;
assign n6084 =  ( n5682 ) | ( n5691 )  ;
assign n6085 =  ( n6084 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6086 =  ( n6083 ) ^ ( n6085 )  ;
assign n6087 = ~ ( n6086 ) ;
assign n6088 =  ( n5713 ) | ( n5722 )  ;
assign n6089 =  ( n6088 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6090 = ~ ( n6089 ) ;
assign n6091 =  ( n6087 ) | ( n6090 )  ;
assign n6092 = ~ ( n6091 ) ;
assign n6093 =  ( n6074 ) | ( n6092 )  ;
assign n6094 = ~ ( n6093 ) ;
assign n6095 =  ( n6030 ) | ( n6039 )  ;
assign n6096 =  ( n6095 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6097 =  ( n5802 ) | ( n5811 )  ;
assign n6098 =  ( n6097 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6099 = ~ ( n6098 ) ;
assign n6100 =  ( n6096 ) | ( n6099 )  ;
assign n6101 = ~ ( n6100 ) ;
assign n6102 = ~ ( n5902 ) ;
assign n6103 =  ( n6101 ) | ( n6102 )  ;
assign n6104 = ~ ( n6103 ) ;
assign n6105 =  ( n6094 ) | ( n6104 )  ;
assign n6106 = ~ ( n6105 ) ;
assign n6107 = ~ ( n6100 ) ;
assign n6108 = ~ ( n5902 ) ;
assign n6109 =  ( n6107 ) | ( n6108 )  ;
assign n6110 =  ( n6093 ) ^ ( n6109 )  ;
assign n6111 = ~ ( n6110 ) ;
assign n6112 =  ( n5802 ) | ( n5811 )  ;
assign n6113 =  ( n6112 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6114 =  ( bv_1_1_n5 ) ^ ( n6113 )  ;
assign n6115 =  ( n5832 ) | ( n5841 )  ;
assign n6116 =  ( n6115 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6117 =  ( n6114 ) ^ ( n6116 )  ;
assign n6118 =  ( n5682 ) | ( n5691 )  ;
assign n6119 =  ( n6118 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6120 =  ( n6117 ) ^ ( n6119 )  ;
assign n6121 =  ( n5713 ) | ( n5722 )  ;
assign n6122 =  ( n6121 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6123 =  ( n6120 ) ^ ( n6122 )  ;
assign n6124 = ~ ( n6123 ) ;
assign n6125 =  ( n6111 ) | ( n6124 )  ;
assign n6126 = ~ ( n6125 ) ;
assign n6127 =  ( n6106 ) | ( n6126 )  ;
assign n6128 = ~ ( n6127 ) ;
assign n6129 =  ( n5802 ) | ( n5811 )  ;
assign n6130 =  ( n6129 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6131 = ~ ( n6130 ) ;
assign n6132 =  ( n5832 ) | ( n5841 )  ;
assign n6133 =  ( n6132 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6134 = ~ ( n6133 ) ;
assign n6135 =  ( n6131 ) | ( n6134 )  ;
assign n6136 =  ( n5682 ) | ( n5691 )  ;
assign n6137 =  ( n6136 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6138 = ~ ( n6137 ) ;
assign n6139 =  ( n6135 ) | ( n6138 )  ;
assign n6140 =  ( n5713 ) | ( n5722 )  ;
assign n6141 =  ( n6140 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6142 = ~ ( n6141 ) ;
assign n6143 =  ( n6139 ) | ( n6142 )  ;
assign n6144 = ~ ( n6143 ) ;
assign n6145 =  ( n5802 ) | ( n5811 )  ;
assign n6146 =  ( n6145 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6147 =  ( n5832 ) | ( n5841 )  ;
assign n6148 =  ( n6147 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6149 =  ( n6146 ) ^ ( n6148 )  ;
assign n6150 = ~ ( n6149 ) ;
assign n6151 = ~ ( n5742 ) ;
assign n6152 =  ( n6150 ) | ( n6151 )  ;
assign n6153 = ~ ( n6152 ) ;
assign n6154 =  ( n6144 ) | ( n6153 )  ;
assign n6155 =  ( n5802 ) | ( n5811 )  ;
assign n6156 =  ( n6155 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6157 =  ( n5832 ) | ( n5841 )  ;
assign n6158 =  ( n6157 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6159 =  ( n6156 ) ^ ( n6158 )  ;
assign n6160 =  ( n5682 ) | ( n5691 )  ;
assign n6161 =  ( n6160 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6162 =  ( n6159 ) ^ ( n6161 )  ;
assign n6163 =  ( n5713 ) | ( n5722 )  ;
assign n6164 =  ( n6163 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6165 =  ( n6162 ) ^ ( n6164 )  ;
assign n6166 =  ( n6154 ) | ( n6165 )  ;
assign n6167 =  ( n5802 ) | ( n5811 )  ;
assign n6168 =  ( n6167 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6169 = ~ ( n6168 ) ;
assign n6170 =  ( n5832 ) | ( n5841 )  ;
assign n6171 =  ( n6170 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6172 = ~ ( n6171 ) ;
assign n6173 =  ( n6169 ) | ( n6172 )  ;
assign n6174 = ~ ( n6173 ) ;
assign n6175 = ~ ( n5736 ) ;
assign n6176 =  ( n6174 ) | ( n6175 )  ;
assign n6177 =  ( n6166 ) ^ ( n6176 )  ;
assign n6178 =  ( n5802 ) | ( n5811 )  ;
assign n6179 =  ( n6178 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6180 = ~ ( n6179 ) ;
assign n6181 =  ( n6177 ) ^ ( n6180 )  ;
assign n6182 =  ( n5832 ) | ( n5841 )  ;
assign n6183 =  ( n6182 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6184 =  ( n6181 ) ^ ( n6183 )  ;
assign n6185 =  ( n5682 ) | ( n5691 )  ;
assign n6186 =  ( n6185 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6187 =  ( n6184 ) ^ ( n6186 )  ;
assign n6188 = ~ ( n6187 ) ;
assign n6189 =  ( n6128 ) | ( n6188 )  ;
assign n6190 = ~ ( n6189 ) ;
assign n6191 = ~ ( n6105 ) ;
assign n6192 =  ( n6111 ) | ( n6124 )  ;
assign n6193 = ~ ( n6192 ) ;
assign n6194 =  ( n6191 ) | ( n6193 )  ;
assign n6195 =  ( n6194 ) ^ ( n6166 )  ;
assign n6196 = ~ ( n6173 ) ;
assign n6197 = ~ ( n5736 ) ;
assign n6198 =  ( n6196 ) | ( n6197 )  ;
assign n6199 =  ( n6195 ) ^ ( n6198 )  ;
assign n6200 =  ( n5802 ) | ( n5811 )  ;
assign n6201 =  ( n6200 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6202 = ~ ( n6201 ) ;
assign n6203 =  ( n6199 ) ^ ( n6202 )  ;
assign n6204 =  ( n5832 ) | ( n5841 )  ;
assign n6205 =  ( n6204 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6206 =  ( n6203 ) ^ ( n6205 )  ;
assign n6207 =  ( n5682 ) | ( n5691 )  ;
assign n6208 =  ( n6207 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6209 =  ( n6206 ) ^ ( n6208 )  ;
assign n6210 = ~ ( n6209 ) ;
assign n6211 =  ( n5713 ) | ( n5722 )  ;
assign n6212 =  ( n6211 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6213 = ~ ( n6212 ) ;
assign n6214 =  ( n6210 ) | ( n6213 )  ;
assign n6215 = ~ ( n6214 ) ;
assign n6216 =  ( n6190 ) | ( n6215 )  ;
assign n6217 = ~ ( n6216 ) ;
assign n6218 = ~ ( n6166 ) ;
assign n6219 = ~ ( n6173 ) ;
assign n6220 = ~ ( n5736 ) ;
assign n6221 =  ( n6219 ) | ( n6220 )  ;
assign n6222 = ~ ( n6221 ) ;
assign n6223 =  ( n6218 ) | ( n6222 )  ;
assign n6224 = ~ ( n6223 ) ;
assign n6225 = ~ ( n6173 ) ;
assign n6226 = ~ ( n5736 ) ;
assign n6227 =  ( n6225 ) | ( n6226 )  ;
assign n6228 =  ( n6166 ) ^ ( n6227 )  ;
assign n6229 = ~ ( n6228 ) ;
assign n6230 =  ( n5802 ) | ( n5811 )  ;
assign n6231 =  ( n6230 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6232 = ~ ( n6231 ) ;
assign n6233 =  ( n5832 ) | ( n5841 )  ;
assign n6234 =  ( n6233 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6235 =  ( n6232 ) ^ ( n6234 )  ;
assign n6236 =  ( n5682 ) | ( n5691 )  ;
assign n6237 =  ( n6236 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6238 =  ( n6235 ) ^ ( n6237 )  ;
assign n6239 = ~ ( n6238 ) ;
assign n6240 =  ( n6229 ) | ( n6239 )  ;
assign n6241 = ~ ( n6240 ) ;
assign n6242 =  ( n6224 ) | ( n6241 )  ;
assign n6243 = ~ ( n6242 ) ;
assign n6244 =  ( n6217 ) | ( n6243 )  ;
assign n6245 = ~ ( n6244 ) ;
assign n6246 =  ( n6216 ) ^ ( n6242 )  ;
assign n6247 = ~ ( n6246 ) ;
assign n6248 = ~ ( n5855 ) ;
assign n6249 = ~ ( n5867 ) ;
assign n6250 =  ( n6248 ) | ( n6249 )  ;
assign n6251 =  ( bv_1_1_n5 ) ^ ( n6250 )  ;
assign n6252 =  ( n5832 ) | ( n5841 )  ;
assign n6253 =  ( n6252 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6254 =  ( n6251 ) ^ ( n6253 )  ;
assign n6255 =  ( n5682 ) | ( n5691 )  ;
assign n6256 =  ( n6255 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6257 =  ( n6254 ) ^ ( n6256 )  ;
assign n6258 =  ( n5713 ) | ( n5722 )  ;
assign n6259 =  ( n6258 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6260 =  ( n6257 ) ^ ( n6259 )  ;
assign n6261 = ~ ( n6260 ) ;
assign n6262 =  ( n6247 ) | ( n6261 )  ;
assign n6263 = ~ ( n6262 ) ;
assign n6264 =  ( n6245 ) | ( n6263 )  ;
assign n6265 = ~ ( n6264 ) ;
assign n6266 = ~ ( n5902 ) ;
assign n6267 = ~ ( n5913 ) ;
assign n6268 =  ( n6266 ) | ( n6267 )  ;
assign n6269 =  ( n5894 ) ^ ( n6268 )  ;
assign n6270 =  ( n5832 ) | ( n5841 )  ;
assign n6271 =  ( n6270 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6272 = ~ ( n6271 ) ;
assign n6273 =  ( n6269 ) ^ ( n6272 )  ;
assign n6274 =  ( n5682 ) | ( n5691 )  ;
assign n6275 =  ( n6274 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6276 =  ( n6273 ) ^ ( n6275 )  ;
assign n6277 =  ( n5713 ) | ( n5722 )  ;
assign n6278 =  ( n6277 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6279 =  ( n6276 ) ^ ( n6278 )  ;
assign n6280 = ~ ( n6279 ) ;
assign n6281 =  ( n6265 ) | ( n6280 )  ;
assign n6282 = ~ ( n6281 ) ;
assign n6283 =  ( n6264 ) ^ ( n5894 )  ;
assign n6284 = ~ ( n5902 ) ;
assign n6285 = ~ ( n5913 ) ;
assign n6286 =  ( n6284 ) | ( n6285 )  ;
assign n6287 =  ( n6283 ) ^ ( n6286 )  ;
assign n6288 =  ( n5832 ) | ( n5841 )  ;
assign n6289 =  ( n6288 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6290 = ~ ( n6289 ) ;
assign n6291 =  ( n6287 ) ^ ( n6290 )  ;
assign n6292 =  ( n5682 ) | ( n5691 )  ;
assign n6293 =  ( n6292 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6294 =  ( n6291 ) ^ ( n6293 )  ;
assign n6295 =  ( n5713 ) | ( n5722 )  ;
assign n6296 =  ( n6295 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6297 =  ( n6294 ) ^ ( n6296 )  ;
assign n6298 = ~ ( n6297 ) ;
assign n6299 =  ( bv_1_1_n5 ) ^ ( n6216 )  ;
assign n6300 =  ( n6299 ) ^ ( n6242 )  ;
assign n6301 = ~ ( n5855 ) ;
assign n6302 = ~ ( n5867 ) ;
assign n6303 =  ( n6301 ) | ( n6302 )  ;
assign n6304 =  ( n6300 ) ^ ( n6303 )  ;
assign n6305 =  ( n5832 ) | ( n5841 )  ;
assign n6306 =  ( n6305 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6307 =  ( n6304 ) ^ ( n6306 )  ;
assign n6308 =  ( n5682 ) | ( n5691 )  ;
assign n6309 =  ( n6308 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6310 =  ( n6307 ) ^ ( n6309 )  ;
assign n6311 =  ( n5713 ) | ( n5722 )  ;
assign n6312 =  ( n6311 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6313 =  ( n6310 ) ^ ( n6312 )  ;
assign n6314 = ~ ( n6313 ) ;
assign n6315 =  ( n6298 ) | ( n6314 )  ;
assign n6316 =  ( n6030 ) | ( n6039 )  ;
assign n6317 =  ( n6316 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6318 = ~ ( n6317 ) ;
assign n6319 =  ( n5802 ) | ( n5811 )  ;
assign n6320 =  ( n6319 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6321 = ~ ( n6320 ) ;
assign n6322 =  ( n6318 ) | ( n6321 )  ;
assign n6323 =  ( n5832 ) | ( n5841 )  ;
assign n6324 =  ( n6323 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6325 = ~ ( n6324 ) ;
assign n6326 =  ( n6322 ) | ( n6325 )  ;
assign n6327 =  ( n5682 ) | ( n5691 )  ;
assign n6328 =  ( n6327 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6329 = ~ ( n6328 ) ;
assign n6330 =  ( n6326 ) | ( n6329 )  ;
assign n6331 = ~ ( n6330 ) ;
assign n6332 =  ( n6030 ) | ( n6039 )  ;
assign n6333 =  ( n6332 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6334 =  ( n5802 ) | ( n5811 )  ;
assign n6335 =  ( n6334 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6336 =  ( n6333 ) ^ ( n6335 )  ;
assign n6337 = ~ ( n6336 ) ;
assign n6338 =  ( n6337 ) | ( n5909 )  ;
assign n6339 = ~ ( n6338 ) ;
assign n6340 =  ( n6331 ) | ( n6339 )  ;
assign n6341 =  ( n6030 ) | ( n6039 )  ;
assign n6342 =  ( n6341 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6343 =  ( n5802 ) | ( n5811 )  ;
assign n6344 =  ( n6343 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6345 =  ( n6342 ) ^ ( n6344 )  ;
assign n6346 =  ( n5832 ) | ( n5841 )  ;
assign n6347 =  ( n6346 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6348 =  ( n6345 ) ^ ( n6347 )  ;
assign n6349 =  ( n5682 ) | ( n5691 )  ;
assign n6350 =  ( n6349 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6351 =  ( n6348 ) ^ ( n6350 )  ;
assign n6352 = ~ ( n6351 ) ;
assign n6353 =  ( n5713 ) | ( n5722 )  ;
assign n6354 =  ( n6353 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6355 = ~ ( n6354 ) ;
assign n6356 =  ( n6352 ) | ( n6355 )  ;
assign n6357 = ~ ( n6356 ) ;
assign n6358 =  ( n6340 ) | ( n6357 )  ;
assign n6359 = ~ ( n6358 ) ;
assign n6360 =  ( n6030 ) | ( n6039 )  ;
assign n6361 =  ( n6360 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6362 = ~ ( n6361 ) ;
assign n6363 =  ( n5802 ) | ( n5811 )  ;
assign n6364 =  ( n6363 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6365 = ~ ( n6364 ) ;
assign n6366 =  ( n6362 ) | ( n6365 )  ;
assign n6367 = ~ ( n6366 ) ;
assign n6368 = ~ ( n5902 ) ;
assign n6369 =  ( n6367 ) | ( n6368 )  ;
assign n6370 = ~ ( n6369 ) ;
assign n6371 =  ( n6359 ) | ( n6370 )  ;
assign n6372 = ~ ( n6371 ) ;
assign n6373 = ~ ( n6330 ) ;
assign n6374 =  ( n6337 ) | ( n5909 )  ;
assign n6375 = ~ ( n6374 ) ;
assign n6376 =  ( n6373 ) | ( n6375 )  ;
assign n6377 = ~ ( n6356 ) ;
assign n6378 =  ( n6376 ) | ( n6377 )  ;
assign n6379 = ~ ( n6366 ) ;
assign n6380 = ~ ( n5902 ) ;
assign n6381 =  ( n6379 ) | ( n6380 )  ;
assign n6382 =  ( n6378 ) ^ ( n6381 )  ;
assign n6383 = ~ ( n6382 ) ;
assign n6384 =  ( n6030 ) | ( n6039 )  ;
assign n6385 =  ( n6384 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6386 = ~ ( n6385 ) ;
assign n6387 =  ( n5802 ) | ( n5811 )  ;
assign n6388 =  ( n6387 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6389 =  ( n6386 ) ^ ( n6388 )  ;
assign n6390 =  ( n5832 ) | ( n5841 )  ;
assign n6391 =  ( n6390 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6392 =  ( n6389 ) ^ ( n6391 )  ;
assign n6393 =  ( n5682 ) | ( n5691 )  ;
assign n6394 =  ( n6393 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6395 =  ( n6392 ) ^ ( n6394 )  ;
assign n6396 =  ( n5713 ) | ( n5722 )  ;
assign n6397 =  ( n6396 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6398 =  ( n6395 ) ^ ( n6397 )  ;
assign n6399 = ~ ( n6398 ) ;
assign n6400 =  ( n6383 ) | ( n6399 )  ;
assign n6401 = ~ ( n6400 ) ;
assign n6402 =  ( n6372 ) | ( n6401 )  ;
assign n6403 = ~ ( n6402 ) ;
assign n6404 =  ( bv_1_1_n5 ) ^ ( n6093 )  ;
assign n6405 = ~ ( n6100 ) ;
assign n6406 = ~ ( n5902 ) ;
assign n6407 =  ( n6405 ) | ( n6406 )  ;
assign n6408 =  ( n6404 ) ^ ( n6407 )  ;
assign n6409 =  ( n5802 ) | ( n5811 )  ;
assign n6410 =  ( n6409 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6411 =  ( n6408 ) ^ ( n6410 )  ;
assign n6412 =  ( n5832 ) | ( n5841 )  ;
assign n6413 =  ( n6412 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6414 =  ( n6411 ) ^ ( n6413 )  ;
assign n6415 =  ( n5682 ) | ( n5691 )  ;
assign n6416 =  ( n6415 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6417 =  ( n6414 ) ^ ( n6416 )  ;
assign n6418 =  ( n5713 ) | ( n5722 )  ;
assign n6419 =  ( n6418 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6420 =  ( n6417 ) ^ ( n6419 )  ;
assign n6421 = ~ ( n6420 ) ;
assign n6422 =  ( n6403 ) | ( n6421 )  ;
assign n6423 = ~ ( n6105 ) ;
assign n6424 =  ( n6111 ) | ( n6124 )  ;
assign n6425 = ~ ( n6424 ) ;
assign n6426 =  ( n6423 ) | ( n6425 )  ;
assign n6427 =  ( n6426 ) ^ ( n6166 )  ;
assign n6428 = ~ ( n6173 ) ;
assign n6429 = ~ ( n5736 ) ;
assign n6430 =  ( n6428 ) | ( n6429 )  ;
assign n6431 =  ( n6427 ) ^ ( n6430 )  ;
assign n6432 =  ( n5802 ) | ( n5811 )  ;
assign n6433 =  ( n6432 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6434 = ~ ( n6433 ) ;
assign n6435 =  ( n6431 ) ^ ( n6434 )  ;
assign n6436 =  ( n5832 ) | ( n5841 )  ;
assign n6437 =  ( n6436 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6438 =  ( n6435 ) ^ ( n6437 )  ;
assign n6439 =  ( n5682 ) | ( n5691 )  ;
assign n6440 =  ( n6439 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6441 =  ( n6438 ) ^ ( n6440 )  ;
assign n6442 =  ( n5713 ) | ( n5722 )  ;
assign n6443 =  ( n6442 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6444 =  ( n6441 ) ^ ( n6443 )  ;
assign n6445 = ~ ( n6444 ) ;
assign n6446 =  ( n6422 ) | ( n6445 )  ;
assign n6447 = ~ ( n6446 ) ;
assign n6448 = ~ ( n6402 ) ;
assign n6449 =  ( n6448 ) | ( n6421 )  ;
assign n6450 = ~ ( n6449 ) ;
assign n6451 = ~ ( n6105 ) ;
assign n6452 =  ( n6111 ) | ( n6124 )  ;
assign n6453 = ~ ( n6452 ) ;
assign n6454 =  ( n6451 ) | ( n6453 )  ;
assign n6455 =  ( n6450 ) ^ ( n6454 )  ;
assign n6456 =  ( n6455 ) ^ ( n6166 )  ;
assign n6457 = ~ ( n6173 ) ;
assign n6458 = ~ ( n5736 ) ;
assign n6459 =  ( n6457 ) | ( n6458 )  ;
assign n6460 =  ( n6456 ) ^ ( n6459 )  ;
assign n6461 =  ( n5802 ) | ( n5811 )  ;
assign n6462 =  ( n6461 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6463 = ~ ( n6462 ) ;
assign n6464 =  ( n6460 ) ^ ( n6463 )  ;
assign n6465 =  ( n5832 ) | ( n5841 )  ;
assign n6466 =  ( n6465 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6467 =  ( n6464 ) ^ ( n6466 )  ;
assign n6468 =  ( n5682 ) | ( n5691 )  ;
assign n6469 =  ( n6468 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6470 =  ( n6467 ) ^ ( n6469 )  ;
assign n6471 =  ( n5713 ) | ( n5722 )  ;
assign n6472 =  ( n6471 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6473 =  ( n6470 ) ^ ( n6472 )  ;
assign n6474 = ~ ( n6473 ) ;
assign n6475 = kd[5:5] ;
assign n6476 =  ( n6475 ) == ( bv_1_0_n2 )  ;
assign n6477 = kd[4:4] ;
assign n6478 =  ( n6477 ) == ( bv_1_0_n2 )  ;
assign n6479 =  ( n6476 ) | ( n6478 )  ;
assign n6480 = kd[3:3] ;
assign n6481 =  ( n6480 ) == ( bv_1_0_n2 )  ;
assign n6482 =  ( n6479 ) | ( n6481 )  ;
assign n6483 = ~ ( n6482 )  ;
assign n6484 = kd[5:5] ;
assign n6485 =  ( n6484 ) == ( bv_1_1_n5 )  ;
assign n6486 = kd[4:4] ;
assign n6487 =  ( n6486 ) == ( bv_1_1_n5 )  ;
assign n6488 =  ( n6485 ) | ( n6487 )  ;
assign n6489 = kd[3:3] ;
assign n6490 =  ( n6489 ) == ( bv_1_1_n5 )  ;
assign n6491 =  ( n6488 ) | ( n6490 )  ;
assign n6492 = ~ ( n6491 )  ;
assign n6493 =  ( n6483 ) | ( n6492 )  ;
assign n6494 = kd[5:5] ;
assign n6495 =  ( n6494 ) == ( bv_1_0_n2 )  ;
assign n6496 = kd[4:4] ;
assign n6497 =  ( n6496 ) == ( bv_1_0_n2 )  ;
assign n6498 = kd[3:3] ;
assign n6499 =  ( n6498 ) == ( bv_1_0_n2 )  ;
assign n6500 =  ( n6497 ) | ( n6499 )  ;
assign n6501 = ~ ( n6500 )  ;
assign n6502 =  ( n6495 ) | ( n6501 )  ;
assign n6503 =  ( n6502 ) ? ( bv_1_0_n2 ) : ( bv_1_1_n5 ) ;
assign n6504 =  ( n6493 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6505 = ~ ( n6504 ) ;
assign n6506 =  ( n6030 ) | ( n6039 )  ;
assign n6507 =  ( n6506 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6508 = ~ ( n6507 ) ;
assign n6509 =  ( n6505 ) | ( n6508 )  ;
assign n6510 =  ( n5802 ) | ( n5811 )  ;
assign n6511 =  ( n6510 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6512 = ~ ( n6511 ) ;
assign n6513 =  ( n6509 ) | ( n6512 )  ;
assign n6514 =  ( n5832 ) | ( n5841 )  ;
assign n6515 =  ( n6514 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6516 = ~ ( n6515 ) ;
assign n6517 =  ( n6513 ) | ( n6516 )  ;
assign n6518 = ~ ( n6517 ) ;
assign n6519 =  ( n6483 ) | ( n6492 )  ;
assign n6520 =  ( n6519 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6521 =  ( n6030 ) | ( n6039 )  ;
assign n6522 =  ( n6521 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6523 =  ( n6520 ) ^ ( n6522 )  ;
assign n6524 = ~ ( n6523 ) ;
assign n6525 =  ( n6524 ) | ( n6150 )  ;
assign n6526 = ~ ( n6525 ) ;
assign n6527 =  ( n6518 ) | ( n6526 )  ;
assign n6528 =  ( n6483 ) | ( n6492 )  ;
assign n6529 =  ( n6528 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6530 =  ( n6030 ) | ( n6039 )  ;
assign n6531 =  ( n6530 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6532 =  ( n6529 ) ^ ( n6531 )  ;
assign n6533 =  ( n5802 ) | ( n5811 )  ;
assign n6534 =  ( n6533 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6535 =  ( n6532 ) ^ ( n6534 )  ;
assign n6536 =  ( n5832 ) | ( n5841 )  ;
assign n6537 =  ( n6536 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6538 =  ( n6535 ) ^ ( n6537 )  ;
assign n6539 = ~ ( n6538 ) ;
assign n6540 =  ( n5682 ) | ( n5691 )  ;
assign n6541 =  ( n6540 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6542 = ~ ( n6541 ) ;
assign n6543 =  ( n6539 ) | ( n6542 )  ;
assign n6544 = ~ ( n6543 ) ;
assign n6545 =  ( n6527 ) | ( n6544 )  ;
assign n6546 = ~ ( n6545 ) ;
assign n6547 =  ( n6483 ) | ( n6492 )  ;
assign n6548 =  ( n6547 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6549 = ~ ( n6548 ) ;
assign n6550 =  ( n6030 ) | ( n6039 )  ;
assign n6551 =  ( n6550 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6552 = ~ ( n6551 ) ;
assign n6553 =  ( n6549 ) | ( n6552 )  ;
assign n6554 = ~ ( n6553 ) ;
assign n6555 = ~ ( n6173 ) ;
assign n6556 =  ( n6554 ) | ( n6555 )  ;
assign n6557 = ~ ( n6556 ) ;
assign n6558 =  ( n6546 ) | ( n6557 )  ;
assign n6559 = ~ ( n6558 ) ;
assign n6560 = ~ ( n6517 ) ;
assign n6561 =  ( n6524 ) | ( n6150 )  ;
assign n6562 = ~ ( n6561 ) ;
assign n6563 =  ( n6560 ) | ( n6562 )  ;
assign n6564 = ~ ( n6543 ) ;
assign n6565 =  ( n6563 ) | ( n6564 )  ;
assign n6566 = ~ ( n6553 ) ;
assign n6567 = ~ ( n6173 ) ;
assign n6568 =  ( n6566 ) | ( n6567 )  ;
assign n6569 =  ( n6565 ) ^ ( n6568 )  ;
assign n6570 = ~ ( n6569 ) ;
assign n6571 =  ( n6483 ) | ( n6492 )  ;
assign n6572 =  ( n6571 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6573 = ~ ( n6572 ) ;
assign n6574 =  ( n6030 ) | ( n6039 )  ;
assign n6575 =  ( n6574 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6576 =  ( n6573 ) ^ ( n6575 )  ;
assign n6577 =  ( n5802 ) | ( n5811 )  ;
assign n6578 =  ( n6577 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6579 =  ( n6576 ) ^ ( n6578 )  ;
assign n6580 =  ( n5832 ) | ( n5841 )  ;
assign n6581 =  ( n6580 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6582 =  ( n6579 ) ^ ( n6581 )  ;
assign n6583 =  ( n5682 ) | ( n5691 )  ;
assign n6584 =  ( n6583 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6585 =  ( n6582 ) ^ ( n6584 )  ;
assign n6586 = ~ ( n6585 ) ;
assign n6587 =  ( n6570 ) | ( n6586 )  ;
assign n6588 = ~ ( n6587 ) ;
assign n6589 =  ( n6559 ) | ( n6588 )  ;
assign n6590 = ~ ( n6589 ) ;
assign n6591 =  ( n6483 ) | ( n6492 )  ;
assign n6592 =  ( n6591 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6593 =  ( n6030 ) | ( n6039 )  ;
assign n6594 =  ( n6593 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6595 = ~ ( n6594 ) ;
assign n6596 =  ( n6592 ) | ( n6595 )  ;
assign n6597 =  ( n5802 ) | ( n5811 )  ;
assign n6598 =  ( n6597 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6599 = ~ ( n6598 ) ;
assign n6600 =  ( n6596 ) | ( n6599 )  ;
assign n6601 =  ( n5832 ) | ( n5841 )  ;
assign n6602 =  ( n6601 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6603 = ~ ( n6602 ) ;
assign n6604 =  ( n6600 ) | ( n6603 )  ;
assign n6605 = ~ ( n6604 ) ;
assign n6606 =  ( n6483 ) | ( n6492 )  ;
assign n6607 =  ( n6606 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6608 = ~ ( n6607 ) ;
assign n6609 =  ( n6030 ) | ( n6039 )  ;
assign n6610 =  ( n6609 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6611 =  ( n6608 ) ^ ( n6610 )  ;
assign n6612 = ~ ( n6611 ) ;
assign n6613 =  ( n6612 ) | ( n6150 )  ;
assign n6614 = ~ ( n6613 ) ;
assign n6615 =  ( n6605 ) | ( n6614 )  ;
assign n6616 =  ( n6483 ) | ( n6492 )  ;
assign n6617 =  ( n6616 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6618 = ~ ( n6617 ) ;
assign n6619 =  ( n6030 ) | ( n6039 )  ;
assign n6620 =  ( n6619 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6621 =  ( n6618 ) ^ ( n6620 )  ;
assign n6622 =  ( n5802 ) | ( n5811 )  ;
assign n6623 =  ( n6622 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6624 =  ( n6621 ) ^ ( n6623 )  ;
assign n6625 =  ( n5832 ) | ( n5841 )  ;
assign n6626 =  ( n6625 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6627 =  ( n6624 ) ^ ( n6626 )  ;
assign n6628 = ~ ( n6627 ) ;
assign n6629 =  ( n5682 ) | ( n5691 )  ;
assign n6630 =  ( n6629 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6631 = ~ ( n6630 ) ;
assign n6632 =  ( n6628 ) | ( n6631 )  ;
assign n6633 = ~ ( n6632 ) ;
assign n6634 =  ( n6615 ) | ( n6633 )  ;
assign n6635 =  ( n6483 ) | ( n6492 )  ;
assign n6636 =  ( n6635 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6637 =  ( n6030 ) | ( n6039 )  ;
assign n6638 =  ( n6637 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6639 = ~ ( n6638 ) ;
assign n6640 =  ( n6636 ) | ( n6639 )  ;
assign n6641 = ~ ( n6640 ) ;
assign n6642 = ~ ( n6173 ) ;
assign n6643 =  ( n6641 ) | ( n6642 )  ;
assign n6644 =  ( n6634 ) ^ ( n6643 )  ;
assign n6645 =  ( n6030 ) | ( n6039 )  ;
assign n6646 =  ( n6645 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6647 =  ( n6644 ) ^ ( n6646 )  ;
assign n6648 =  ( n5802 ) | ( n5811 )  ;
assign n6649 =  ( n6648 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6650 =  ( n6647 ) ^ ( n6649 )  ;
assign n6651 =  ( n5832 ) | ( n5841 )  ;
assign n6652 =  ( n6651 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6653 =  ( n6650 ) ^ ( n6652 )  ;
assign n6654 =  ( n5682 ) | ( n5691 )  ;
assign n6655 =  ( n6654 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6656 =  ( n6653 ) ^ ( n6655 )  ;
assign n6657 =  ( n5713 ) | ( n5722 )  ;
assign n6658 =  ( n6657 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6659 =  ( n6656 ) ^ ( n6658 )  ;
assign n6660 = ~ ( n6659 ) ;
assign n6661 =  ( n6590 ) | ( n6660 )  ;
assign n6662 = ~ ( n6661 ) ;
assign n6663 =  ( n6589 ) ^ ( n6634 )  ;
assign n6664 = ~ ( n6640 ) ;
assign n6665 = ~ ( n6173 ) ;
assign n6666 =  ( n6664 ) | ( n6665 )  ;
assign n6667 =  ( n6663 ) ^ ( n6666 )  ;
assign n6668 =  ( n6030 ) | ( n6039 )  ;
assign n6669 =  ( n6668 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6670 =  ( n6667 ) ^ ( n6669 )  ;
assign n6671 =  ( n5802 ) | ( n5811 )  ;
assign n6672 =  ( n6671 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6673 =  ( n6670 ) ^ ( n6672 )  ;
assign n6674 =  ( n5832 ) | ( n5841 )  ;
assign n6675 =  ( n6674 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6676 =  ( n6673 ) ^ ( n6675 )  ;
assign n6677 =  ( n5682 ) | ( n5691 )  ;
assign n6678 =  ( n6677 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6679 =  ( n6676 ) ^ ( n6678 )  ;
assign n6680 =  ( n5713 ) | ( n5722 )  ;
assign n6681 =  ( n6680 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6682 =  ( n6679 ) ^ ( n6681 )  ;
assign n6683 =  ( n6662 ) | ( n6682 )  ;
assign n6684 = ~ ( n6683 ) ;
assign n6685 = ~ ( n6634 ) ;
assign n6686 = ~ ( n6640 ) ;
assign n6687 = ~ ( n6173 ) ;
assign n6688 =  ( n6686 ) | ( n6687 )  ;
assign n6689 = ~ ( n6688 ) ;
assign n6690 =  ( n6685 ) | ( n6689 )  ;
assign n6691 = ~ ( n6690 ) ;
assign n6692 = ~ ( n6640 ) ;
assign n6693 = ~ ( n6173 ) ;
assign n6694 =  ( n6692 ) | ( n6693 )  ;
assign n6695 =  ( n6634 ) ^ ( n6694 )  ;
assign n6696 = ~ ( n6695 ) ;
assign n6697 =  ( n6030 ) | ( n6039 )  ;
assign n6698 =  ( n6697 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6699 =  ( n5802 ) | ( n5811 )  ;
assign n6700 =  ( n6699 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6701 =  ( n6698 ) ^ ( n6700 )  ;
assign n6702 =  ( n5832 ) | ( n5841 )  ;
assign n6703 =  ( n6702 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6704 =  ( n6701 ) ^ ( n6703 )  ;
assign n6705 =  ( n5682 ) | ( n5691 )  ;
assign n6706 =  ( n6705 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6707 =  ( n6704 ) ^ ( n6706 )  ;
assign n6708 =  ( n5713 ) | ( n5722 )  ;
assign n6709 =  ( n6708 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6710 =  ( n6707 ) ^ ( n6709 )  ;
assign n6711 = ~ ( n6710 ) ;
assign n6712 =  ( n6696 ) | ( n6711 )  ;
assign n6713 = ~ ( n6712 ) ;
assign n6714 =  ( n6691 ) | ( n6713 )  ;
assign n6715 = ~ ( n6714 ) ;
assign n6716 =  ( n6684 ) | ( n6715 )  ;
assign n6717 = ~ ( n6716 ) ;
assign n6718 = ~ ( n6690 ) ;
assign n6719 =  ( n6696 ) | ( n6711 )  ;
assign n6720 = ~ ( n6719 ) ;
assign n6721 =  ( n6718 ) | ( n6720 )  ;
assign n6722 =  ( n6683 ) ^ ( n6721 )  ;
assign n6723 = ~ ( n6722 ) ;
assign n6724 = ~ ( n6330 ) ;
assign n6725 =  ( n6337 ) | ( n5909 )  ;
assign n6726 = ~ ( n6725 ) ;
assign n6727 =  ( n6724 ) | ( n6726 )  ;
assign n6728 = ~ ( n6356 ) ;
assign n6729 =  ( n6727 ) | ( n6728 )  ;
assign n6730 = ~ ( n6366 ) ;
assign n6731 = ~ ( n5902 ) ;
assign n6732 =  ( n6730 ) | ( n6731 )  ;
assign n6733 =  ( n6729 ) ^ ( n6732 )  ;
assign n6734 =  ( n6030 ) | ( n6039 )  ;
assign n6735 =  ( n6734 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6736 = ~ ( n6735 ) ;
assign n6737 =  ( n6733 ) ^ ( n6736 )  ;
assign n6738 =  ( n5802 ) | ( n5811 )  ;
assign n6739 =  ( n6738 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6740 =  ( n6737 ) ^ ( n6739 )  ;
assign n6741 =  ( n5832 ) | ( n5841 )  ;
assign n6742 =  ( n6741 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6743 =  ( n6740 ) ^ ( n6742 )  ;
assign n6744 =  ( n5682 ) | ( n5691 )  ;
assign n6745 =  ( n6744 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6746 =  ( n6743 ) ^ ( n6745 )  ;
assign n6747 =  ( n5713 ) | ( n5722 )  ;
assign n6748 =  ( n6747 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6749 =  ( n6746 ) ^ ( n6748 )  ;
assign n6750 = ~ ( n6749 ) ;
assign n6751 =  ( n6723 ) | ( n6750 )  ;
assign n6752 = ~ ( n6751 ) ;
assign n6753 =  ( n6717 ) | ( n6752 )  ;
assign n6754 = ~ ( n6753 ) ;
assign n6755 =  ( n6474 ) | ( n6754 )  ;
assign n6756 =  ( bv_1_1_n5 ) ^ ( n6402 )  ;
assign n6757 =  ( n6756 ) ^ ( n6093 )  ;
assign n6758 = ~ ( n6100 ) ;
assign n6759 = ~ ( n5902 ) ;
assign n6760 =  ( n6758 ) | ( n6759 )  ;
assign n6761 =  ( n6757 ) ^ ( n6760 )  ;
assign n6762 =  ( n5802 ) | ( n5811 )  ;
assign n6763 =  ( n6762 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6764 =  ( n6761 ) ^ ( n6763 )  ;
assign n6765 =  ( n5832 ) | ( n5841 )  ;
assign n6766 =  ( n6765 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6767 =  ( n6764 ) ^ ( n6766 )  ;
assign n6768 =  ( n5682 ) | ( n5691 )  ;
assign n6769 =  ( n6768 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6770 =  ( n6767 ) ^ ( n6769 )  ;
assign n6771 =  ( n5713 ) | ( n5722 )  ;
assign n6772 =  ( n6771 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6773 =  ( n6770 ) ^ ( n6772 )  ;
assign n6774 = ~ ( n6773 ) ;
assign n6775 =  ( n6755 ) | ( n6774 )  ;
assign n6776 = ~ ( n6775 ) ;
assign n6777 =  ( n6447 ) | ( n6776 )  ;
assign n6778 = ~ ( n6777 ) ;
assign n6779 =  ( n6315 ) | ( n6778 )  ;
assign n6780 = ~ ( n6779 ) ;
assign n6781 =  ( n6282 ) | ( n6780 )  ;
assign n6782 = ~ ( n6781 ) ;
assign n6783 =  ( n6021 ) | ( n6782 )  ;
assign n6784 = ~ ( n6783 ) ;
assign n6785 =  ( n5990 ) | ( n6784 )  ;
assign n6786 = ~ ( n5783 ) ;
assign n6787 =  ( n6786 ) | ( n5792 )  ;
assign n6788 = ~ ( n6006 ) ;
assign n6789 =  ( n6787 ) | ( n6788 )  ;
assign n6790 =  ( n6789 ) | ( n6020 )  ;
assign n6791 = ~ ( n6297 ) ;
assign n6792 =  ( n6790 ) | ( n6791 )  ;
assign n6793 =  ( n6792 ) | ( n6314 )  ;
assign n6794 = ~ ( n6473 ) ;
assign n6795 =  ( n6793 ) | ( n6794 )  ;
assign n6796 =  ( bv_1_1_n5 ) ^ ( n6753 )  ;
assign n6797 =  ( n6796 ) ^ ( n6402 )  ;
assign n6798 =  ( n6797 ) ^ ( n6093 )  ;
assign n6799 = ~ ( n6100 ) ;
assign n6800 = ~ ( n5902 ) ;
assign n6801 =  ( n6799 ) | ( n6800 )  ;
assign n6802 =  ( n6798 ) ^ ( n6801 )  ;
assign n6803 =  ( n5802 ) | ( n5811 )  ;
assign n6804 =  ( n6803 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6805 =  ( n6802 ) ^ ( n6804 )  ;
assign n6806 =  ( n5832 ) | ( n5841 )  ;
assign n6807 =  ( n6806 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6808 =  ( n6805 ) ^ ( n6807 )  ;
assign n6809 =  ( n5682 ) | ( n5691 )  ;
assign n6810 =  ( n6809 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6811 =  ( n6808 ) ^ ( n6810 )  ;
assign n6812 =  ( n5713 ) | ( n5722 )  ;
assign n6813 =  ( n6812 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6814 =  ( n6811 ) ^ ( n6813 )  ;
assign n6815 = ~ ( n6814 ) ;
assign n6816 =  ( n6795 ) | ( n6815 )  ;
assign n6817 = kd[3:3] ;
assign n6818 =  ( n6817 ) == ( bv_1_0_n2 )  ;
assign n6819 = kd[2:2] ;
assign n6820 =  ( n6819 ) == ( bv_1_0_n2 )  ;
assign n6821 =  ( n6818 ) | ( n6820 )  ;
assign n6822 = kd[1:1] ;
assign n6823 =  ( n6822 ) == ( bv_1_0_n2 )  ;
assign n6824 =  ( n6821 ) | ( n6823 )  ;
assign n6825 = ~ ( n6824 )  ;
assign n6826 = kd[3:3] ;
assign n6827 =  ( n6826 ) == ( bv_1_1_n5 )  ;
assign n6828 = kd[2:2] ;
assign n6829 =  ( n6828 ) == ( bv_1_1_n5 )  ;
assign n6830 =  ( n6827 ) | ( n6829 )  ;
assign n6831 = kd[1:1] ;
assign n6832 =  ( n6831 ) == ( bv_1_1_n5 )  ;
assign n6833 =  ( n6830 ) | ( n6832 )  ;
assign n6834 = ~ ( n6833 )  ;
assign n6835 =  ( n6825 ) | ( n6834 )  ;
assign n6836 = kd[3:3] ;
assign n6837 =  ( n6836 ) == ( bv_1_0_n2 )  ;
assign n6838 = kd[2:2] ;
assign n6839 =  ( n6838 ) == ( bv_1_0_n2 )  ;
assign n6840 = kd[1:1] ;
assign n6841 =  ( n6840 ) == ( bv_1_0_n2 )  ;
assign n6842 =  ( n6839 ) | ( n6841 )  ;
assign n6843 = ~ ( n6842 )  ;
assign n6844 =  ( n6837 ) | ( n6843 )  ;
assign n6845 =  ( n6844 ) ? ( bv_1_0_n2 ) : ( bv_1_1_n5 ) ;
assign n6846 =  ( n6835 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n6847 =  ( n6483 ) | ( n6492 )  ;
assign n6848 =  ( n6847 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6849 = ~ ( n6848 ) ;
assign n6850 =  ( n6846 ) | ( n6849 )  ;
assign n6851 =  ( n6030 ) | ( n6039 )  ;
assign n6852 =  ( n6851 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6853 = ~ ( n6852 ) ;
assign n6854 =  ( n6850 ) | ( n6853 )  ;
assign n6855 =  ( n5802 ) | ( n5811 )  ;
assign n6856 =  ( n6855 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6857 = ~ ( n6856 ) ;
assign n6858 =  ( n6854 ) | ( n6857 )  ;
assign n6859 = ~ ( n6858 ) ;
assign n6860 =  ( n6825 ) | ( n6834 )  ;
assign n6861 =  ( n6860 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n6862 = ~ ( n6861 ) ;
assign n6863 =  ( n6483 ) | ( n6492 )  ;
assign n6864 =  ( n6863 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6865 =  ( n6862 ) ^ ( n6864 )  ;
assign n6866 = ~ ( n6865 ) ;
assign n6867 =  ( n6866 ) | ( n6337 )  ;
assign n6868 = ~ ( n6867 ) ;
assign n6869 =  ( n6859 ) | ( n6868 )  ;
assign n6870 =  ( n6825 ) | ( n6834 )  ;
assign n6871 =  ( n6870 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n6872 = ~ ( n6871 ) ;
assign n6873 =  ( n6483 ) | ( n6492 )  ;
assign n6874 =  ( n6873 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6875 =  ( n6872 ) ^ ( n6874 )  ;
assign n6876 =  ( n6030 ) | ( n6039 )  ;
assign n6877 =  ( n6876 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6878 =  ( n6875 ) ^ ( n6877 )  ;
assign n6879 =  ( n5802 ) | ( n5811 )  ;
assign n6880 =  ( n6879 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6881 =  ( n6878 ) ^ ( n6880 )  ;
assign n6882 = ~ ( n6881 ) ;
assign n6883 =  ( n5832 ) | ( n5841 )  ;
assign n6884 =  ( n6883 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6885 = ~ ( n6884 ) ;
assign n6886 =  ( n6882 ) | ( n6885 )  ;
assign n6887 = ~ ( n6886 ) ;
assign n6888 =  ( n6869 ) | ( n6887 )  ;
assign n6889 = ~ ( n6888 ) ;
assign n6890 =  ( n6825 ) | ( n6834 )  ;
assign n6891 =  ( n6890 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n6892 =  ( n6483 ) | ( n6492 )  ;
assign n6893 =  ( n6892 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6894 = ~ ( n6893 ) ;
assign n6895 =  ( n6891 ) | ( n6894 )  ;
assign n6896 = ~ ( n6895 ) ;
assign n6897 = ~ ( n6366 ) ;
assign n6898 =  ( n6896 ) | ( n6897 )  ;
assign n6899 = ~ ( n6898 ) ;
assign n6900 =  ( n6889 ) | ( n6899 )  ;
assign n6901 =  ( n6483 ) | ( n6492 )  ;
assign n6902 =  ( n6901 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6903 =  ( n6030 ) | ( n6039 )  ;
assign n6904 =  ( n6903 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6905 =  ( n6902 ) ^ ( n6904 )  ;
assign n6906 =  ( n5802 ) | ( n5811 )  ;
assign n6907 =  ( n6906 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6908 =  ( n6905 ) ^ ( n6907 )  ;
assign n6909 =  ( n5832 ) | ( n5841 )  ;
assign n6910 =  ( n6909 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6911 =  ( n6908 ) ^ ( n6910 )  ;
assign n6912 =  ( n5682 ) | ( n5691 )  ;
assign n6913 =  ( n6912 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6914 =  ( n6911 ) ^ ( n6913 )  ;
assign n6915 = ~ ( n6914 ) ;
assign n6916 =  ( n6900 ) | ( n6915 )  ;
assign n6917 =  ( n5713 ) | ( n5722 )  ;
assign n6918 =  ( n6917 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6919 = ~ ( n6918 ) ;
assign n6920 =  ( n6916 ) | ( n6919 )  ;
assign n6921 = ~ ( n6920 ) ;
assign n6922 = ~ ( n6895 ) ;
assign n6923 = ~ ( n6366 ) ;
assign n6924 =  ( n6922 ) | ( n6923 )  ;
assign n6925 =  ( n6888 ) ^ ( n6924 )  ;
assign n6926 = ~ ( n6925 ) ;
assign n6927 =  ( n6483 ) | ( n6492 )  ;
assign n6928 =  ( n6927 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6929 =  ( n6030 ) | ( n6039 )  ;
assign n6930 =  ( n6929 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6931 =  ( n6928 ) ^ ( n6930 )  ;
assign n6932 =  ( n5802 ) | ( n5811 )  ;
assign n6933 =  ( n6932 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6934 =  ( n6931 ) ^ ( n6933 )  ;
assign n6935 =  ( n5832 ) | ( n5841 )  ;
assign n6936 =  ( n6935 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6937 =  ( n6934 ) ^ ( n6936 )  ;
assign n6938 =  ( n5682 ) | ( n5691 )  ;
assign n6939 =  ( n6938 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6940 =  ( n6937 ) ^ ( n6939 )  ;
assign n6941 =  ( n5713 ) | ( n5722 )  ;
assign n6942 =  ( n6941 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6943 =  ( n6940 ) ^ ( n6942 )  ;
assign n6944 = ~ ( n6943 ) ;
assign n6945 =  ( n6926 ) | ( n6944 )  ;
assign n6946 = ~ ( n6945 ) ;
assign n6947 =  ( n6921 ) | ( n6946 )  ;
assign n6948 = ~ ( n6895 ) ;
assign n6949 = ~ ( n6366 ) ;
assign n6950 =  ( n6948 ) | ( n6949 )  ;
assign n6951 =  ( n6888 ) ^ ( n6950 )  ;
assign n6952 =  ( n6483 ) | ( n6492 )  ;
assign n6953 =  ( n6952 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n6954 =  ( n6951 ) ^ ( n6953 )  ;
assign n6955 =  ( n6030 ) | ( n6039 )  ;
assign n6956 =  ( n6955 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n6957 =  ( n6954 ) ^ ( n6956 )  ;
assign n6958 =  ( n5802 ) | ( n5811 )  ;
assign n6959 =  ( n6958 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n6960 =  ( n6957 ) ^ ( n6959 )  ;
assign n6961 =  ( n5832 ) | ( n5841 )  ;
assign n6962 =  ( n6961 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n6963 =  ( n6960 ) ^ ( n6962 )  ;
assign n6964 =  ( n5682 ) | ( n5691 )  ;
assign n6965 =  ( n6964 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n6966 =  ( n6963 ) ^ ( n6965 )  ;
assign n6967 =  ( n5713 ) | ( n5722 )  ;
assign n6968 =  ( n6967 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6969 =  ( n6966 ) ^ ( n6968 )  ;
assign n6970 =  ( n6947 ) | ( n6969 )  ;
assign n6971 = ~ ( n6970 ) ;
assign n6972 = ~ ( n6888 ) ;
assign n6973 = ~ ( n6895 ) ;
assign n6974 = ~ ( n6366 ) ;
assign n6975 =  ( n6973 ) | ( n6974 )  ;
assign n6976 = ~ ( n6975 ) ;
assign n6977 =  ( n6972 ) | ( n6976 )  ;
assign n6978 = ~ ( n6977 ) ;
assign n6979 =  ( n5713 ) | ( n5722 )  ;
assign n6980 =  ( n6979 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n6981 = ~ ( n6980 ) ;
assign n6982 =  ( n6915 ) | ( n6981 )  ;
assign n6983 = ~ ( n6982 ) ;
assign n6984 =  ( n6978 ) | ( n6983 )  ;
assign n6985 = ~ ( n6984 ) ;
assign n6986 =  ( n6971 ) | ( n6985 )  ;
assign n6987 = ~ ( n6986 ) ;
assign n6988 = ~ ( n6977 ) ;
assign n6989 = ~ ( n6982 ) ;
assign n6990 =  ( n6988 ) | ( n6989 )  ;
assign n6991 =  ( n6970 ) ^ ( n6990 )  ;
assign n6992 = ~ ( n6991 ) ;
assign n6993 = ~ ( n6517 ) ;
assign n6994 =  ( n6524 ) | ( n6150 )  ;
assign n6995 = ~ ( n6994 ) ;
assign n6996 =  ( n6993 ) | ( n6995 )  ;
assign n6997 = ~ ( n6543 ) ;
assign n6998 =  ( n6996 ) | ( n6997 )  ;
assign n6999 = ~ ( n6553 ) ;
assign n7000 = ~ ( n6173 ) ;
assign n7001 =  ( n6999 ) | ( n7000 )  ;
assign n7002 =  ( n6998 ) ^ ( n7001 )  ;
assign n7003 =  ( n6483 ) | ( n6492 )  ;
assign n7004 =  ( n7003 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7005 = ~ ( n7004 ) ;
assign n7006 =  ( n7002 ) ^ ( n7005 )  ;
assign n7007 =  ( n6030 ) | ( n6039 )  ;
assign n7008 =  ( n7007 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7009 =  ( n7006 ) ^ ( n7008 )  ;
assign n7010 =  ( n5802 ) | ( n5811 )  ;
assign n7011 =  ( n7010 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7012 =  ( n7009 ) ^ ( n7011 )  ;
assign n7013 =  ( n5832 ) | ( n5841 )  ;
assign n7014 =  ( n7013 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7015 =  ( n7012 ) ^ ( n7014 )  ;
assign n7016 =  ( n5682 ) | ( n5691 )  ;
assign n7017 =  ( n7016 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7018 =  ( n7015 ) ^ ( n7017 )  ;
assign n7019 = ~ ( n7018 ) ;
assign n7020 =  ( n6992 ) | ( n7019 )  ;
assign n7021 = ~ ( n7020 ) ;
assign n7022 =  ( n6987 ) | ( n7021 )  ;
assign n7023 = ~ ( n7022 ) ;
assign n7024 =  ( bv_1_1_n5 ) ^ ( n6589 )  ;
assign n7025 =  ( n7024 ) ^ ( n6634 )  ;
assign n7026 = ~ ( n6640 ) ;
assign n7027 = ~ ( n6173 ) ;
assign n7028 =  ( n7026 ) | ( n7027 )  ;
assign n7029 =  ( n7025 ) ^ ( n7028 )  ;
assign n7030 =  ( n6030 ) | ( n6039 )  ;
assign n7031 =  ( n7030 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7032 =  ( n7029 ) ^ ( n7031 )  ;
assign n7033 =  ( n5802 ) | ( n5811 )  ;
assign n7034 =  ( n7033 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7035 =  ( n7032 ) ^ ( n7034 )  ;
assign n7036 =  ( n5832 ) | ( n5841 )  ;
assign n7037 =  ( n7036 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7038 =  ( n7035 ) ^ ( n7037 )  ;
assign n7039 =  ( n5682 ) | ( n5691 )  ;
assign n7040 =  ( n7039 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7041 =  ( n7038 ) ^ ( n7040 )  ;
assign n7042 =  ( n5713 ) | ( n5722 )  ;
assign n7043 =  ( n7042 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7044 =  ( n7041 ) ^ ( n7043 )  ;
assign n7045 = ~ ( n7044 ) ;
assign n7046 =  ( n7023 ) | ( n7045 )  ;
assign n7047 = ~ ( n6690 ) ;
assign n7048 =  ( n6696 ) | ( n6711 )  ;
assign n7049 = ~ ( n7048 ) ;
assign n7050 =  ( n7047 ) | ( n7049 )  ;
assign n7051 =  ( n6683 ) ^ ( n7050 )  ;
assign n7052 = ~ ( n6330 ) ;
assign n7053 =  ( n6337 ) | ( n5909 )  ;
assign n7054 = ~ ( n7053 ) ;
assign n7055 =  ( n7052 ) | ( n7054 )  ;
assign n7056 = ~ ( n6356 ) ;
assign n7057 =  ( n7055 ) | ( n7056 )  ;
assign n7058 =  ( n7051 ) ^ ( n7057 )  ;
assign n7059 = ~ ( n6366 ) ;
assign n7060 = ~ ( n5902 ) ;
assign n7061 =  ( n7059 ) | ( n7060 )  ;
assign n7062 =  ( n7058 ) ^ ( n7061 )  ;
assign n7063 =  ( n6030 ) | ( n6039 )  ;
assign n7064 =  ( n7063 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7065 = ~ ( n7064 ) ;
assign n7066 =  ( n7062 ) ^ ( n7065 )  ;
assign n7067 =  ( n5802 ) | ( n5811 )  ;
assign n7068 =  ( n7067 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7069 =  ( n7066 ) ^ ( n7068 )  ;
assign n7070 =  ( n5832 ) | ( n5841 )  ;
assign n7071 =  ( n7070 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7072 =  ( n7069 ) ^ ( n7071 )  ;
assign n7073 =  ( n5682 ) | ( n5691 )  ;
assign n7074 =  ( n7073 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7075 =  ( n7072 ) ^ ( n7074 )  ;
assign n7076 =  ( n5713 ) | ( n5722 )  ;
assign n7077 =  ( n7076 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7078 =  ( n7075 ) ^ ( n7077 )  ;
assign n7079 = ~ ( n7078 ) ;
assign n7080 =  ( n7046 ) | ( n7079 )  ;
assign n7081 = ~ ( n7080 ) ;
assign n7082 = ~ ( n7022 ) ;
assign n7083 =  ( n7082 ) | ( n7045 )  ;
assign n7084 = ~ ( n7083 ) ;
assign n7085 =  ( n7084 ) ^ ( n6683 )  ;
assign n7086 = ~ ( n6690 ) ;
assign n7087 =  ( n6696 ) | ( n6711 )  ;
assign n7088 = ~ ( n7087 ) ;
assign n7089 =  ( n7086 ) | ( n7088 )  ;
assign n7090 =  ( n7085 ) ^ ( n7089 )  ;
assign n7091 = ~ ( n6330 ) ;
assign n7092 =  ( n6337 ) | ( n5909 )  ;
assign n7093 = ~ ( n7092 ) ;
assign n7094 =  ( n7091 ) | ( n7093 )  ;
assign n7095 = ~ ( n6356 ) ;
assign n7096 =  ( n7094 ) | ( n7095 )  ;
assign n7097 =  ( n7090 ) ^ ( n7096 )  ;
assign n7098 = ~ ( n6366 ) ;
assign n7099 = ~ ( n5902 ) ;
assign n7100 =  ( n7098 ) | ( n7099 )  ;
assign n7101 =  ( n7097 ) ^ ( n7100 )  ;
assign n7102 =  ( n6030 ) | ( n6039 )  ;
assign n7103 =  ( n7102 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7104 = ~ ( n7103 ) ;
assign n7105 =  ( n7101 ) ^ ( n7104 )  ;
assign n7106 =  ( n5802 ) | ( n5811 )  ;
assign n7107 =  ( n7106 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7108 =  ( n7105 ) ^ ( n7107 )  ;
assign n7109 =  ( n5832 ) | ( n5841 )  ;
assign n7110 =  ( n7109 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7111 =  ( n7108 ) ^ ( n7110 )  ;
assign n7112 =  ( n5682 ) | ( n5691 )  ;
assign n7113 =  ( n7112 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7114 =  ( n7111 ) ^ ( n7113 )  ;
assign n7115 =  ( n5713 ) | ( n5722 )  ;
assign n7116 =  ( n7115 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7117 =  ( n7114 ) ^ ( n7116 )  ;
assign n7118 = ~ ( n7117 ) ;
assign n7119 =  ( n6825 ) | ( n6834 )  ;
assign n7120 =  ( n7119 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7121 = ~ ( n7120 ) ;
assign n7122 =  ( n6483 ) | ( n6492 )  ;
assign n7123 =  ( n7122 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7124 = ~ ( n7123 ) ;
assign n7125 =  ( n7121 ) | ( n7124 )  ;
assign n7126 =  ( n6030 ) | ( n6039 )  ;
assign n7127 =  ( n7126 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7128 = ~ ( n7127 ) ;
assign n7129 =  ( n7125 ) | ( n7128 )  ;
assign n7130 =  ( n5802 ) | ( n5811 )  ;
assign n7131 =  ( n7130 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7132 = ~ ( n7131 ) ;
assign n7133 =  ( n7129 ) | ( n7132 )  ;
assign n7134 = ~ ( n7133 ) ;
assign n7135 =  ( n6825 ) | ( n6834 )  ;
assign n7136 =  ( n7135 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7137 =  ( n6483 ) | ( n6492 )  ;
assign n7138 =  ( n7137 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7139 =  ( n7136 ) ^ ( n7138 )  ;
assign n7140 = ~ ( n7139 ) ;
assign n7141 =  ( n7140 ) | ( n6337 )  ;
assign n7142 = ~ ( n7141 ) ;
assign n7143 =  ( n7134 ) | ( n7142 )  ;
assign n7144 =  ( n6825 ) | ( n6834 )  ;
assign n7145 =  ( n7144 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7146 =  ( n6483 ) | ( n6492 )  ;
assign n7147 =  ( n7146 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7148 =  ( n7145 ) ^ ( n7147 )  ;
assign n7149 =  ( n6030 ) | ( n6039 )  ;
assign n7150 =  ( n7149 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7151 =  ( n7148 ) ^ ( n7150 )  ;
assign n7152 =  ( n5802 ) | ( n5811 )  ;
assign n7153 =  ( n7152 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7154 =  ( n7151 ) ^ ( n7153 )  ;
assign n7155 = ~ ( n7154 ) ;
assign n7156 =  ( n5832 ) | ( n5841 )  ;
assign n7157 =  ( n7156 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7158 = ~ ( n7157 ) ;
assign n7159 =  ( n7155 ) | ( n7158 )  ;
assign n7160 = ~ ( n7159 ) ;
assign n7161 =  ( n7143 ) | ( n7160 )  ;
assign n7162 = ~ ( n7161 ) ;
assign n7163 =  ( n6825 ) | ( n6834 )  ;
assign n7164 =  ( n7163 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7165 = ~ ( n7164 ) ;
assign n7166 =  ( n6483 ) | ( n6492 )  ;
assign n7167 =  ( n7166 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7168 = ~ ( n7167 ) ;
assign n7169 =  ( n7165 ) | ( n7168 )  ;
assign n7170 = ~ ( n7169 ) ;
assign n7171 = ~ ( n6366 ) ;
assign n7172 =  ( n7170 ) | ( n7171 )  ;
assign n7173 = ~ ( n7172 ) ;
assign n7174 =  ( n7162 ) | ( n7173 )  ;
assign n7175 = ~ ( n5736 ) ;
assign n7176 =  ( n7175 ) | ( n5742 )  ;
assign n7177 = ~ ( n7176 ) ;
assign n7178 =  ( n7174 ) | ( n7177 )  ;
assign n7179 =  ( n6825 ) | ( n6834 )  ;
assign n7180 =  ( n7179 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7181 = ~ ( n7180 ) ;
assign n7182 =  ( n6483 ) | ( n6492 )  ;
assign n7183 =  ( n7182 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7184 =  ( n7181 ) ^ ( n7183 )  ;
assign n7185 =  ( n6030 ) | ( n6039 )  ;
assign n7186 =  ( n7185 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7187 =  ( n7184 ) ^ ( n7186 )  ;
assign n7188 =  ( n5802 ) | ( n5811 )  ;
assign n7189 =  ( n7188 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7190 =  ( n7187 ) ^ ( n7189 )  ;
assign n7191 =  ( n5832 ) | ( n5841 )  ;
assign n7192 =  ( n7191 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7193 =  ( n7190 ) ^ ( n7192 )  ;
assign n7194 = ~ ( n7193 ) ;
assign n7195 =  ( n7178 ) | ( n7194 )  ;
assign n7196 = ~ ( n7195 ) ;
assign n7197 = ~ ( n7133 ) ;
assign n7198 =  ( n7140 ) | ( n6337 )  ;
assign n7199 = ~ ( n7198 ) ;
assign n7200 =  ( n7197 ) | ( n7199 )  ;
assign n7201 = ~ ( n7159 ) ;
assign n7202 =  ( n7200 ) | ( n7201 )  ;
assign n7203 = ~ ( n7169 ) ;
assign n7204 = ~ ( n6366 ) ;
assign n7205 =  ( n7203 ) | ( n7204 )  ;
assign n7206 =  ( n7202 ) ^ ( n7205 )  ;
assign n7207 = ~ ( n7206 ) ;
assign n7208 = ~ ( n5736 ) ;
assign n7209 =  ( n7208 ) | ( n5742 )  ;
assign n7210 =  ( n6825 ) | ( n6834 )  ;
assign n7211 =  ( n7210 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7212 = ~ ( n7211 ) ;
assign n7213 =  ( n7209 ) ^ ( n7212 )  ;
assign n7214 =  ( n6483 ) | ( n6492 )  ;
assign n7215 =  ( n7214 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7216 =  ( n7213 ) ^ ( n7215 )  ;
assign n7217 =  ( n6030 ) | ( n6039 )  ;
assign n7218 =  ( n7217 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7219 =  ( n7216 ) ^ ( n7218 )  ;
assign n7220 =  ( n5802 ) | ( n5811 )  ;
assign n7221 =  ( n7220 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7222 =  ( n7219 ) ^ ( n7221 )  ;
assign n7223 =  ( n5832 ) | ( n5841 )  ;
assign n7224 =  ( n7223 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7225 =  ( n7222 ) ^ ( n7224 )  ;
assign n7226 = ~ ( n7225 ) ;
assign n7227 =  ( n7207 ) | ( n7226 )  ;
assign n7228 = ~ ( n7227 ) ;
assign n7229 =  ( n7196 ) | ( n7228 )  ;
assign n7230 = ~ ( n7133 ) ;
assign n7231 =  ( n7140 ) | ( n6337 )  ;
assign n7232 = ~ ( n7231 ) ;
assign n7233 =  ( n7230 ) | ( n7232 )  ;
assign n7234 = ~ ( n7159 ) ;
assign n7235 =  ( n7233 ) | ( n7234 )  ;
assign n7236 = ~ ( n7169 ) ;
assign n7237 = ~ ( n6366 ) ;
assign n7238 =  ( n7236 ) | ( n7237 )  ;
assign n7239 =  ( n7235 ) ^ ( n7238 )  ;
assign n7240 = ~ ( n5736 ) ;
assign n7241 =  ( n7240 ) | ( n5742 )  ;
assign n7242 =  ( n7239 ) ^ ( n7241 )  ;
assign n7243 =  ( n6825 ) | ( n6834 )  ;
assign n7244 =  ( n7243 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7245 = ~ ( n7244 ) ;
assign n7246 =  ( n7242 ) ^ ( n7245 )  ;
assign n7247 =  ( n6483 ) | ( n6492 )  ;
assign n7248 =  ( n7247 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7249 =  ( n7246 ) ^ ( n7248 )  ;
assign n7250 =  ( n6030 ) | ( n6039 )  ;
assign n7251 =  ( n7250 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7252 =  ( n7249 ) ^ ( n7251 )  ;
assign n7253 =  ( n5802 ) | ( n5811 )  ;
assign n7254 =  ( n7253 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7255 =  ( n7252 ) ^ ( n7254 )  ;
assign n7256 =  ( n5832 ) | ( n5841 )  ;
assign n7257 =  ( n7256 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7258 =  ( n7255 ) ^ ( n7257 )  ;
assign n7259 = ~ ( n7258 ) ;
assign n7260 =  ( n5682 ) | ( n5691 )  ;
assign n7261 =  ( n7260 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7262 = ~ ( n7261 ) ;
assign n7263 =  ( n7259 ) | ( n7262 )  ;
assign n7264 = ~ ( n7263 ) ;
assign n7265 =  ( n7229 ) | ( n7264 )  ;
assign n7266 = ~ ( n7265 ) ;
assign n7267 = ~ ( n7169 ) ;
assign n7268 = ~ ( n6366 ) ;
assign n7269 =  ( n7267 ) | ( n7268 )  ;
assign n7270 = ~ ( n7269 ) ;
assign n7271 =  ( n7162 ) | ( n7270 )  ;
assign n7272 = ~ ( n7271 ) ;
assign n7273 = ~ ( n5736 ) ;
assign n7274 =  ( n7273 ) | ( n5742 )  ;
assign n7275 = ~ ( n7274 ) ;
assign n7276 = ~ ( n7193 ) ;
assign n7277 =  ( n7275 ) | ( n7276 )  ;
assign n7278 = ~ ( n7277 ) ;
assign n7279 =  ( n7272 ) | ( n7278 )  ;
assign n7280 = ~ ( n7279 ) ;
assign n7281 =  ( n7266 ) | ( n7280 )  ;
assign n7282 = ~ ( n7281 ) ;
assign n7283 = ~ ( n7271 ) ;
assign n7284 = ~ ( n7277 ) ;
assign n7285 =  ( n7283 ) | ( n7284 )  ;
assign n7286 =  ( n7265 ) ^ ( n7285 )  ;
assign n7287 = ~ ( n7286 ) ;
assign n7288 =  ( bv_1_1_n5 ) ^ ( n6888 )  ;
assign n7289 = ~ ( n6895 ) ;
assign n7290 = ~ ( n6366 ) ;
assign n7291 =  ( n7289 ) | ( n7290 )  ;
assign n7292 =  ( n7288 ) ^ ( n7291 )  ;
assign n7293 =  ( n6483 ) | ( n6492 )  ;
assign n7294 =  ( n7293 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7295 =  ( n7292 ) ^ ( n7294 )  ;
assign n7296 =  ( n6030 ) | ( n6039 )  ;
assign n7297 =  ( n7296 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7298 =  ( n7295 ) ^ ( n7297 )  ;
assign n7299 =  ( n5802 ) | ( n5811 )  ;
assign n7300 =  ( n7299 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7301 =  ( n7298 ) ^ ( n7300 )  ;
assign n7302 =  ( n5832 ) | ( n5841 )  ;
assign n7303 =  ( n7302 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7304 =  ( n7301 ) ^ ( n7303 )  ;
assign n7305 =  ( n5682 ) | ( n5691 )  ;
assign n7306 =  ( n7305 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7307 =  ( n7304 ) ^ ( n7306 )  ;
assign n7308 =  ( n5713 ) | ( n5722 )  ;
assign n7309 =  ( n7308 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7310 =  ( n7307 ) ^ ( n7309 )  ;
assign n7311 = ~ ( n7310 ) ;
assign n7312 =  ( n7287 ) | ( n7311 )  ;
assign n7313 = ~ ( n7312 ) ;
assign n7314 =  ( n7282 ) | ( n7313 )  ;
assign n7315 = ~ ( n7314 ) ;
assign n7316 = ~ ( n6977 ) ;
assign n7317 = ~ ( n6982 ) ;
assign n7318 =  ( n7316 ) | ( n7317 )  ;
assign n7319 =  ( n6970 ) ^ ( n7318 )  ;
assign n7320 = ~ ( n6517 ) ;
assign n7321 =  ( n6524 ) | ( n6150 )  ;
assign n7322 = ~ ( n7321 ) ;
assign n7323 =  ( n7320 ) | ( n7322 )  ;
assign n7324 = ~ ( n6543 ) ;
assign n7325 =  ( n7323 ) | ( n7324 )  ;
assign n7326 =  ( n7319 ) ^ ( n7325 )  ;
assign n7327 = ~ ( n6553 ) ;
assign n7328 = ~ ( n6173 ) ;
assign n7329 =  ( n7327 ) | ( n7328 )  ;
assign n7330 =  ( n7326 ) ^ ( n7329 )  ;
assign n7331 =  ( n6483 ) | ( n6492 )  ;
assign n7332 =  ( n7331 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7333 = ~ ( n7332 ) ;
assign n7334 =  ( n7330 ) ^ ( n7333 )  ;
assign n7335 =  ( n6030 ) | ( n6039 )  ;
assign n7336 =  ( n7335 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7337 =  ( n7334 ) ^ ( n7336 )  ;
assign n7338 =  ( n5802 ) | ( n5811 )  ;
assign n7339 =  ( n7338 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7340 =  ( n7337 ) ^ ( n7339 )  ;
assign n7341 =  ( n5832 ) | ( n5841 )  ;
assign n7342 =  ( n7341 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7343 =  ( n7340 ) ^ ( n7342 )  ;
assign n7344 =  ( n5682 ) | ( n5691 )  ;
assign n7345 =  ( n7344 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7346 =  ( n7343 ) ^ ( n7345 )  ;
assign n7347 = ~ ( n7346 ) ;
assign n7348 =  ( n7315 ) | ( n7347 )  ;
assign n7349 = ~ ( n7348 ) ;
assign n7350 = ~ ( n7281 ) ;
assign n7351 =  ( n7287 ) | ( n7311 )  ;
assign n7352 = ~ ( n7351 ) ;
assign n7353 =  ( n7350 ) | ( n7352 )  ;
assign n7354 =  ( n7353 ) ^ ( n6970 )  ;
assign n7355 = ~ ( n6977 ) ;
assign n7356 = ~ ( n6982 ) ;
assign n7357 =  ( n7355 ) | ( n7356 )  ;
assign n7358 =  ( n7354 ) ^ ( n7357 )  ;
assign n7359 = ~ ( n6517 ) ;
assign n7360 =  ( n6524 ) | ( n6150 )  ;
assign n7361 = ~ ( n7360 ) ;
assign n7362 =  ( n7359 ) | ( n7361 )  ;
assign n7363 = ~ ( n6543 ) ;
assign n7364 =  ( n7362 ) | ( n7363 )  ;
assign n7365 =  ( n7358 ) ^ ( n7364 )  ;
assign n7366 = ~ ( n6553 ) ;
assign n7367 = ~ ( n6173 ) ;
assign n7368 =  ( n7366 ) | ( n7367 )  ;
assign n7369 =  ( n7365 ) ^ ( n7368 )  ;
assign n7370 =  ( n6483 ) | ( n6492 )  ;
assign n7371 =  ( n7370 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7372 = ~ ( n7371 ) ;
assign n7373 =  ( n7369 ) ^ ( n7372 )  ;
assign n7374 =  ( n6030 ) | ( n6039 )  ;
assign n7375 =  ( n7374 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7376 =  ( n7373 ) ^ ( n7375 )  ;
assign n7377 =  ( n5802 ) | ( n5811 )  ;
assign n7378 =  ( n7377 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7379 =  ( n7376 ) ^ ( n7378 )  ;
assign n7380 =  ( n5832 ) | ( n5841 )  ;
assign n7381 =  ( n7380 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7382 =  ( n7379 ) ^ ( n7381 )  ;
assign n7383 =  ( n5682 ) | ( n5691 )  ;
assign n7384 =  ( n7383 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7385 =  ( n7382 ) ^ ( n7384 )  ;
assign n7386 = ~ ( n7385 ) ;
assign n7387 =  ( n5713 ) | ( n5722 )  ;
assign n7388 =  ( n7387 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7389 = ~ ( n7388 ) ;
assign n7390 =  ( n7386 ) | ( n7389 )  ;
assign n7391 = ~ ( n7390 ) ;
assign n7392 =  ( n7349 ) | ( n7391 )  ;
assign n7393 = ~ ( n7392 ) ;
assign n7394 =  ( n7118 ) | ( n7393 )  ;
assign n7395 =  ( bv_1_1_n5 ) ^ ( n7022 )  ;
assign n7396 =  ( n7395 ) ^ ( n6589 )  ;
assign n7397 =  ( n7396 ) ^ ( n6634 )  ;
assign n7398 = ~ ( n6640 ) ;
assign n7399 = ~ ( n6173 ) ;
assign n7400 =  ( n7398 ) | ( n7399 )  ;
assign n7401 =  ( n7397 ) ^ ( n7400 )  ;
assign n7402 =  ( n6030 ) | ( n6039 )  ;
assign n7403 =  ( n7402 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7404 =  ( n7401 ) ^ ( n7403 )  ;
assign n7405 =  ( n5802 ) | ( n5811 )  ;
assign n7406 =  ( n7405 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7407 =  ( n7404 ) ^ ( n7406 )  ;
assign n7408 =  ( n5832 ) | ( n5841 )  ;
assign n7409 =  ( n7408 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7410 =  ( n7407 ) ^ ( n7409 )  ;
assign n7411 =  ( n5682 ) | ( n5691 )  ;
assign n7412 =  ( n7411 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7413 =  ( n7410 ) ^ ( n7412 )  ;
assign n7414 =  ( n5713 ) | ( n5722 )  ;
assign n7415 =  ( n7414 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7416 =  ( n7413 ) ^ ( n7415 )  ;
assign n7417 = ~ ( n7416 ) ;
assign n7418 =  ( n7394 ) | ( n7417 )  ;
assign n7419 = ~ ( n7418 ) ;
assign n7420 =  ( n7081 ) | ( n7419 )  ;
assign n7421 = ~ ( n7117 ) ;
assign n7422 =  ( bv_1_1_n5 ) ^ ( n7392 )  ;
assign n7423 =  ( n7422 ) ^ ( n7022 )  ;
assign n7424 =  ( n7423 ) ^ ( n6589 )  ;
assign n7425 =  ( n7424 ) ^ ( n6634 )  ;
assign n7426 = ~ ( n6640 ) ;
assign n7427 = ~ ( n6173 ) ;
assign n7428 =  ( n7426 ) | ( n7427 )  ;
assign n7429 =  ( n7425 ) ^ ( n7428 )  ;
assign n7430 =  ( n6030 ) | ( n6039 )  ;
assign n7431 =  ( n7430 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7432 =  ( n7429 ) ^ ( n7431 )  ;
assign n7433 =  ( n5802 ) | ( n5811 )  ;
assign n7434 =  ( n7433 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7435 =  ( n7432 ) ^ ( n7434 )  ;
assign n7436 =  ( n5832 ) | ( n5841 )  ;
assign n7437 =  ( n7436 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7438 =  ( n7435 ) ^ ( n7437 )  ;
assign n7439 =  ( n5682 ) | ( n5691 )  ;
assign n7440 =  ( n7439 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7441 =  ( n7438 ) ^ ( n7440 )  ;
assign n7442 =  ( n5713 ) | ( n5722 )  ;
assign n7443 =  ( n7442 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7444 =  ( n7441 ) ^ ( n7443 )  ;
assign n7445 = ~ ( n7444 ) ;
assign n7446 =  ( n7421 ) | ( n7445 )  ;
assign n7447 = kd[1:1] ;
assign n7448 =  ( n7447 ) == ( bv_1_1_n5 )  ;
assign n7449 = kd[0:0] ;
assign n7450 =  ( n7449 ) == ( bv_1_1_n5 )  ;
assign n7451 =  ( n7448 ) | ( n7450 )  ;
assign n7452 = kd[1:1] ;
assign n7453 =  ( n7452 ) == ( bv_1_1_n5 )  ;
assign n7454 =  ( n7453 ) ? ( bv_1_1_n5 ) : ( bv_1_0_n2 ) ;
assign n7455 =  ( n7451 ) ? ( n7454 ) : ( bv_1_0_n2 ) ;
assign n7456 =  ( n6825 ) | ( n6834 )  ;
assign n7457 =  ( n7456 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7458 = ~ ( n7457 ) ;
assign n7459 =  ( n7455 ) | ( n7458 )  ;
assign n7460 =  ( n6483 ) | ( n6492 )  ;
assign n7461 =  ( n7460 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7462 = ~ ( n7461 ) ;
assign n7463 =  ( n7459 ) | ( n7462 )  ;
assign n7464 =  ( n6030 ) | ( n6039 )  ;
assign n7465 =  ( n7464 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7466 = ~ ( n7465 ) ;
assign n7467 =  ( n7463 ) | ( n7466 )  ;
assign n7468 = ~ ( n7467 ) ;
assign n7469 = ~ ( n7455 ) ;
assign n7470 =  ( n6825 ) | ( n6834 )  ;
assign n7471 =  ( n7470 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7472 =  ( n7469 ) ^ ( n7471 )  ;
assign n7473 = ~ ( n7472 ) ;
assign n7474 =  ( n7473 ) | ( n6524 )  ;
assign n7475 = ~ ( n7474 ) ;
assign n7476 =  ( n7468 ) | ( n7475 )  ;
assign n7477 = ~ ( n7455 ) ;
assign n7478 =  ( n6825 ) | ( n6834 )  ;
assign n7479 =  ( n7478 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7480 =  ( n7477 ) ^ ( n7479 )  ;
assign n7481 =  ( n6483 ) | ( n6492 )  ;
assign n7482 =  ( n7481 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7483 =  ( n7480 ) ^ ( n7482 )  ;
assign n7484 =  ( n6030 ) | ( n6039 )  ;
assign n7485 =  ( n7484 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7486 =  ( n7483 ) ^ ( n7485 )  ;
assign n7487 = ~ ( n7486 ) ;
assign n7488 =  ( n5802 ) | ( n5811 )  ;
assign n7489 =  ( n7488 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7490 = ~ ( n7489 ) ;
assign n7491 =  ( n7487 ) | ( n7490 )  ;
assign n7492 = ~ ( n7491 ) ;
assign n7493 =  ( n7476 ) | ( n7492 )  ;
assign n7494 = ~ ( n7493 ) ;
assign n7495 =  ( n6825 ) | ( n6834 )  ;
assign n7496 =  ( n7495 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7497 = ~ ( n7496 ) ;
assign n7498 =  ( n7455 ) | ( n7497 )  ;
assign n7499 = ~ ( n7498 ) ;
assign n7500 = ~ ( n6553 ) ;
assign n7501 =  ( n7499 ) | ( n7500 )  ;
assign n7502 = ~ ( n7501 ) ;
assign n7503 =  ( n7494 ) | ( n7502 )  ;
assign n7504 = ~ ( n5902 ) ;
assign n7505 = ~ ( n5913 ) ;
assign n7506 =  ( n7504 ) | ( n7505 )  ;
assign n7507 = ~ ( n7506 ) ;
assign n7508 =  ( n7503 ) | ( n7507 )  ;
assign n7509 =  ( n6825 ) | ( n6834 )  ;
assign n7510 =  ( n7509 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7511 =  ( n6483 ) | ( n6492 )  ;
assign n7512 =  ( n7511 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7513 =  ( n7510 ) ^ ( n7512 )  ;
assign n7514 =  ( n6030 ) | ( n6039 )  ;
assign n7515 =  ( n7514 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7516 =  ( n7513 ) ^ ( n7515 )  ;
assign n7517 =  ( n5802 ) | ( n5811 )  ;
assign n7518 =  ( n7517 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7519 =  ( n7516 ) ^ ( n7518 )  ;
assign n7520 =  ( n5832 ) | ( n5841 )  ;
assign n7521 =  ( n7520 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7522 =  ( n7519 ) ^ ( n7521 )  ;
assign n7523 = ~ ( n7522 ) ;
assign n7524 =  ( n7508 ) | ( n7523 )  ;
assign n7525 = ~ ( n7524 ) ;
assign n7526 = ~ ( n7467 ) ;
assign n7527 =  ( n7473 ) | ( n6524 )  ;
assign n7528 = ~ ( n7527 ) ;
assign n7529 =  ( n7526 ) | ( n7528 )  ;
assign n7530 = ~ ( n7491 ) ;
assign n7531 =  ( n7529 ) | ( n7530 )  ;
assign n7532 = ~ ( n7498 ) ;
assign n7533 = ~ ( n6553 ) ;
assign n7534 =  ( n7532 ) | ( n7533 )  ;
assign n7535 =  ( n7531 ) ^ ( n7534 )  ;
assign n7536 = ~ ( n7535 ) ;
assign n7537 = ~ ( n5902 ) ;
assign n7538 = ~ ( n5913 ) ;
assign n7539 =  ( n7537 ) | ( n7538 )  ;
assign n7540 =  ( n6825 ) | ( n6834 )  ;
assign n7541 =  ( n7540 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7542 =  ( n7539 ) ^ ( n7541 )  ;
assign n7543 =  ( n6483 ) | ( n6492 )  ;
assign n7544 =  ( n7543 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7545 =  ( n7542 ) ^ ( n7544 )  ;
assign n7546 =  ( n6030 ) | ( n6039 )  ;
assign n7547 =  ( n7546 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7548 =  ( n7545 ) ^ ( n7547 )  ;
assign n7549 =  ( n5802 ) | ( n5811 )  ;
assign n7550 =  ( n7549 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7551 =  ( n7548 ) ^ ( n7550 )  ;
assign n7552 =  ( n5832 ) | ( n5841 )  ;
assign n7553 =  ( n7552 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7554 =  ( n7551 ) ^ ( n7553 )  ;
assign n7555 = ~ ( n7554 ) ;
assign n7556 =  ( n7536 ) | ( n7555 )  ;
assign n7557 = ~ ( n7556 ) ;
assign n7558 =  ( n7525 ) | ( n7557 )  ;
assign n7559 = ~ ( n7467 ) ;
assign n7560 =  ( n7473 ) | ( n6524 )  ;
assign n7561 = ~ ( n7560 ) ;
assign n7562 =  ( n7559 ) | ( n7561 )  ;
assign n7563 = ~ ( n7491 ) ;
assign n7564 =  ( n7562 ) | ( n7563 )  ;
assign n7565 = ~ ( n7498 ) ;
assign n7566 = ~ ( n6553 ) ;
assign n7567 =  ( n7565 ) | ( n7566 )  ;
assign n7568 =  ( n7564 ) ^ ( n7567 )  ;
assign n7569 = ~ ( n5902 ) ;
assign n7570 = ~ ( n5913 ) ;
assign n7571 =  ( n7569 ) | ( n7570 )  ;
assign n7572 =  ( n7568 ) ^ ( n7571 )  ;
assign n7573 =  ( n6825 ) | ( n6834 )  ;
assign n7574 =  ( n7573 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7575 =  ( n7572 ) ^ ( n7574 )  ;
assign n7576 =  ( n6483 ) | ( n6492 )  ;
assign n7577 =  ( n7576 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7578 =  ( n7575 ) ^ ( n7577 )  ;
assign n7579 =  ( n6030 ) | ( n6039 )  ;
assign n7580 =  ( n7579 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7581 =  ( n7578 ) ^ ( n7580 )  ;
assign n7582 =  ( n5802 ) | ( n5811 )  ;
assign n7583 =  ( n7582 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7584 =  ( n7581 ) ^ ( n7583 )  ;
assign n7585 =  ( n5832 ) | ( n5841 )  ;
assign n7586 =  ( n7585 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7587 =  ( n7584 ) ^ ( n7586 )  ;
assign n7588 = ~ ( n7587 ) ;
assign n7589 =  ( n7588 ) | ( n5972 )  ;
assign n7590 = ~ ( n7589 ) ;
assign n7591 =  ( n7558 ) | ( n7590 )  ;
assign n7592 = ~ ( n7591 ) ;
assign n7593 = ~ ( n7498 ) ;
assign n7594 = ~ ( n6553 ) ;
assign n7595 =  ( n7593 ) | ( n7594 )  ;
assign n7596 = ~ ( n7595 ) ;
assign n7597 =  ( n7494 ) | ( n7596 )  ;
assign n7598 = ~ ( n7597 ) ;
assign n7599 = ~ ( n5902 ) ;
assign n7600 = ~ ( n5913 ) ;
assign n7601 =  ( n7599 ) | ( n7600 )  ;
assign n7602 = ~ ( n7601 ) ;
assign n7603 =  ( n7602 ) | ( n7523 )  ;
assign n7604 = ~ ( n7603 ) ;
assign n7605 =  ( n7598 ) | ( n7604 )  ;
assign n7606 = ~ ( n7605 ) ;
assign n7607 =  ( n7592 ) | ( n7606 )  ;
assign n7608 = ~ ( n7607 ) ;
assign n7609 = ~ ( n7597 ) ;
assign n7610 = ~ ( n7603 ) ;
assign n7611 =  ( n7609 ) | ( n7610 )  ;
assign n7612 =  ( n7591 ) ^ ( n7611 )  ;
assign n7613 = ~ ( n7612 ) ;
assign n7614 = ~ ( n7133 ) ;
assign n7615 =  ( n7140 ) | ( n6337 )  ;
assign n7616 = ~ ( n7615 ) ;
assign n7617 =  ( n7614 ) | ( n7616 )  ;
assign n7618 = ~ ( n7159 ) ;
assign n7619 =  ( n7617 ) | ( n7618 )  ;
assign n7620 = ~ ( n7169 ) ;
assign n7621 = ~ ( n6366 ) ;
assign n7622 =  ( n7620 ) | ( n7621 )  ;
assign n7623 =  ( n7619 ) ^ ( n7622 )  ;
assign n7624 = ~ ( n5736 ) ;
assign n7625 =  ( n7624 ) | ( n5742 )  ;
assign n7626 =  ( n7623 ) ^ ( n7625 )  ;
assign n7627 =  ( n6825 ) | ( n6834 )  ;
assign n7628 =  ( n7627 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7629 = ~ ( n7628 ) ;
assign n7630 =  ( n7626 ) ^ ( n7629 )  ;
assign n7631 =  ( n6483 ) | ( n6492 )  ;
assign n7632 =  ( n7631 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7633 =  ( n7630 ) ^ ( n7632 )  ;
assign n7634 =  ( n6030 ) | ( n6039 )  ;
assign n7635 =  ( n7634 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7636 =  ( n7633 ) ^ ( n7635 )  ;
assign n7637 =  ( n5802 ) | ( n5811 )  ;
assign n7638 =  ( n7637 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7639 =  ( n7636 ) ^ ( n7638 )  ;
assign n7640 =  ( n5832 ) | ( n5841 )  ;
assign n7641 =  ( n7640 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7642 =  ( n7639 ) ^ ( n7641 )  ;
assign n7643 =  ( n5682 ) | ( n5691 )  ;
assign n7644 =  ( n7643 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7645 =  ( n7642 ) ^ ( n7644 )  ;
assign n7646 = ~ ( n7645 ) ;
assign n7647 =  ( n7613 ) | ( n7646 )  ;
assign n7648 = ~ ( n7647 ) ;
assign n7649 =  ( n7608 ) | ( n7648 )  ;
assign n7650 = ~ ( n7649 ) ;
assign n7651 =  ( bv_1_1_n5 ) ^ ( n7265 )  ;
assign n7652 = ~ ( n7271 ) ;
assign n7653 = ~ ( n7277 ) ;
assign n7654 =  ( n7652 ) | ( n7653 )  ;
assign n7655 =  ( n7651 ) ^ ( n7654 )  ;
assign n7656 =  ( n7655 ) ^ ( n6888 )  ;
assign n7657 = ~ ( n6895 ) ;
assign n7658 = ~ ( n6366 ) ;
assign n7659 =  ( n7657 ) | ( n7658 )  ;
assign n7660 =  ( n7656 ) ^ ( n7659 )  ;
assign n7661 =  ( n6483 ) | ( n6492 )  ;
assign n7662 =  ( n7661 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7663 =  ( n7660 ) ^ ( n7662 )  ;
assign n7664 =  ( n6030 ) | ( n6039 )  ;
assign n7665 =  ( n7664 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7666 =  ( n7663 ) ^ ( n7665 )  ;
assign n7667 =  ( n5802 ) | ( n5811 )  ;
assign n7668 =  ( n7667 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7669 =  ( n7666 ) ^ ( n7668 )  ;
assign n7670 =  ( n5832 ) | ( n5841 )  ;
assign n7671 =  ( n7670 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7672 =  ( n7669 ) ^ ( n7671 )  ;
assign n7673 =  ( n5682 ) | ( n5691 )  ;
assign n7674 =  ( n7673 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7675 =  ( n7672 ) ^ ( n7674 )  ;
assign n7676 =  ( n5713 ) | ( n5722 )  ;
assign n7677 =  ( n7676 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7678 =  ( n7675 ) ^ ( n7677 )  ;
assign n7679 = ~ ( n7678 ) ;
assign n7680 =  ( n7650 ) | ( n7679 )  ;
assign n7681 = ~ ( n7281 ) ;
assign n7682 =  ( n7287 ) | ( n7311 )  ;
assign n7683 = ~ ( n7682 ) ;
assign n7684 =  ( n7681 ) | ( n7683 )  ;
assign n7685 =  ( n7684 ) ^ ( n6970 )  ;
assign n7686 = ~ ( n6977 ) ;
assign n7687 = ~ ( n6982 ) ;
assign n7688 =  ( n7686 ) | ( n7687 )  ;
assign n7689 =  ( n7685 ) ^ ( n7688 )  ;
assign n7690 = ~ ( n6517 ) ;
assign n7691 =  ( n6524 ) | ( n6150 )  ;
assign n7692 = ~ ( n7691 ) ;
assign n7693 =  ( n7690 ) | ( n7692 )  ;
assign n7694 = ~ ( n6543 ) ;
assign n7695 =  ( n7693 ) | ( n7694 )  ;
assign n7696 =  ( n7689 ) ^ ( n7695 )  ;
assign n7697 = ~ ( n6553 ) ;
assign n7698 = ~ ( n6173 ) ;
assign n7699 =  ( n7697 ) | ( n7698 )  ;
assign n7700 =  ( n7696 ) ^ ( n7699 )  ;
assign n7701 =  ( n6483 ) | ( n6492 )  ;
assign n7702 =  ( n7701 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7703 = ~ ( n7702 ) ;
assign n7704 =  ( n7700 ) ^ ( n7703 )  ;
assign n7705 =  ( n6030 ) | ( n6039 )  ;
assign n7706 =  ( n7705 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7707 =  ( n7704 ) ^ ( n7706 )  ;
assign n7708 =  ( n5802 ) | ( n5811 )  ;
assign n7709 =  ( n7708 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7710 =  ( n7707 ) ^ ( n7709 )  ;
assign n7711 =  ( n5832 ) | ( n5841 )  ;
assign n7712 =  ( n7711 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7713 =  ( n7710 ) ^ ( n7712 )  ;
assign n7714 =  ( n5682 ) | ( n5691 )  ;
assign n7715 =  ( n7714 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7716 =  ( n7713 ) ^ ( n7715 )  ;
assign n7717 =  ( n5713 ) | ( n5722 )  ;
assign n7718 =  ( n7717 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7719 =  ( n7716 ) ^ ( n7718 )  ;
assign n7720 = ~ ( n7719 ) ;
assign n7721 =  ( n7680 ) | ( n7720 )  ;
assign n7722 = ~ ( n7721 ) ;
assign n7723 = ~ ( n7649 ) ;
assign n7724 =  ( n7723 ) | ( n7679 )  ;
assign n7725 = ~ ( n7724 ) ;
assign n7726 = ~ ( n7281 ) ;
assign n7727 =  ( n7287 ) | ( n7311 )  ;
assign n7728 = ~ ( n7727 ) ;
assign n7729 =  ( n7726 ) | ( n7728 )  ;
assign n7730 =  ( n7725 ) ^ ( n7729 )  ;
assign n7731 =  ( n7730 ) ^ ( n6970 )  ;
assign n7732 = ~ ( n6977 ) ;
assign n7733 = ~ ( n6982 ) ;
assign n7734 =  ( n7732 ) | ( n7733 )  ;
assign n7735 =  ( n7731 ) ^ ( n7734 )  ;
assign n7736 = ~ ( n6517 ) ;
assign n7737 =  ( n6524 ) | ( n6150 )  ;
assign n7738 = ~ ( n7737 ) ;
assign n7739 =  ( n7736 ) | ( n7738 )  ;
assign n7740 = ~ ( n6543 ) ;
assign n7741 =  ( n7739 ) | ( n7740 )  ;
assign n7742 =  ( n7735 ) ^ ( n7741 )  ;
assign n7743 = ~ ( n6553 ) ;
assign n7744 = ~ ( n6173 ) ;
assign n7745 =  ( n7743 ) | ( n7744 )  ;
assign n7746 =  ( n7742 ) ^ ( n7745 )  ;
assign n7747 =  ( n6483 ) | ( n6492 )  ;
assign n7748 =  ( n7747 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7749 = ~ ( n7748 ) ;
assign n7750 =  ( n7746 ) ^ ( n7749 )  ;
assign n7751 =  ( n6030 ) | ( n6039 )  ;
assign n7752 =  ( n7751 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7753 =  ( n7750 ) ^ ( n7752 )  ;
assign n7754 =  ( n5802 ) | ( n5811 )  ;
assign n7755 =  ( n7754 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7756 =  ( n7753 ) ^ ( n7755 )  ;
assign n7757 =  ( n5832 ) | ( n5841 )  ;
assign n7758 =  ( n7757 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7759 =  ( n7756 ) ^ ( n7758 )  ;
assign n7760 =  ( n5682 ) | ( n5691 )  ;
assign n7761 =  ( n7760 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7762 =  ( n7759 ) ^ ( n7761 )  ;
assign n7763 =  ( n5713 ) | ( n5722 )  ;
assign n7764 =  ( n7763 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7765 =  ( n7762 ) ^ ( n7764 )  ;
assign n7766 = ~ ( n7765 ) ;
assign n7767 = ~ ( n7455 ) ;
assign n7768 =  ( n6825 ) | ( n6834 )  ;
assign n7769 =  ( n7768 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7770 = ~ ( n7769 ) ;
assign n7771 =  ( n7767 ) | ( n7770 )  ;
assign n7772 =  ( n6483 ) | ( n6492 )  ;
assign n7773 =  ( n7772 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7774 = ~ ( n7773 ) ;
assign n7775 =  ( n7771 ) | ( n7774 )  ;
assign n7776 =  ( n6030 ) | ( n6039 )  ;
assign n7777 =  ( n7776 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7778 = ~ ( n7777 ) ;
assign n7779 =  ( n7775 ) | ( n7778 )  ;
assign n7780 = ~ ( n7779 ) ;
assign n7781 =  ( n6825 ) | ( n6834 )  ;
assign n7782 =  ( n7781 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7783 =  ( n7455 ) ^ ( n7782 )  ;
assign n7784 = ~ ( n7783 ) ;
assign n7785 =  ( n7784 ) | ( n6524 )  ;
assign n7786 = ~ ( n7785 ) ;
assign n7787 =  ( n7780 ) | ( n7786 )  ;
assign n7788 =  ( n6825 ) | ( n6834 )  ;
assign n7789 =  ( n7788 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7790 =  ( n7455 ) ^ ( n7789 )  ;
assign n7791 =  ( n6483 ) | ( n6492 )  ;
assign n7792 =  ( n7791 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7793 =  ( n7790 ) ^ ( n7792 )  ;
assign n7794 =  ( n6030 ) | ( n6039 )  ;
assign n7795 =  ( n7794 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7796 =  ( n7793 ) ^ ( n7795 )  ;
assign n7797 = ~ ( n7796 ) ;
assign n7798 =  ( n5802 ) | ( n5811 )  ;
assign n7799 =  ( n7798 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7800 = ~ ( n7799 ) ;
assign n7801 =  ( n7797 ) | ( n7800 )  ;
assign n7802 = ~ ( n7801 ) ;
assign n7803 =  ( n7787 ) | ( n7802 )  ;
assign n7804 = ~ ( n7803 ) ;
assign n7805 = ~ ( n7455 ) ;
assign n7806 =  ( n6825 ) | ( n6834 )  ;
assign n7807 =  ( n7806 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7808 = ~ ( n7807 ) ;
assign n7809 =  ( n7805 ) | ( n7808 )  ;
assign n7810 = ~ ( n7809 ) ;
assign n7811 = ~ ( n6553 ) ;
assign n7812 =  ( n7810 ) | ( n7811 )  ;
assign n7813 = ~ ( n7812 ) ;
assign n7814 =  ( n7804 ) | ( n7813 )  ;
assign n7815 = ~ ( n5902 ) ;
assign n7816 = ~ ( n5913 ) ;
assign n7817 =  ( n7815 ) | ( n7816 )  ;
assign n7818 = ~ ( n7817 ) ;
assign n7819 =  ( n7814 ) | ( n7818 )  ;
assign n7820 = ~ ( n7455 ) ;
assign n7821 =  ( n6825 ) | ( n6834 )  ;
assign n7822 =  ( n7821 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7823 =  ( n7820 ) ^ ( n7822 )  ;
assign n7824 =  ( n6483 ) | ( n6492 )  ;
assign n7825 =  ( n7824 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7826 =  ( n7823 ) ^ ( n7825 )  ;
assign n7827 =  ( n6030 ) | ( n6039 )  ;
assign n7828 =  ( n7827 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7829 =  ( n7826 ) ^ ( n7828 )  ;
assign n7830 =  ( n5802 ) | ( n5811 )  ;
assign n7831 =  ( n7830 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7832 =  ( n7829 ) ^ ( n7831 )  ;
assign n7833 = ~ ( n7832 ) ;
assign n7834 =  ( n7819 ) | ( n7833 )  ;
assign n7835 = ~ ( n7834 ) ;
assign n7836 = ~ ( n7779 ) ;
assign n7837 =  ( n7784 ) | ( n6524 )  ;
assign n7838 = ~ ( n7837 ) ;
assign n7839 =  ( n7836 ) | ( n7838 )  ;
assign n7840 = ~ ( n7801 ) ;
assign n7841 =  ( n7839 ) | ( n7840 )  ;
assign n7842 = ~ ( n7809 ) ;
assign n7843 = ~ ( n6553 ) ;
assign n7844 =  ( n7842 ) | ( n7843 )  ;
assign n7845 =  ( n7841 ) ^ ( n7844 )  ;
assign n7846 = ~ ( n7845 ) ;
assign n7847 = ~ ( n5902 ) ;
assign n7848 = ~ ( n5913 ) ;
assign n7849 =  ( n7847 ) | ( n7848 )  ;
assign n7850 = ~ ( n7455 ) ;
assign n7851 =  ( n7849 ) ^ ( n7850 )  ;
assign n7852 =  ( n6825 ) | ( n6834 )  ;
assign n7853 =  ( n7852 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7854 =  ( n7851 ) ^ ( n7853 )  ;
assign n7855 =  ( n6483 ) | ( n6492 )  ;
assign n7856 =  ( n7855 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7857 =  ( n7854 ) ^ ( n7856 )  ;
assign n7858 =  ( n6030 ) | ( n6039 )  ;
assign n7859 =  ( n7858 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7860 =  ( n7857 ) ^ ( n7859 )  ;
assign n7861 =  ( n5802 ) | ( n5811 )  ;
assign n7862 =  ( n7861 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7863 =  ( n7860 ) ^ ( n7862 )  ;
assign n7864 = ~ ( n7863 ) ;
assign n7865 =  ( n7846 ) | ( n7864 )  ;
assign n7866 = ~ ( n7865 ) ;
assign n7867 =  ( n7835 ) | ( n7866 )  ;
assign n7868 = ~ ( n7779 ) ;
assign n7869 =  ( n7784 ) | ( n6524 )  ;
assign n7870 = ~ ( n7869 ) ;
assign n7871 =  ( n7868 ) | ( n7870 )  ;
assign n7872 = ~ ( n7801 ) ;
assign n7873 =  ( n7871 ) | ( n7872 )  ;
assign n7874 = ~ ( n7809 ) ;
assign n7875 = ~ ( n6553 ) ;
assign n7876 =  ( n7874 ) | ( n7875 )  ;
assign n7877 =  ( n7873 ) ^ ( n7876 )  ;
assign n7878 = ~ ( n5902 ) ;
assign n7879 = ~ ( n5913 ) ;
assign n7880 =  ( n7878 ) | ( n7879 )  ;
assign n7881 =  ( n7877 ) ^ ( n7880 )  ;
assign n7882 = ~ ( n7455 ) ;
assign n7883 =  ( n7881 ) ^ ( n7882 )  ;
assign n7884 =  ( n6825 ) | ( n6834 )  ;
assign n7885 =  ( n7884 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7886 =  ( n7883 ) ^ ( n7885 )  ;
assign n7887 =  ( n6483 ) | ( n6492 )  ;
assign n7888 =  ( n7887 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7889 =  ( n7886 ) ^ ( n7888 )  ;
assign n7890 =  ( n6030 ) | ( n6039 )  ;
assign n7891 =  ( n7890 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7892 =  ( n7889 ) ^ ( n7891 )  ;
assign n7893 =  ( n5802 ) | ( n5811 )  ;
assign n7894 =  ( n7893 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7895 =  ( n7892 ) ^ ( n7894 )  ;
assign n7896 = ~ ( n7895 ) ;
assign n7897 =  ( n7896 ) | ( n5879 )  ;
assign n7898 = ~ ( n7897 ) ;
assign n7899 =  ( n7867 ) | ( n7898 )  ;
assign n7900 = ~ ( n7899 ) ;
assign n7901 = ~ ( n7809 ) ;
assign n7902 = ~ ( n6553 ) ;
assign n7903 =  ( n7901 ) | ( n7902 )  ;
assign n7904 = ~ ( n7903 ) ;
assign n7905 =  ( n7804 ) | ( n7904 )  ;
assign n7906 = ~ ( n7905 ) ;
assign n7907 = ~ ( n5902 ) ;
assign n7908 = ~ ( n5913 ) ;
assign n7909 =  ( n7907 ) | ( n7908 )  ;
assign n7910 = ~ ( n7909 ) ;
assign n7911 =  ( n7910 ) | ( n7833 )  ;
assign n7912 = ~ ( n7911 ) ;
assign n7913 =  ( n7906 ) | ( n7912 )  ;
assign n7914 = ~ ( n7913 ) ;
assign n7915 =  ( n7900 ) | ( n7914 )  ;
assign n7916 = ~ ( n7915 ) ;
assign n7917 = ~ ( n7905 ) ;
assign n7918 = ~ ( n7911 ) ;
assign n7919 =  ( n7917 ) | ( n7918 )  ;
assign n7920 =  ( n7899 ) ^ ( n7919 )  ;
assign n7921 = ~ ( n7920 ) ;
assign n7922 = ~ ( n7467 ) ;
assign n7923 =  ( n7473 ) | ( n6524 )  ;
assign n7924 = ~ ( n7923 ) ;
assign n7925 =  ( n7922 ) | ( n7924 )  ;
assign n7926 = ~ ( n7491 ) ;
assign n7927 =  ( n7925 ) | ( n7926 )  ;
assign n7928 =  ( bv_1_1_n5 ) ^ ( n7927 )  ;
assign n7929 = ~ ( n7498 ) ;
assign n7930 = ~ ( n6553 ) ;
assign n7931 =  ( n7929 ) | ( n7930 )  ;
assign n7932 =  ( n7928 ) ^ ( n7931 )  ;
assign n7933 = ~ ( n5902 ) ;
assign n7934 = ~ ( n5913 ) ;
assign n7935 =  ( n7933 ) | ( n7934 )  ;
assign n7936 =  ( n7932 ) ^ ( n7935 )  ;
assign n7937 =  ( n6825 ) | ( n6834 )  ;
assign n7938 =  ( n7937 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7939 =  ( n7936 ) ^ ( n7938 )  ;
assign n7940 =  ( n6483 ) | ( n6492 )  ;
assign n7941 =  ( n7940 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7942 =  ( n7939 ) ^ ( n7941 )  ;
assign n7943 =  ( n6030 ) | ( n6039 )  ;
assign n7944 =  ( n7943 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7945 =  ( n7942 ) ^ ( n7944 )  ;
assign n7946 =  ( n5802 ) | ( n5811 )  ;
assign n7947 =  ( n7946 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7948 =  ( n7945 ) ^ ( n7947 )  ;
assign n7949 =  ( n5832 ) | ( n5841 )  ;
assign n7950 =  ( n7949 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7951 =  ( n7948 ) ^ ( n7950 )  ;
assign n7952 =  ( n5682 ) | ( n5691 )  ;
assign n7953 =  ( n7952 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7954 =  ( n7951 ) ^ ( n7953 )  ;
assign n7955 =  ( n5713 ) | ( n5722 )  ;
assign n7956 =  ( n7955 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n7957 =  ( n7954 ) ^ ( n7956 )  ;
assign n7958 = ~ ( n7957 ) ;
assign n7959 =  ( n7921 ) | ( n7958 )  ;
assign n7960 = ~ ( n7959 ) ;
assign n7961 =  ( n7916 ) | ( n7960 )  ;
assign n7962 = ~ ( n7961 ) ;
assign n7963 = ~ ( n7597 ) ;
assign n7964 = ~ ( n7603 ) ;
assign n7965 =  ( n7963 ) | ( n7964 )  ;
assign n7966 =  ( n7591 ) ^ ( n7965 )  ;
assign n7967 = ~ ( n7133 ) ;
assign n7968 =  ( n7140 ) | ( n6337 )  ;
assign n7969 = ~ ( n7968 ) ;
assign n7970 =  ( n7967 ) | ( n7969 )  ;
assign n7971 = ~ ( n7159 ) ;
assign n7972 =  ( n7970 ) | ( n7971 )  ;
assign n7973 =  ( n7966 ) ^ ( n7972 )  ;
assign n7974 = ~ ( n7169 ) ;
assign n7975 = ~ ( n6366 ) ;
assign n7976 =  ( n7974 ) | ( n7975 )  ;
assign n7977 =  ( n7973 ) ^ ( n7976 )  ;
assign n7978 = ~ ( n5736 ) ;
assign n7979 =  ( n7978 ) | ( n5742 )  ;
assign n7980 =  ( n7977 ) ^ ( n7979 )  ;
assign n7981 =  ( n6825 ) | ( n6834 )  ;
assign n7982 =  ( n7981 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n7983 = ~ ( n7982 ) ;
assign n7984 =  ( n7980 ) ^ ( n7983 )  ;
assign n7985 =  ( n6483 ) | ( n6492 )  ;
assign n7986 =  ( n7985 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n7987 =  ( n7984 ) ^ ( n7986 )  ;
assign n7988 =  ( n6030 ) | ( n6039 )  ;
assign n7989 =  ( n7988 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n7990 =  ( n7987 ) ^ ( n7989 )  ;
assign n7991 =  ( n5802 ) | ( n5811 )  ;
assign n7992 =  ( n7991 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n7993 =  ( n7990 ) ^ ( n7992 )  ;
assign n7994 =  ( n5832 ) | ( n5841 )  ;
assign n7995 =  ( n7994 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n7996 =  ( n7993 ) ^ ( n7995 )  ;
assign n7997 =  ( n5682 ) | ( n5691 )  ;
assign n7998 =  ( n7997 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n7999 =  ( n7996 ) ^ ( n7998 )  ;
assign n8000 = ~ ( n7999 ) ;
assign n8001 =  ( n7962 ) | ( n8000 )  ;
assign n8002 = ~ ( n8001 ) ;
assign n8003 =  ( n7961 ) ^ ( n7591 )  ;
assign n8004 = ~ ( n7597 ) ;
assign n8005 = ~ ( n7603 ) ;
assign n8006 =  ( n8004 ) | ( n8005 )  ;
assign n8007 =  ( n8003 ) ^ ( n8006 )  ;
assign n8008 = ~ ( n7133 ) ;
assign n8009 =  ( n7140 ) | ( n6337 )  ;
assign n8010 = ~ ( n8009 ) ;
assign n8011 =  ( n8008 ) | ( n8010 )  ;
assign n8012 = ~ ( n7159 ) ;
assign n8013 =  ( n8011 ) | ( n8012 )  ;
assign n8014 =  ( n8007 ) ^ ( n8013 )  ;
assign n8015 = ~ ( n7169 ) ;
assign n8016 = ~ ( n6366 ) ;
assign n8017 =  ( n8015 ) | ( n8016 )  ;
assign n8018 =  ( n8014 ) ^ ( n8017 )  ;
assign n8019 = ~ ( n5736 ) ;
assign n8020 =  ( n8019 ) | ( n5742 )  ;
assign n8021 =  ( n8018 ) ^ ( n8020 )  ;
assign n8022 =  ( n6825 ) | ( n6834 )  ;
assign n8023 =  ( n8022 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8024 = ~ ( n8023 ) ;
assign n8025 =  ( n8021 ) ^ ( n8024 )  ;
assign n8026 =  ( n6483 ) | ( n6492 )  ;
assign n8027 =  ( n8026 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8028 =  ( n8025 ) ^ ( n8027 )  ;
assign n8029 =  ( n6030 ) | ( n6039 )  ;
assign n8030 =  ( n8029 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8031 =  ( n8028 ) ^ ( n8030 )  ;
assign n8032 =  ( n5802 ) | ( n5811 )  ;
assign n8033 =  ( n8032 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8034 =  ( n8031 ) ^ ( n8033 )  ;
assign n8035 =  ( n5832 ) | ( n5841 )  ;
assign n8036 =  ( n8035 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8037 =  ( n8034 ) ^ ( n8036 )  ;
assign n8038 =  ( n5682 ) | ( n5691 )  ;
assign n8039 =  ( n8038 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8040 =  ( n8037 ) ^ ( n8039 )  ;
assign n8041 = ~ ( n8040 ) ;
assign n8042 =  ( n5713 ) | ( n5722 )  ;
assign n8043 =  ( n8042 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8044 = ~ ( n8043 ) ;
assign n8045 =  ( n8041 ) | ( n8044 )  ;
assign n8046 = ~ ( n8045 ) ;
assign n8047 =  ( n8002 ) | ( n8046 )  ;
assign n8048 = ~ ( n8047 ) ;
assign n8049 =  ( n7766 ) | ( n8048 )  ;
assign n8050 =  ( bv_1_1_n5 ) ^ ( n7649 )  ;
assign n8051 =  ( n8050 ) ^ ( n7265 )  ;
assign n8052 = ~ ( n7271 ) ;
assign n8053 = ~ ( n7277 ) ;
assign n8054 =  ( n8052 ) | ( n8053 )  ;
assign n8055 =  ( n8051 ) ^ ( n8054 )  ;
assign n8056 =  ( n8055 ) ^ ( n6888 )  ;
assign n8057 = ~ ( n6895 ) ;
assign n8058 = ~ ( n6366 ) ;
assign n8059 =  ( n8057 ) | ( n8058 )  ;
assign n8060 =  ( n8056 ) ^ ( n8059 )  ;
assign n8061 =  ( n6483 ) | ( n6492 )  ;
assign n8062 =  ( n8061 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8063 =  ( n8060 ) ^ ( n8062 )  ;
assign n8064 =  ( n6030 ) | ( n6039 )  ;
assign n8065 =  ( n8064 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8066 =  ( n8063 ) ^ ( n8065 )  ;
assign n8067 =  ( n5802 ) | ( n5811 )  ;
assign n8068 =  ( n8067 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8069 =  ( n8066 ) ^ ( n8068 )  ;
assign n8070 =  ( n5832 ) | ( n5841 )  ;
assign n8071 =  ( n8070 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8072 =  ( n8069 ) ^ ( n8071 )  ;
assign n8073 =  ( n5682 ) | ( n5691 )  ;
assign n8074 =  ( n8073 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8075 =  ( n8072 ) ^ ( n8074 )  ;
assign n8076 =  ( n5713 ) | ( n5722 )  ;
assign n8077 =  ( n8076 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8078 =  ( n8075 ) ^ ( n8077 )  ;
assign n8079 = ~ ( n8078 ) ;
assign n8080 =  ( n8049 ) | ( n8079 )  ;
assign n8081 = ~ ( n8080 ) ;
assign n8082 =  ( n7722 ) | ( n8081 )  ;
assign n8083 = ~ ( n8082 ) ;
assign n8084 =  ( n7446 ) | ( n8083 )  ;
assign n8085 = ~ ( n8084 ) ;
assign n8086 =  ( n7420 ) | ( n8085 )  ;
assign n8087 = ~ ( n7117 ) ;
assign n8088 =  ( n8087 ) | ( n7445 )  ;
assign n8089 = ~ ( n7765 ) ;
assign n8090 =  ( n8088 ) | ( n8089 )  ;
assign n8091 =  ( bv_1_1_n5 ) ^ ( n8047 )  ;
assign n8092 =  ( n8091 ) ^ ( n7649 )  ;
assign n8093 =  ( n8092 ) ^ ( n7265 )  ;
assign n8094 = ~ ( n7271 ) ;
assign n8095 = ~ ( n7277 ) ;
assign n8096 =  ( n8094 ) | ( n8095 )  ;
assign n8097 =  ( n8093 ) ^ ( n8096 )  ;
assign n8098 =  ( n8097 ) ^ ( n6888 )  ;
assign n8099 = ~ ( n6895 ) ;
assign n8100 = ~ ( n6366 ) ;
assign n8101 =  ( n8099 ) | ( n8100 )  ;
assign n8102 =  ( n8098 ) ^ ( n8101 )  ;
assign n8103 =  ( n6483 ) | ( n6492 )  ;
assign n8104 =  ( n8103 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8105 =  ( n8102 ) ^ ( n8104 )  ;
assign n8106 =  ( n6030 ) | ( n6039 )  ;
assign n8107 =  ( n8106 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8108 =  ( n8105 ) ^ ( n8107 )  ;
assign n8109 =  ( n5802 ) | ( n5811 )  ;
assign n8110 =  ( n8109 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8111 =  ( n8108 ) ^ ( n8110 )  ;
assign n8112 =  ( n5832 ) | ( n5841 )  ;
assign n8113 =  ( n8112 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8114 =  ( n8111 ) ^ ( n8113 )  ;
assign n8115 =  ( n5682 ) | ( n5691 )  ;
assign n8116 =  ( n8115 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8117 =  ( n8114 ) ^ ( n8116 )  ;
assign n8118 =  ( n5713 ) | ( n5722 )  ;
assign n8119 =  ( n8118 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8120 =  ( n8117 ) ^ ( n8119 )  ;
assign n8121 = ~ ( n8120 ) ;
assign n8122 =  ( n8090 ) | ( n8121 )  ;
assign n8123 = ~ ( n7809 ) ;
assign n8124 = ~ ( n6553 ) ;
assign n8125 =  ( n8123 ) | ( n8124 )  ;
assign n8126 = ~ ( n8125 ) ;
assign n8127 =  ( n7804 ) | ( n8126 )  ;
assign n8128 = ~ ( n5902 ) ;
assign n8129 = kd[14:14] ;
assign n8130 =  ( n8129 ) == ( bv_1_1_n5 )  ;
assign n8131 = kd[13:13] ;
assign n8132 =  ( n8131 ) == ( bv_1_1_n5 )  ;
assign n8133 =  ( n8130 ) | ( n8132 )  ;
assign n8134 = kd[15:15] ;
assign n8135 =  ( n8134 ) == ( bv_1_0_n2 )  ;
assign n8136 =  ( n8133 ) | ( n8135 )  ;
assign n8137 = ~ ( n8136 )  ;
assign n8138 = kd[15:15] ;
assign n8139 =  ( n8138 ) == ( bv_1_1_n5 )  ;
assign n8140 = kd[14:14] ;
assign n8141 =  ( n8140 ) == ( bv_1_0_n2 )  ;
assign n8142 =  ( n8139 ) | ( n8141 )  ;
assign n8143 = kd[13:13] ;
assign n8144 =  ( n8143 ) == ( bv_1_0_n2 )  ;
assign n8145 =  ( n8142 ) | ( n8144 )  ;
assign n8146 = ~ ( n8145 )  ;
assign n8147 =  ( n8137 ) | ( n8146 )  ;
assign n8148 = kd[15:15] ;
assign n8149 = ~ ( n8148 ) ;
assign n8150 = kd[14:14] ;
assign n8151 = ~ ( n8150 ) ;
assign n8152 = kd[13:13] ;
assign n8153 = ~ ( n8152 ) ;
assign n8154 =  ( n8151 ) | ( n8153 )  ;
assign n8155 = ~ ( n8154 ) ;
assign n8156 =  ( n8149 ) | ( n8155 )  ;
assign n8157 = ~ ( n8156 ) ;
assign n8158 =  ( n5713 ) | ( n5722 )  ;
assign n8159 =  ( n8158 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8160 =  ( n8147 ) ? ( n8157 ) : ( n8159 ) ;
assign n8161 = ~ ( n8160 ) ;
assign n8162 =  ( n5909 ) | ( n8161 )  ;
assign n8163 = ~ ( n8162 ) ;
assign n8164 =  ( n8128 ) | ( n8163 )  ;
assign n8165 = ~ ( n8164 ) ;
assign n8166 =  ( n8127 ) | ( n8165 )  ;
assign n8167 =  ( n6825 ) | ( n6834 )  ;
assign n8168 =  ( n8167 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8169 =  ( n7455 ) ^ ( n8168 )  ;
assign n8170 =  ( n6483 ) | ( n6492 )  ;
assign n8171 =  ( n8170 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8172 =  ( n8169 ) ^ ( n8171 )  ;
assign n8173 =  ( n6030 ) | ( n6039 )  ;
assign n8174 =  ( n8173 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8175 =  ( n8172 ) ^ ( n8174 )  ;
assign n8176 =  ( n5802 ) | ( n5811 )  ;
assign n8177 =  ( n8176 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8178 =  ( n8175 ) ^ ( n8177 )  ;
assign n8179 = ~ ( n8178 ) ;
assign n8180 =  ( n8166 ) | ( n8179 )  ;
assign n8181 = ~ ( n8180 ) ;
assign n8182 = ~ ( n7845 ) ;
assign n8183 =  ( n8164 ) ^ ( n7455 )  ;
assign n8184 =  ( n6825 ) | ( n6834 )  ;
assign n8185 =  ( n8184 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8186 =  ( n8183 ) ^ ( n8185 )  ;
assign n8187 =  ( n6483 ) | ( n6492 )  ;
assign n8188 =  ( n8187 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8189 =  ( n8186 ) ^ ( n8188 )  ;
assign n8190 =  ( n6030 ) | ( n6039 )  ;
assign n8191 =  ( n8190 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8192 =  ( n8189 ) ^ ( n8191 )  ;
assign n8193 =  ( n5802 ) | ( n5811 )  ;
assign n8194 =  ( n8193 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8195 =  ( n8192 ) ^ ( n8194 )  ;
assign n8196 = ~ ( n8195 ) ;
assign n8197 =  ( n8182 ) | ( n8196 )  ;
assign n8198 = ~ ( n8197 ) ;
assign n8199 =  ( n8181 ) | ( n8198 )  ;
assign n8200 = ~ ( n7779 ) ;
assign n8201 =  ( n7784 ) | ( n6524 )  ;
assign n8202 = ~ ( n8201 ) ;
assign n8203 =  ( n8200 ) | ( n8202 )  ;
assign n8204 = ~ ( n7801 ) ;
assign n8205 =  ( n8203 ) | ( n8204 )  ;
assign n8206 = ~ ( n7809 ) ;
assign n8207 = ~ ( n6553 ) ;
assign n8208 =  ( n8206 ) | ( n8207 )  ;
assign n8209 =  ( n8205 ) ^ ( n8208 )  ;
assign n8210 =  ( n8209 ) ^ ( n8164 )  ;
assign n8211 =  ( n8210 ) ^ ( n7455 )  ;
assign n8212 =  ( n6825 ) | ( n6834 )  ;
assign n8213 =  ( n8212 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8214 =  ( n8211 ) ^ ( n8213 )  ;
assign n8215 =  ( n6483 ) | ( n6492 )  ;
assign n8216 =  ( n8215 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8217 =  ( n8214 ) ^ ( n8216 )  ;
assign n8218 =  ( n6030 ) | ( n6039 )  ;
assign n8219 =  ( n8218 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8220 =  ( n8217 ) ^ ( n8219 )  ;
assign n8221 =  ( n5802 ) | ( n5811 )  ;
assign n8222 =  ( n8221 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8223 =  ( n8220 ) ^ ( n8222 )  ;
assign n8224 = ~ ( n8223 ) ;
assign n8225 =  ( n8224 ) | ( n5879 )  ;
assign n8226 = ~ ( n8225 ) ;
assign n8227 =  ( n8199 ) | ( n8226 )  ;
assign n8228 = ~ ( n8227 ) ;
assign n8229 = ~ ( n7905 ) ;
assign n8230 = ~ ( n8164 ) ;
assign n8231 =  ( n8230 ) | ( n8179 )  ;
assign n8232 = ~ ( n8231 ) ;
assign n8233 =  ( n8229 ) | ( n8232 )  ;
assign n8234 = ~ ( n8233 ) ;
assign n8235 =  ( n8228 ) | ( n8234 )  ;
assign n8236 = ~ ( n8235 ) ;
assign n8237 =  ( n8227 ) ^ ( n8233 )  ;
assign n8238 = ~ ( n8237 ) ;
assign n8239 = ~ ( n7779 ) ;
assign n8240 =  ( n7784 ) | ( n6524 )  ;
assign n8241 = ~ ( n8240 ) ;
assign n8242 =  ( n8239 ) | ( n8241 )  ;
assign n8243 = ~ ( n7801 ) ;
assign n8244 =  ( n8242 ) | ( n8243 )  ;
assign n8245 = ~ ( n7809 ) ;
assign n8246 = ~ ( n6553 ) ;
assign n8247 =  ( n8245 ) | ( n8246 )  ;
assign n8248 =  ( n8244 ) ^ ( n8247 )  ;
assign n8249 = ~ ( n5902 ) ;
assign n8250 = ~ ( n5913 ) ;
assign n8251 =  ( n8249 ) | ( n8250 )  ;
assign n8252 =  ( n8248 ) ^ ( n8251 )  ;
assign n8253 = ~ ( n7455 ) ;
assign n8254 =  ( n8252 ) ^ ( n8253 )  ;
assign n8255 =  ( n6825 ) | ( n6834 )  ;
assign n8256 =  ( n8255 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8257 =  ( n8254 ) ^ ( n8256 )  ;
assign n8258 =  ( n6483 ) | ( n6492 )  ;
assign n8259 =  ( n8258 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8260 =  ( n8257 ) ^ ( n8259 )  ;
assign n8261 =  ( n6030 ) | ( n6039 )  ;
assign n8262 =  ( n8261 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8263 =  ( n8260 ) ^ ( n8262 )  ;
assign n8264 =  ( n5802 ) | ( n5811 )  ;
assign n8265 =  ( n8264 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8266 =  ( n8263 ) ^ ( n8265 )  ;
assign n8267 =  ( n5832 ) | ( n5841 )  ;
assign n8268 =  ( n8267 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8269 =  ( n8266 ) ^ ( n8268 )  ;
assign n8270 =  ( n5682 ) | ( n5691 )  ;
assign n8271 =  ( n8270 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8272 =  ( n8269 ) ^ ( n8271 )  ;
assign n8273 =  ( n5713 ) | ( n5722 )  ;
assign n8274 =  ( n8273 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8275 =  ( n8272 ) ^ ( n8274 )  ;
assign n8276 = ~ ( n8275 ) ;
assign n8277 =  ( n8238 ) | ( n8276 )  ;
assign n8278 = ~ ( n8277 ) ;
assign n8279 =  ( n8236 ) | ( n8278 )  ;
assign n8280 = ~ ( n8279 ) ;
assign n8281 =  ( bv_1_1_n5 ) ^ ( n7899 )  ;
assign n8282 = ~ ( n7905 ) ;
assign n8283 = ~ ( n7911 ) ;
assign n8284 =  ( n8282 ) | ( n8283 )  ;
assign n8285 =  ( n8281 ) ^ ( n8284 )  ;
assign n8286 = ~ ( n7467 ) ;
assign n8287 =  ( n7473 ) | ( n6524 )  ;
assign n8288 = ~ ( n8287 ) ;
assign n8289 =  ( n8286 ) | ( n8288 )  ;
assign n8290 = ~ ( n7491 ) ;
assign n8291 =  ( n8289 ) | ( n8290 )  ;
assign n8292 =  ( n8285 ) ^ ( n8291 )  ;
assign n8293 = ~ ( n7498 ) ;
assign n8294 = ~ ( n6553 ) ;
assign n8295 =  ( n8293 ) | ( n8294 )  ;
assign n8296 =  ( n8292 ) ^ ( n8295 )  ;
assign n8297 = ~ ( n5902 ) ;
assign n8298 = ~ ( n5913 ) ;
assign n8299 =  ( n8297 ) | ( n8298 )  ;
assign n8300 =  ( n8296 ) ^ ( n8299 )  ;
assign n8301 =  ( n6825 ) | ( n6834 )  ;
assign n8302 =  ( n8301 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8303 =  ( n8300 ) ^ ( n8302 )  ;
assign n8304 =  ( n6483 ) | ( n6492 )  ;
assign n8305 =  ( n8304 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8306 =  ( n8303 ) ^ ( n8305 )  ;
assign n8307 =  ( n6030 ) | ( n6039 )  ;
assign n8308 =  ( n8307 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8309 =  ( n8306 ) ^ ( n8308 )  ;
assign n8310 =  ( n5802 ) | ( n5811 )  ;
assign n8311 =  ( n8310 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8312 =  ( n8309 ) ^ ( n8311 )  ;
assign n8313 =  ( n5832 ) | ( n5841 )  ;
assign n8314 =  ( n8313 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8315 =  ( n8312 ) ^ ( n8314 )  ;
assign n8316 =  ( n5682 ) | ( n5691 )  ;
assign n8317 =  ( n8316 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8318 =  ( n8315 ) ^ ( n8317 )  ;
assign n8319 =  ( n5713 ) | ( n5722 )  ;
assign n8320 =  ( n8319 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8321 =  ( n8318 ) ^ ( n8320 )  ;
assign n8322 = ~ ( n8321 ) ;
assign n8323 =  ( n8280 ) | ( n8322 )  ;
assign n8324 =  ( n7961 ) ^ ( n7591 )  ;
assign n8325 = ~ ( n7597 ) ;
assign n8326 = ~ ( n7603 ) ;
assign n8327 =  ( n8325 ) | ( n8326 )  ;
assign n8328 =  ( n8324 ) ^ ( n8327 )  ;
assign n8329 = ~ ( n7133 ) ;
assign n8330 =  ( n7140 ) | ( n6337 )  ;
assign n8331 = ~ ( n8330 ) ;
assign n8332 =  ( n8329 ) | ( n8331 )  ;
assign n8333 = ~ ( n7159 ) ;
assign n8334 =  ( n8332 ) | ( n8333 )  ;
assign n8335 =  ( n8328 ) ^ ( n8334 )  ;
assign n8336 = ~ ( n7169 ) ;
assign n8337 = ~ ( n6366 ) ;
assign n8338 =  ( n8336 ) | ( n8337 )  ;
assign n8339 =  ( n8335 ) ^ ( n8338 )  ;
assign n8340 = ~ ( n5736 ) ;
assign n8341 =  ( n8340 ) | ( n5742 )  ;
assign n8342 =  ( n8339 ) ^ ( n8341 )  ;
assign n8343 =  ( n6825 ) | ( n6834 )  ;
assign n8344 =  ( n8343 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8345 = ~ ( n8344 ) ;
assign n8346 =  ( n8342 ) ^ ( n8345 )  ;
assign n8347 =  ( n6483 ) | ( n6492 )  ;
assign n8348 =  ( n8347 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8349 =  ( n8346 ) ^ ( n8348 )  ;
assign n8350 =  ( n6030 ) | ( n6039 )  ;
assign n8351 =  ( n8350 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8352 =  ( n8349 ) ^ ( n8351 )  ;
assign n8353 =  ( n5802 ) | ( n5811 )  ;
assign n8354 =  ( n8353 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8355 =  ( n8352 ) ^ ( n8354 )  ;
assign n8356 =  ( n5832 ) | ( n5841 )  ;
assign n8357 =  ( n8356 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8358 =  ( n8355 ) ^ ( n8357 )  ;
assign n8359 =  ( n5682 ) | ( n5691 )  ;
assign n8360 =  ( n8359 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8361 =  ( n8358 ) ^ ( n8360 )  ;
assign n8362 =  ( n5713 ) | ( n5722 )  ;
assign n8363 =  ( n8362 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8364 =  ( n8361 ) ^ ( n8363 )  ;
assign n8365 = ~ ( n8364 ) ;
assign n8366 =  ( n8323 ) | ( n8365 )  ;
assign n8367 = ~ ( n8366 ) ;
assign n8368 = ~ ( n8279 ) ;
assign n8369 = ~ ( n8321 ) ;
assign n8370 =  ( n8368 ) | ( n8369 )  ;
assign n8371 = ~ ( n8370 ) ;
assign n8372 =  ( n8371 ) ^ ( n7961 )  ;
assign n8373 =  ( n8372 ) ^ ( n7591 )  ;
assign n8374 = ~ ( n7597 ) ;
assign n8375 = ~ ( n7603 ) ;
assign n8376 =  ( n8374 ) | ( n8375 )  ;
assign n8377 =  ( n8373 ) ^ ( n8376 )  ;
assign n8378 = ~ ( n7133 ) ;
assign n8379 =  ( n7140 ) | ( n6337 )  ;
assign n8380 = ~ ( n8379 ) ;
assign n8381 =  ( n8378 ) | ( n8380 )  ;
assign n8382 = ~ ( n7159 ) ;
assign n8383 =  ( n8381 ) | ( n8382 )  ;
assign n8384 =  ( n8377 ) ^ ( n8383 )  ;
assign n8385 = ~ ( n7169 ) ;
assign n8386 = ~ ( n6366 ) ;
assign n8387 =  ( n8385 ) | ( n8386 )  ;
assign n8388 =  ( n8384 ) ^ ( n8387 )  ;
assign n8389 = ~ ( n5736 ) ;
assign n8390 =  ( n8389 ) | ( n5742 )  ;
assign n8391 =  ( n8388 ) ^ ( n8390 )  ;
assign n8392 =  ( n6825 ) | ( n6834 )  ;
assign n8393 =  ( n8392 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8394 = ~ ( n8393 ) ;
assign n8395 =  ( n8391 ) ^ ( n8394 )  ;
assign n8396 =  ( n6483 ) | ( n6492 )  ;
assign n8397 =  ( n8396 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8398 =  ( n8395 ) ^ ( n8397 )  ;
assign n8399 =  ( n6030 ) | ( n6039 )  ;
assign n8400 =  ( n8399 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8401 =  ( n8398 ) ^ ( n8400 )  ;
assign n8402 =  ( n5802 ) | ( n5811 )  ;
assign n8403 =  ( n8402 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8404 =  ( n8401 ) ^ ( n8403 )  ;
assign n8405 =  ( n5832 ) | ( n5841 )  ;
assign n8406 =  ( n8405 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8407 =  ( n8404 ) ^ ( n8406 )  ;
assign n8408 =  ( n5682 ) | ( n5691 )  ;
assign n8409 =  ( n8408 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8410 =  ( n8407 ) ^ ( n8409 )  ;
assign n8411 =  ( n5713 ) | ( n5722 )  ;
assign n8412 =  ( n8411 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8413 =  ( n8410 ) ^ ( n8412 )  ;
assign n8414 = ~ ( n8413 ) ;
assign n8415 = ~ ( n7809 ) ;
assign n8416 = ~ ( n6553 ) ;
assign n8417 =  ( n8415 ) | ( n8416 )  ;
assign n8418 = ~ ( n8417 ) ;
assign n8419 =  ( n7804 ) | ( n8418 )  ;
assign n8420 =  ( n8419 ) | ( n8179 )  ;
assign n8421 =  ( n5832 ) | ( n5841 )  ;
assign n8422 =  ( n8421 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8423 =  ( n5682 ) | ( n5691 )  ;
assign n8424 =  ( n8423 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8425 =  ( n8422 ) ^ ( n8424 )  ;
assign n8426 =  ( n8425 ) ^ ( n8160 )  ;
assign n8427 = ~ ( n8426 ) ;
assign n8428 =  ( n8420 ) | ( n8427 )  ;
assign n8429 = ~ ( n8428 ) ;
assign n8430 = ~ ( n7845 ) ;
assign n8431 =  ( n6825 ) | ( n6834 )  ;
assign n8432 =  ( n8431 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8433 =  ( n7455 ) ^ ( n8432 )  ;
assign n8434 =  ( n6483 ) | ( n6492 )  ;
assign n8435 =  ( n8434 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8436 =  ( n8433 ) ^ ( n8435 )  ;
assign n8437 =  ( n6030 ) | ( n6039 )  ;
assign n8438 =  ( n8437 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8439 =  ( n8436 ) ^ ( n8438 )  ;
assign n8440 =  ( n5802 ) | ( n5811 )  ;
assign n8441 =  ( n8440 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8442 =  ( n8439 ) ^ ( n8441 )  ;
assign n8443 =  ( n5832 ) | ( n5841 )  ;
assign n8444 =  ( n8443 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8445 =  ( n8442 ) ^ ( n8444 )  ;
assign n8446 =  ( n5682 ) | ( n5691 )  ;
assign n8447 =  ( n8446 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8448 =  ( n8445 ) ^ ( n8447 )  ;
assign n8449 =  ( n8448 ) ^ ( n8160 )  ;
assign n8450 = ~ ( n8449 ) ;
assign n8451 =  ( n8430 ) | ( n8450 )  ;
assign n8452 = ~ ( n8451 ) ;
assign n8453 =  ( n8429 ) | ( n8452 )  ;
assign n8454 = ~ ( n7779 ) ;
assign n8455 =  ( n7784 ) | ( n6524 )  ;
assign n8456 = ~ ( n8455 ) ;
assign n8457 =  ( n8454 ) | ( n8456 )  ;
assign n8458 = ~ ( n7801 ) ;
assign n8459 =  ( n8457 ) | ( n8458 )  ;
assign n8460 = ~ ( n7809 ) ;
assign n8461 = ~ ( n6553 ) ;
assign n8462 =  ( n8460 ) | ( n8461 )  ;
assign n8463 =  ( n8459 ) ^ ( n8462 )  ;
assign n8464 =  ( n8463 ) ^ ( n7455 )  ;
assign n8465 =  ( n6825 ) | ( n6834 )  ;
assign n8466 =  ( n8465 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8467 =  ( n8464 ) ^ ( n8466 )  ;
assign n8468 =  ( n6483 ) | ( n6492 )  ;
assign n8469 =  ( n8468 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8470 =  ( n8467 ) ^ ( n8469 )  ;
assign n8471 =  ( n6030 ) | ( n6039 )  ;
assign n8472 =  ( n8471 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8473 =  ( n8470 ) ^ ( n8472 )  ;
assign n8474 =  ( n5802 ) | ( n5811 )  ;
assign n8475 =  ( n8474 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8476 =  ( n8473 ) ^ ( n8475 )  ;
assign n8477 =  ( n5832 ) | ( n5841 )  ;
assign n8478 =  ( n8477 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8479 =  ( n8476 ) ^ ( n8478 )  ;
assign n8480 =  ( n5682 ) | ( n5691 )  ;
assign n8481 =  ( n8480 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8482 =  ( n8479 ) ^ ( n8481 )  ;
assign n8483 =  ( n8482 ) ^ ( n8160 )  ;
assign n8484 = ~ ( n8483 ) ;
assign n8485 = kd[15:15] ;
assign n8486 = ~ ( n8485 ) ;
assign n8487 =  ( n8484 ) | ( n8486 )  ;
assign n8488 =  ( n8487 ) | ( n8155 )  ;
assign n8489 = ~ ( n8488 ) ;
assign n8490 =  ( n8453 ) | ( n8489 )  ;
assign n8491 = ~ ( n8490 ) ;
assign n8492 = ~ ( n7905 ) ;
assign n8493 =  ( n8179 ) | ( n8427 )  ;
assign n8494 = ~ ( n8493 ) ;
assign n8495 =  ( n8492 ) | ( n8494 )  ;
assign n8496 = ~ ( n8495 ) ;
assign n8497 =  ( n8491 ) | ( n8496 )  ;
assign n8498 = ~ ( n8497 ) ;
assign n8499 = ~ ( n7905 ) ;
assign n8500 =  ( n8179 ) | ( n8427 )  ;
assign n8501 = ~ ( n8500 ) ;
assign n8502 =  ( n8499 ) | ( n8501 )  ;
assign n8503 =  ( n8490 ) ^ ( n8502 )  ;
assign n8504 = ~ ( n8503 ) ;
assign n8505 = ~ ( n7779 ) ;
assign n8506 =  ( n7784 ) | ( n6524 )  ;
assign n8507 = ~ ( n8506 ) ;
assign n8508 =  ( n8505 ) | ( n8507 )  ;
assign n8509 = ~ ( n7801 ) ;
assign n8510 =  ( n8508 ) | ( n8509 )  ;
assign n8511 = ~ ( n7809 ) ;
assign n8512 = ~ ( n6553 ) ;
assign n8513 =  ( n8511 ) | ( n8512 )  ;
assign n8514 =  ( n8510 ) ^ ( n8513 )  ;
assign n8515 =  ( n8514 ) ^ ( n8164 )  ;
assign n8516 =  ( n8515 ) ^ ( n7455 )  ;
assign n8517 =  ( n6825 ) | ( n6834 )  ;
assign n8518 =  ( n8517 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8519 =  ( n8516 ) ^ ( n8518 )  ;
assign n8520 =  ( n6483 ) | ( n6492 )  ;
assign n8521 =  ( n8520 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8522 =  ( n8519 ) ^ ( n8521 )  ;
assign n8523 =  ( n6030 ) | ( n6039 )  ;
assign n8524 =  ( n8523 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8525 =  ( n8522 ) ^ ( n8524 )  ;
assign n8526 =  ( n5802 ) | ( n5811 )  ;
assign n8527 =  ( n8526 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8528 =  ( n8525 ) ^ ( n8527 )  ;
assign n8529 =  ( n5832 ) | ( n5841 )  ;
assign n8530 =  ( n8529 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8531 =  ( n8528 ) ^ ( n8530 )  ;
assign n8532 =  ( n5682 ) | ( n5691 )  ;
assign n8533 =  ( n8532 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8534 =  ( n8531 ) ^ ( n8533 )  ;
assign n8535 =  ( n5713 ) | ( n5722 )  ;
assign n8536 =  ( n8535 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8537 =  ( n8534 ) ^ ( n8536 )  ;
assign n8538 = ~ ( n8537 ) ;
assign n8539 =  ( n8504 ) | ( n8538 )  ;
assign n8540 = ~ ( n8539 ) ;
assign n8541 =  ( n8498 ) | ( n8540 )  ;
assign n8542 = ~ ( n8541 ) ;
assign n8543 =  ( n8227 ) ^ ( n8233 )  ;
assign n8544 = ~ ( n7779 ) ;
assign n8545 =  ( n7784 ) | ( n6524 )  ;
assign n8546 = ~ ( n8545 ) ;
assign n8547 =  ( n8544 ) | ( n8546 )  ;
assign n8548 = ~ ( n7801 ) ;
assign n8549 =  ( n8547 ) | ( n8548 )  ;
assign n8550 =  ( n8543 ) ^ ( n8549 )  ;
assign n8551 = ~ ( n7809 ) ;
assign n8552 = ~ ( n6553 ) ;
assign n8553 =  ( n8551 ) | ( n8552 )  ;
assign n8554 =  ( n8550 ) ^ ( n8553 )  ;
assign n8555 = ~ ( n5902 ) ;
assign n8556 = ~ ( n5913 ) ;
assign n8557 =  ( n8555 ) | ( n8556 )  ;
assign n8558 =  ( n8554 ) ^ ( n8557 )  ;
assign n8559 = ~ ( n7455 ) ;
assign n8560 =  ( n8558 ) ^ ( n8559 )  ;
assign n8561 =  ( n6825 ) | ( n6834 )  ;
assign n8562 =  ( n8561 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8563 =  ( n8560 ) ^ ( n8562 )  ;
assign n8564 =  ( n6483 ) | ( n6492 )  ;
assign n8565 =  ( n8564 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8566 =  ( n8563 ) ^ ( n8565 )  ;
assign n8567 =  ( n6030 ) | ( n6039 )  ;
assign n8568 =  ( n8567 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8569 =  ( n8566 ) ^ ( n8568 )  ;
assign n8570 =  ( n5802 ) | ( n5811 )  ;
assign n8571 =  ( n8570 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8572 =  ( n8569 ) ^ ( n8571 )  ;
assign n8573 =  ( n5832 ) | ( n5841 )  ;
assign n8574 =  ( n8573 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8575 =  ( n8572 ) ^ ( n8574 )  ;
assign n8576 =  ( n5682 ) | ( n5691 )  ;
assign n8577 =  ( n8576 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8578 =  ( n8575 ) ^ ( n8577 )  ;
assign n8579 =  ( n5713 ) | ( n5722 )  ;
assign n8580 =  ( n8579 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8581 =  ( n8578 ) ^ ( n8580 )  ;
assign n8582 = ~ ( n8581 ) ;
assign n8583 =  ( n8542 ) | ( n8582 )  ;
assign n8584 = ~ ( n8583 ) ;
assign n8585 =  ( n8541 ) ^ ( n8227 )  ;
assign n8586 =  ( n8585 ) ^ ( n8233 )  ;
assign n8587 = ~ ( n7779 ) ;
assign n8588 =  ( n7784 ) | ( n6524 )  ;
assign n8589 = ~ ( n8588 ) ;
assign n8590 =  ( n8587 ) | ( n8589 )  ;
assign n8591 = ~ ( n7801 ) ;
assign n8592 =  ( n8590 ) | ( n8591 )  ;
assign n8593 =  ( n8586 ) ^ ( n8592 )  ;
assign n8594 = ~ ( n7809 ) ;
assign n8595 = ~ ( n6553 ) ;
assign n8596 =  ( n8594 ) | ( n8595 )  ;
assign n8597 =  ( n8593 ) ^ ( n8596 )  ;
assign n8598 = ~ ( n5902 ) ;
assign n8599 = ~ ( n5913 ) ;
assign n8600 =  ( n8598 ) | ( n8599 )  ;
assign n8601 =  ( n8597 ) ^ ( n8600 )  ;
assign n8602 = ~ ( n7455 ) ;
assign n8603 =  ( n8601 ) ^ ( n8602 )  ;
assign n8604 =  ( n6825 ) | ( n6834 )  ;
assign n8605 =  ( n8604 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8606 =  ( n8603 ) ^ ( n8605 )  ;
assign n8607 =  ( n6483 ) | ( n6492 )  ;
assign n8608 =  ( n8607 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8609 =  ( n8606 ) ^ ( n8608 )  ;
assign n8610 =  ( n6030 ) | ( n6039 )  ;
assign n8611 =  ( n8610 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8612 =  ( n8609 ) ^ ( n8611 )  ;
assign n8613 =  ( n5802 ) | ( n5811 )  ;
assign n8614 =  ( n8613 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8615 =  ( n8612 ) ^ ( n8614 )  ;
assign n8616 =  ( n5832 ) | ( n5841 )  ;
assign n8617 =  ( n8616 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8618 =  ( n8615 ) ^ ( n8617 )  ;
assign n8619 =  ( n5682 ) | ( n5691 )  ;
assign n8620 =  ( n8619 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8621 =  ( n8618 ) ^ ( n8620 )  ;
assign n8622 =  ( n5713 ) | ( n5722 )  ;
assign n8623 =  ( n8622 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8624 =  ( n8621 ) ^ ( n8623 )  ;
assign n8625 =  ( n8584 ) | ( n8624 )  ;
assign n8626 = ~ ( n8625 ) ;
assign n8627 =  ( n8414 ) | ( n8626 )  ;
assign n8628 =  ( bv_1_1_n5 ) ^ ( n8279 )  ;
assign n8629 =  ( n8628 ) ^ ( n7899 )  ;
assign n8630 = ~ ( n7905 ) ;
assign n8631 = ~ ( n7911 ) ;
assign n8632 =  ( n8630 ) | ( n8631 )  ;
assign n8633 =  ( n8629 ) ^ ( n8632 )  ;
assign n8634 = ~ ( n7467 ) ;
assign n8635 =  ( n7473 ) | ( n6524 )  ;
assign n8636 = ~ ( n8635 ) ;
assign n8637 =  ( n8634 ) | ( n8636 )  ;
assign n8638 = ~ ( n7491 ) ;
assign n8639 =  ( n8637 ) | ( n8638 )  ;
assign n8640 =  ( n8633 ) ^ ( n8639 )  ;
assign n8641 = ~ ( n7498 ) ;
assign n8642 = ~ ( n6553 ) ;
assign n8643 =  ( n8641 ) | ( n8642 )  ;
assign n8644 =  ( n8640 ) ^ ( n8643 )  ;
assign n8645 = ~ ( n5902 ) ;
assign n8646 = ~ ( n5913 ) ;
assign n8647 =  ( n8645 ) | ( n8646 )  ;
assign n8648 =  ( n8644 ) ^ ( n8647 )  ;
assign n8649 =  ( n6825 ) | ( n6834 )  ;
assign n8650 =  ( n8649 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8651 =  ( n8648 ) ^ ( n8650 )  ;
assign n8652 =  ( n6483 ) | ( n6492 )  ;
assign n8653 =  ( n8652 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8654 =  ( n8651 ) ^ ( n8653 )  ;
assign n8655 =  ( n6030 ) | ( n6039 )  ;
assign n8656 =  ( n8655 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8657 =  ( n8654 ) ^ ( n8656 )  ;
assign n8658 =  ( n5802 ) | ( n5811 )  ;
assign n8659 =  ( n8658 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8660 =  ( n8657 ) ^ ( n8659 )  ;
assign n8661 =  ( n5832 ) | ( n5841 )  ;
assign n8662 =  ( n8661 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8663 =  ( n8660 ) ^ ( n8662 )  ;
assign n8664 =  ( n5682 ) | ( n5691 )  ;
assign n8665 =  ( n8664 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8666 =  ( n8663 ) ^ ( n8665 )  ;
assign n8667 =  ( n5713 ) | ( n5722 )  ;
assign n8668 =  ( n8667 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8669 =  ( n8666 ) ^ ( n8668 )  ;
assign n8670 = ~ ( n8669 ) ;
assign n8671 =  ( n8627 ) | ( n8670 )  ;
assign n8672 = ~ ( n8671 ) ;
assign n8673 =  ( n8367 ) | ( n8672 )  ;
assign n8674 = ~ ( n8413 ) ;
assign n8675 =  ( bv_1_1_n5 ) ^ ( n8625 )  ;
assign n8676 =  ( n8675 ) ^ ( n8279 )  ;
assign n8677 =  ( n8676 ) ^ ( n7899 )  ;
assign n8678 = ~ ( n7905 ) ;
assign n8679 = ~ ( n7911 ) ;
assign n8680 =  ( n8678 ) | ( n8679 )  ;
assign n8681 =  ( n8677 ) ^ ( n8680 )  ;
assign n8682 = ~ ( n7467 ) ;
assign n8683 =  ( n7473 ) | ( n6524 )  ;
assign n8684 = ~ ( n8683 ) ;
assign n8685 =  ( n8682 ) | ( n8684 )  ;
assign n8686 = ~ ( n7491 ) ;
assign n8687 =  ( n8685 ) | ( n8686 )  ;
assign n8688 =  ( n8681 ) ^ ( n8687 )  ;
assign n8689 = ~ ( n7498 ) ;
assign n8690 = ~ ( n6553 ) ;
assign n8691 =  ( n8689 ) | ( n8690 )  ;
assign n8692 =  ( n8688 ) ^ ( n8691 )  ;
assign n8693 = ~ ( n5902 ) ;
assign n8694 = ~ ( n5913 ) ;
assign n8695 =  ( n8693 ) | ( n8694 )  ;
assign n8696 =  ( n8692 ) ^ ( n8695 )  ;
assign n8697 =  ( n6825 ) | ( n6834 )  ;
assign n8698 =  ( n8697 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8699 =  ( n8696 ) ^ ( n8698 )  ;
assign n8700 =  ( n6483 ) | ( n6492 )  ;
assign n8701 =  ( n8700 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8702 =  ( n8699 ) ^ ( n8701 )  ;
assign n8703 =  ( n6030 ) | ( n6039 )  ;
assign n8704 =  ( n8703 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8705 =  ( n8702 ) ^ ( n8704 )  ;
assign n8706 =  ( n5802 ) | ( n5811 )  ;
assign n8707 =  ( n8706 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8708 =  ( n8705 ) ^ ( n8707 )  ;
assign n8709 =  ( n5832 ) | ( n5841 )  ;
assign n8710 =  ( n8709 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8711 =  ( n8708 ) ^ ( n8710 )  ;
assign n8712 =  ( n5682 ) | ( n5691 )  ;
assign n8713 =  ( n8712 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8714 =  ( n8711 ) ^ ( n8713 )  ;
assign n8715 =  ( n5713 ) | ( n5722 )  ;
assign n8716 =  ( n8715 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8717 =  ( n8714 ) ^ ( n8716 )  ;
assign n8718 = ~ ( n8717 ) ;
assign n8719 =  ( n8674 ) | ( n8718 )  ;
assign n8720 = ~ ( n7809 ) ;
assign n8721 = ~ ( n6553 ) ;
assign n8722 =  ( n8720 ) | ( n8721 )  ;
assign n8723 = ~ ( n8722 ) ;
assign n8724 =  ( n7804 ) | ( n8723 )  ;
assign n8725 =  ( n5832 ) | ( n5841 )  ;
assign n8726 =  ( n8725 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8727 = ~ ( n8726 ) ;
assign n8728 = kd[13:13] ;
assign n8729 =  ( n8728 ) == ( bv_1_0_n2 )  ;
assign n8730 = kd[12:12] ;
assign n8731 =  ( n8730 ) == ( bv_1_1_n5 )  ;
assign n8732 =  ( n8729 ) | ( n8731 )  ;
assign n8733 = kd[11:11] ;
assign n8734 =  ( n8733 ) == ( bv_1_1_n5 )  ;
assign n8735 =  ( n8732 ) | ( n8734 )  ;
assign n8736 = ~ ( n8735 )  ;
assign n8737 = kd[13:13] ;
assign n8738 =  ( n8737 ) == ( bv_1_1_n5 )  ;
assign n8739 = kd[12:12] ;
assign n8740 =  ( n8739 ) == ( bv_1_0_n2 )  ;
assign n8741 =  ( n8738 ) | ( n8740 )  ;
assign n8742 = kd[11:11] ;
assign n8743 =  ( n8742 ) == ( bv_1_0_n2 )  ;
assign n8744 =  ( n8741 ) | ( n8743 )  ;
assign n8745 = ~ ( n8744 )  ;
assign n8746 =  ( n8736 ) | ( n8745 )  ;
assign n8747 = kd[13:13] ;
assign n8748 = ~ ( n8747 ) ;
assign n8749 = kd[12:12] ;
assign n8750 = ~ ( n8749 ) ;
assign n8751 = kd[11:11] ;
assign n8752 = ~ ( n8751 ) ;
assign n8753 =  ( n8750 ) | ( n8752 )  ;
assign n8754 = ~ ( n8753 ) ;
assign n8755 =  ( n8748 ) | ( n8754 )  ;
assign n8756 = ~ ( n8755 ) ;
assign n8757 =  ( n5682 ) | ( n5691 )  ;
assign n8758 =  ( n8757 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8759 =  ( n8746 ) ? ( n8756 ) : ( n8758 ) ;
assign n8760 = ~ ( n8759 ) ;
assign n8761 =  ( n8727 ) | ( n8760 )  ;
assign n8762 = ~ ( n8761 ) ;
assign n8763 =  ( n5832 ) | ( n5841 )  ;
assign n8764 =  ( n8763 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8765 =  ( n8764 ) ^ ( n8759 )  ;
assign n8766 = ~ ( n8765 ) ;
assign n8767 = kd[13:13] ;
assign n8768 = ~ ( n8767 ) ;
assign n8769 =  ( n8766 ) | ( n8768 )  ;
assign n8770 =  ( n8769 ) | ( n8754 )  ;
assign n8771 = ~ ( n8770 ) ;
assign n8772 =  ( n8762 ) | ( n8771 )  ;
assign n8773 = ~ ( n8772 ) ;
assign n8774 =  ( n8724 ) | ( n8773 )  ;
assign n8775 =  ( n8774 ) | ( n8179 )  ;
assign n8776 = ~ ( n8775 ) ;
assign n8777 = ~ ( n7845 ) ;
assign n8778 = ~ ( n8761 ) ;
assign n8779 =  ( n8778 ) | ( n8771 )  ;
assign n8780 =  ( n8779 ) ^ ( n7455 )  ;
assign n8781 =  ( n6825 ) | ( n6834 )  ;
assign n8782 =  ( n8781 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8783 =  ( n8780 ) ^ ( n8782 )  ;
assign n8784 =  ( n6483 ) | ( n6492 )  ;
assign n8785 =  ( n8784 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8786 =  ( n8783 ) ^ ( n8785 )  ;
assign n8787 =  ( n6030 ) | ( n6039 )  ;
assign n8788 =  ( n8787 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8789 =  ( n8786 ) ^ ( n8788 )  ;
assign n8790 =  ( n5802 ) | ( n5811 )  ;
assign n8791 =  ( n8790 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8792 =  ( n8789 ) ^ ( n8791 )  ;
assign n8793 = ~ ( n8792 ) ;
assign n8794 =  ( n8777 ) | ( n8793 )  ;
assign n8795 = ~ ( n8794 ) ;
assign n8796 =  ( n8776 ) | ( n8795 )  ;
assign n8797 = ~ ( n7779 ) ;
assign n8798 =  ( n7784 ) | ( n6524 )  ;
assign n8799 = ~ ( n8798 ) ;
assign n8800 =  ( n8797 ) | ( n8799 )  ;
assign n8801 = ~ ( n7801 ) ;
assign n8802 =  ( n8800 ) | ( n8801 )  ;
assign n8803 = ~ ( n7809 ) ;
assign n8804 = ~ ( n6553 ) ;
assign n8805 =  ( n8803 ) | ( n8804 )  ;
assign n8806 =  ( n8802 ) ^ ( n8805 )  ;
assign n8807 = ~ ( n8761 ) ;
assign n8808 =  ( n8807 ) | ( n8771 )  ;
assign n8809 =  ( n8806 ) ^ ( n8808 )  ;
assign n8810 =  ( n8809 ) ^ ( n7455 )  ;
assign n8811 =  ( n6825 ) | ( n6834 )  ;
assign n8812 =  ( n8811 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8813 =  ( n8810 ) ^ ( n8812 )  ;
assign n8814 =  ( n6483 ) | ( n6492 )  ;
assign n8815 =  ( n8814 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8816 =  ( n8813 ) ^ ( n8815 )  ;
assign n8817 =  ( n6030 ) | ( n6039 )  ;
assign n8818 =  ( n8817 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8819 =  ( n8816 ) ^ ( n8818 )  ;
assign n8820 =  ( n5802 ) | ( n5811 )  ;
assign n8821 =  ( n8820 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8822 =  ( n8819 ) ^ ( n8821 )  ;
assign n8823 = ~ ( n8822 ) ;
assign n8824 =  ( n5832 ) | ( n5841 )  ;
assign n8825 =  ( n8824 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8826 = ~ ( n8825 ) ;
assign n8827 =  ( n8823 ) | ( n8826 )  ;
assign n8828 = ~ ( n8827 ) ;
assign n8829 =  ( n8796 ) | ( n8828 )  ;
assign n8830 = ~ ( n8829 ) ;
assign n8831 = ~ ( n7905 ) ;
assign n8832 = ~ ( n8761 ) ;
assign n8833 =  ( n8832 ) | ( n8771 )  ;
assign n8834 = ~ ( n8833 ) ;
assign n8835 =  ( n8834 ) | ( n8179 )  ;
assign n8836 = ~ ( n8835 ) ;
assign n8837 =  ( n8831 ) | ( n8836 )  ;
assign n8838 = ~ ( n8837 ) ;
assign n8839 =  ( n8830 ) | ( n8838 )  ;
assign n8840 = ~ ( n8839 ) ;
assign n8841 = ~ ( n7905 ) ;
assign n8842 = ~ ( n8835 ) ;
assign n8843 =  ( n8841 ) | ( n8842 )  ;
assign n8844 =  ( n8829 ) ^ ( n8843 )  ;
assign n8845 = ~ ( n8844 ) ;
assign n8846 = ~ ( n7779 ) ;
assign n8847 =  ( n7784 ) | ( n6524 )  ;
assign n8848 = ~ ( n8847 ) ;
assign n8849 =  ( n8846 ) | ( n8848 )  ;
assign n8850 = ~ ( n7801 ) ;
assign n8851 =  ( n8849 ) | ( n8850 )  ;
assign n8852 = ~ ( n7809 ) ;
assign n8853 = ~ ( n6553 ) ;
assign n8854 =  ( n8852 ) | ( n8853 )  ;
assign n8855 =  ( n8851 ) ^ ( n8854 )  ;
assign n8856 =  ( n8855 ) ^ ( n7455 )  ;
assign n8857 =  ( n6825 ) | ( n6834 )  ;
assign n8858 =  ( n8857 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8859 =  ( n8856 ) ^ ( n8858 )  ;
assign n8860 =  ( n6483 ) | ( n6492 )  ;
assign n8861 =  ( n8860 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8862 =  ( n8859 ) ^ ( n8861 )  ;
assign n8863 =  ( n6030 ) | ( n6039 )  ;
assign n8864 =  ( n8863 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8865 =  ( n8862 ) ^ ( n8864 )  ;
assign n8866 =  ( n5802 ) | ( n5811 )  ;
assign n8867 =  ( n8866 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8868 =  ( n8865 ) ^ ( n8867 )  ;
assign n8869 =  ( n5832 ) | ( n5841 )  ;
assign n8870 =  ( n8869 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8871 =  ( n8868 ) ^ ( n8870 )  ;
assign n8872 =  ( n5682 ) | ( n5691 )  ;
assign n8873 =  ( n8872 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8874 =  ( n8871 ) ^ ( n8873 )  ;
assign n8875 =  ( n8874 ) ^ ( n8160 )  ;
assign n8876 =  ( n8875 ) ^ ( n8157 )  ;
assign n8877 = ~ ( n8876 ) ;
assign n8878 =  ( n8845 ) | ( n8877 )  ;
assign n8879 = ~ ( n8878 ) ;
assign n8880 =  ( n8840 ) | ( n8879 )  ;
assign n8881 = ~ ( n8880 ) ;
assign n8882 = ~ ( n7905 ) ;
assign n8883 =  ( n8179 ) | ( n8427 )  ;
assign n8884 = ~ ( n8883 ) ;
assign n8885 =  ( n8882 ) | ( n8884 )  ;
assign n8886 =  ( n8490 ) ^ ( n8885 )  ;
assign n8887 = ~ ( n7779 ) ;
assign n8888 =  ( n7784 ) | ( n6524 )  ;
assign n8889 = ~ ( n8888 ) ;
assign n8890 =  ( n8887 ) | ( n8889 )  ;
assign n8891 = ~ ( n7801 ) ;
assign n8892 =  ( n8890 ) | ( n8891 )  ;
assign n8893 =  ( n8886 ) ^ ( n8892 )  ;
assign n8894 = ~ ( n7809 ) ;
assign n8895 = ~ ( n6553 ) ;
assign n8896 =  ( n8894 ) | ( n8895 )  ;
assign n8897 =  ( n8893 ) ^ ( n8896 )  ;
assign n8898 =  ( n8897 ) ^ ( n8164 )  ;
assign n8899 =  ( n8898 ) ^ ( n7455 )  ;
assign n8900 =  ( n6825 ) | ( n6834 )  ;
assign n8901 =  ( n8900 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8902 =  ( n8899 ) ^ ( n8901 )  ;
assign n8903 =  ( n6483 ) | ( n6492 )  ;
assign n8904 =  ( n8903 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8905 =  ( n8902 ) ^ ( n8904 )  ;
assign n8906 =  ( n6030 ) | ( n6039 )  ;
assign n8907 =  ( n8906 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8908 =  ( n8905 ) ^ ( n8907 )  ;
assign n8909 =  ( n5802 ) | ( n5811 )  ;
assign n8910 =  ( n8909 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8911 =  ( n8908 ) ^ ( n8910 )  ;
assign n8912 =  ( n5832 ) | ( n5841 )  ;
assign n8913 =  ( n8912 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8914 =  ( n8911 ) ^ ( n8913 )  ;
assign n8915 =  ( n5682 ) | ( n5691 )  ;
assign n8916 =  ( n8915 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8917 =  ( n8914 ) ^ ( n8916 )  ;
assign n8918 =  ( n5713 ) | ( n5722 )  ;
assign n8919 =  ( n8918 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8920 =  ( n8917 ) ^ ( n8919 )  ;
assign n8921 = ~ ( n8920 ) ;
assign n8922 =  ( n8881 ) | ( n8921 )  ;
assign n8923 =  ( bv_1_1_n5 ) ^ ( n8541 )  ;
assign n8924 =  ( n8923 ) ^ ( n8227 )  ;
assign n8925 =  ( n8924 ) ^ ( n8233 )  ;
assign n8926 = ~ ( n7779 ) ;
assign n8927 =  ( n7784 ) | ( n6524 )  ;
assign n8928 = ~ ( n8927 ) ;
assign n8929 =  ( n8926 ) | ( n8928 )  ;
assign n8930 = ~ ( n7801 ) ;
assign n8931 =  ( n8929 ) | ( n8930 )  ;
assign n8932 =  ( n8925 ) ^ ( n8931 )  ;
assign n8933 = ~ ( n7809 ) ;
assign n8934 = ~ ( n6553 ) ;
assign n8935 =  ( n8933 ) | ( n8934 )  ;
assign n8936 =  ( n8932 ) ^ ( n8935 )  ;
assign n8937 = ~ ( n5902 ) ;
assign n8938 = ~ ( n5913 ) ;
assign n8939 =  ( n8937 ) | ( n8938 )  ;
assign n8940 =  ( n8936 ) ^ ( n8939 )  ;
assign n8941 = ~ ( n7455 ) ;
assign n8942 =  ( n8940 ) ^ ( n8941 )  ;
assign n8943 =  ( n6825 ) | ( n6834 )  ;
assign n8944 =  ( n8943 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8945 =  ( n8942 ) ^ ( n8944 )  ;
assign n8946 =  ( n6483 ) | ( n6492 )  ;
assign n8947 =  ( n8946 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8948 =  ( n8945 ) ^ ( n8947 )  ;
assign n8949 =  ( n6030 ) | ( n6039 )  ;
assign n8950 =  ( n8949 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n8951 =  ( n8948 ) ^ ( n8950 )  ;
assign n8952 =  ( n5802 ) | ( n5811 )  ;
assign n8953 =  ( n8952 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n8954 =  ( n8951 ) ^ ( n8953 )  ;
assign n8955 =  ( n5832 ) | ( n5841 )  ;
assign n8956 =  ( n8955 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n8957 =  ( n8954 ) ^ ( n8956 )  ;
assign n8958 =  ( n5682 ) | ( n5691 )  ;
assign n8959 =  ( n8958 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n8960 =  ( n8957 ) ^ ( n8959 )  ;
assign n8961 =  ( n5713 ) | ( n5722 )  ;
assign n8962 =  ( n8961 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n8963 =  ( n8960 ) ^ ( n8962 )  ;
assign n8964 = ~ ( n8963 ) ;
assign n8965 =  ( n8922 ) | ( n8964 )  ;
assign n8966 = ~ ( n8965 ) ;
assign n8967 = ~ ( n8880 ) ;
assign n8968 = ~ ( n8920 ) ;
assign n8969 =  ( n8967 ) | ( n8968 )  ;
assign n8970 = ~ ( n8969 ) ;
assign n8971 =  ( bv_1_1_n5 ) ^ ( n8970 )  ;
assign n8972 =  ( n8971 ) ^ ( n8541 )  ;
assign n8973 =  ( n8972 ) ^ ( n8227 )  ;
assign n8974 =  ( n8973 ) ^ ( n8233 )  ;
assign n8975 = ~ ( n7779 ) ;
assign n8976 =  ( n7784 ) | ( n6524 )  ;
assign n8977 = ~ ( n8976 ) ;
assign n8978 =  ( n8975 ) | ( n8977 )  ;
assign n8979 = ~ ( n7801 ) ;
assign n8980 =  ( n8978 ) | ( n8979 )  ;
assign n8981 =  ( n8974 ) ^ ( n8980 )  ;
assign n8982 = ~ ( n7809 ) ;
assign n8983 = ~ ( n6553 ) ;
assign n8984 =  ( n8982 ) | ( n8983 )  ;
assign n8985 =  ( n8981 ) ^ ( n8984 )  ;
assign n8986 = ~ ( n5902 ) ;
assign n8987 = ~ ( n5913 ) ;
assign n8988 =  ( n8986 ) | ( n8987 )  ;
assign n8989 =  ( n8985 ) ^ ( n8988 )  ;
assign n8990 = ~ ( n7455 ) ;
assign n8991 =  ( n8989 ) ^ ( n8990 )  ;
assign n8992 =  ( n6825 ) | ( n6834 )  ;
assign n8993 =  ( n8992 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n8994 =  ( n8991 ) ^ ( n8993 )  ;
assign n8995 =  ( n6483 ) | ( n6492 )  ;
assign n8996 =  ( n8995 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n8997 =  ( n8994 ) ^ ( n8996 )  ;
assign n8998 =  ( n6030 ) | ( n6039 )  ;
assign n8999 =  ( n8998 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9000 =  ( n8997 ) ^ ( n8999 )  ;
assign n9001 =  ( n5802 ) | ( n5811 )  ;
assign n9002 =  ( n9001 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9003 =  ( n9000 ) ^ ( n9002 )  ;
assign n9004 =  ( n5832 ) | ( n5841 )  ;
assign n9005 =  ( n9004 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9006 =  ( n9003 ) ^ ( n9005 )  ;
assign n9007 =  ( n5682 ) | ( n5691 )  ;
assign n9008 =  ( n9007 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9009 =  ( n9006 ) ^ ( n9008 )  ;
assign n9010 =  ( n5713 ) | ( n5722 )  ;
assign n9011 =  ( n9010 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n9012 =  ( n9009 ) ^ ( n9011 )  ;
assign n9013 = ~ ( n9012 ) ;
assign n9014 = ~ ( n7905 ) ;
assign n9015 = ~ ( n7845 ) ;
assign n9016 =  ( n9015 ) | ( n8179 )  ;
assign n9017 = ~ ( n9016 ) ;
assign n9018 =  ( n9014 ) | ( n9017 )  ;
assign n9019 = ~ ( n9018 ) ;
assign n9020 = ~ ( n7779 ) ;
assign n9021 =  ( n7784 ) | ( n6524 )  ;
assign n9022 = ~ ( n9021 ) ;
assign n9023 =  ( n9020 ) | ( n9022 )  ;
assign n9024 = ~ ( n7801 ) ;
assign n9025 =  ( n9023 ) | ( n9024 )  ;
assign n9026 = ~ ( n7809 ) ;
assign n9027 = ~ ( n6553 ) ;
assign n9028 =  ( n9026 ) | ( n9027 )  ;
assign n9029 =  ( n9025 ) ^ ( n9028 )  ;
assign n9030 = ~ ( n8761 ) ;
assign n9031 =  ( n9030 ) | ( n8771 )  ;
assign n9032 =  ( n9029 ) ^ ( n9031 )  ;
assign n9033 =  ( n9032 ) ^ ( n7455 )  ;
assign n9034 =  ( n6825 ) | ( n6834 )  ;
assign n9035 =  ( n9034 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9036 =  ( n9033 ) ^ ( n9035 )  ;
assign n9037 =  ( n6483 ) | ( n6492 )  ;
assign n9038 =  ( n9037 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9039 =  ( n9036 ) ^ ( n9038 )  ;
assign n9040 =  ( n6030 ) | ( n6039 )  ;
assign n9041 =  ( n9040 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9042 =  ( n9039 ) ^ ( n9041 )  ;
assign n9043 =  ( n5802 ) | ( n5811 )  ;
assign n9044 =  ( n9043 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9045 =  ( n9042 ) ^ ( n9044 )  ;
assign n9046 =  ( n5832 ) | ( n5841 )  ;
assign n9047 =  ( n9046 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9048 =  ( n9045 ) ^ ( n9047 )  ;
assign n9049 = ~ ( n9048 ) ;
assign n9050 =  ( n9019 ) | ( n9049 )  ;
assign n9051 = ~ ( n9050 ) ;
assign n9052 = ~ ( n7779 ) ;
assign n9053 =  ( n7784 ) | ( n6524 )  ;
assign n9054 = ~ ( n9053 ) ;
assign n9055 =  ( n9052 ) | ( n9054 )  ;
assign n9056 = ~ ( n7801 ) ;
assign n9057 =  ( n9055 ) | ( n9056 )  ;
assign n9058 =  ( n9018 ) ^ ( n9057 )  ;
assign n9059 = ~ ( n7809 ) ;
assign n9060 = ~ ( n6553 ) ;
assign n9061 =  ( n9059 ) | ( n9060 )  ;
assign n9062 =  ( n9058 ) ^ ( n9061 )  ;
assign n9063 = ~ ( n8761 ) ;
assign n9064 =  ( n9063 ) | ( n8771 )  ;
assign n9065 =  ( n9062 ) ^ ( n9064 )  ;
assign n9066 =  ( n9065 ) ^ ( n7455 )  ;
assign n9067 =  ( n6825 ) | ( n6834 )  ;
assign n9068 =  ( n9067 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9069 =  ( n9066 ) ^ ( n9068 )  ;
assign n9070 =  ( n6483 ) | ( n6492 )  ;
assign n9071 =  ( n9070 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9072 =  ( n9069 ) ^ ( n9071 )  ;
assign n9073 =  ( n6030 ) | ( n6039 )  ;
assign n9074 =  ( n9073 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9075 =  ( n9072 ) ^ ( n9074 )  ;
assign n9076 =  ( n5802 ) | ( n5811 )  ;
assign n9077 =  ( n9076 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9078 =  ( n9075 ) ^ ( n9077 )  ;
assign n9079 =  ( n5832 ) | ( n5841 )  ;
assign n9080 =  ( n9079 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9081 =  ( n9078 ) ^ ( n9080 )  ;
assign n9082 = ~ ( n9081 ) ;
assign n9083 =  ( n5682 ) | ( n5691 )  ;
assign n9084 =  ( n9083 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9085 = ~ ( n9084 ) ;
assign n9086 =  ( n9082 ) | ( n9085 )  ;
assign n9087 = ~ ( n9086 ) ;
assign n9088 =  ( n9051 ) | ( n9087 )  ;
assign n9089 = ~ ( n9088 ) ;
assign n9090 =  ( n9013 ) | ( n9089 )  ;
assign n9091 = ~ ( n7905 ) ;
assign n9092 = ~ ( n8835 ) ;
assign n9093 =  ( n9091 ) | ( n9092 )  ;
assign n9094 =  ( n8829 ) ^ ( n9093 )  ;
assign n9095 = ~ ( n7779 ) ;
assign n9096 =  ( n7784 ) | ( n6524 )  ;
assign n9097 = ~ ( n9096 ) ;
assign n9098 =  ( n9095 ) | ( n9097 )  ;
assign n9099 = ~ ( n7801 ) ;
assign n9100 =  ( n9098 ) | ( n9099 )  ;
assign n9101 =  ( n9094 ) ^ ( n9100 )  ;
assign n9102 = ~ ( n7809 ) ;
assign n9103 = ~ ( n6553 ) ;
assign n9104 =  ( n9102 ) | ( n9103 )  ;
assign n9105 =  ( n9101 ) ^ ( n9104 )  ;
assign n9106 =  ( n9105 ) ^ ( n7455 )  ;
assign n9107 =  ( n6825 ) | ( n6834 )  ;
assign n9108 =  ( n9107 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9109 =  ( n9106 ) ^ ( n9108 )  ;
assign n9110 =  ( n6483 ) | ( n6492 )  ;
assign n9111 =  ( n9110 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9112 =  ( n9109 ) ^ ( n9111 )  ;
assign n9113 =  ( n6030 ) | ( n6039 )  ;
assign n9114 =  ( n9113 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9115 =  ( n9112 ) ^ ( n9114 )  ;
assign n9116 =  ( n5802 ) | ( n5811 )  ;
assign n9117 =  ( n9116 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9118 =  ( n9115 ) ^ ( n9117 )  ;
assign n9119 =  ( n5832 ) | ( n5841 )  ;
assign n9120 =  ( n9119 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9121 =  ( n9118 ) ^ ( n9120 )  ;
assign n9122 =  ( n5682 ) | ( n5691 )  ;
assign n9123 =  ( n9122 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9124 =  ( n9121 ) ^ ( n9123 )  ;
assign n9125 =  ( n9124 ) ^ ( n8160 )  ;
assign n9126 =  ( n9125 ) ^ ( n8157 )  ;
assign n9127 = ~ ( n9126 ) ;
assign n9128 =  ( n9090 ) | ( n9127 )  ;
assign n9129 =  ( n8880 ) ^ ( n8490 )  ;
assign n9130 = ~ ( n7905 ) ;
assign n9131 =  ( n8179 ) | ( n8427 )  ;
assign n9132 = ~ ( n9131 ) ;
assign n9133 =  ( n9130 ) | ( n9132 )  ;
assign n9134 =  ( n9129 ) ^ ( n9133 )  ;
assign n9135 = ~ ( n7779 ) ;
assign n9136 =  ( n7784 ) | ( n6524 )  ;
assign n9137 = ~ ( n9136 ) ;
assign n9138 =  ( n9135 ) | ( n9137 )  ;
assign n9139 = ~ ( n7801 ) ;
assign n9140 =  ( n9138 ) | ( n9139 )  ;
assign n9141 =  ( n9134 ) ^ ( n9140 )  ;
assign n9142 = ~ ( n7809 ) ;
assign n9143 = ~ ( n6553 ) ;
assign n9144 =  ( n9142 ) | ( n9143 )  ;
assign n9145 =  ( n9141 ) ^ ( n9144 )  ;
assign n9146 =  ( n9145 ) ^ ( n8164 )  ;
assign n9147 =  ( n9146 ) ^ ( n7455 )  ;
assign n9148 =  ( n6825 ) | ( n6834 )  ;
assign n9149 =  ( n9148 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9150 =  ( n9147 ) ^ ( n9149 )  ;
assign n9151 =  ( n6483 ) | ( n6492 )  ;
assign n9152 =  ( n9151 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9153 =  ( n9150 ) ^ ( n9152 )  ;
assign n9154 =  ( n6030 ) | ( n6039 )  ;
assign n9155 =  ( n9154 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9156 =  ( n9153 ) ^ ( n9155 )  ;
assign n9157 =  ( n5802 ) | ( n5811 )  ;
assign n9158 =  ( n9157 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9159 =  ( n9156 ) ^ ( n9158 )  ;
assign n9160 =  ( n5832 ) | ( n5841 )  ;
assign n9161 =  ( n9160 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9162 =  ( n9159 ) ^ ( n9161 )  ;
assign n9163 =  ( n5682 ) | ( n5691 )  ;
assign n9164 =  ( n9163 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9165 =  ( n9162 ) ^ ( n9164 )  ;
assign n9166 =  ( n5713 ) | ( n5722 )  ;
assign n9167 =  ( n9166 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n9168 =  ( n9165 ) ^ ( n9167 )  ;
assign n9169 = ~ ( n9168 ) ;
assign n9170 =  ( n9128 ) | ( n9169 )  ;
assign n9171 = ~ ( n9170 ) ;
assign n9172 =  ( n8966 ) | ( n9171 )  ;
assign n9173 = ~ ( n9172 ) ;
assign n9174 =  ( n8719 ) | ( n9173 )  ;
assign n9175 = ~ ( n9174 ) ;
assign n9176 =  ( n8673 ) | ( n9175 )  ;
assign n9177 = ~ ( n9176 ) ;
assign n9178 =  ( n8122 ) | ( n9177 )  ;
assign n9179 = ~ ( n9178 ) ;
assign n9180 =  ( n8086 ) | ( n9179 )  ;
assign n9181 = ~ ( n9180 ) ;
assign n9182 =  ( n6816 ) | ( n9181 )  ;
assign n9183 = ~ ( n9182 ) ;
assign n9184 =  ( n6785 ) | ( n9183 )  ;
assign n9185 = ~ ( n5783 ) ;
assign n9186 =  ( n9185 ) | ( n5792 )  ;
assign n9187 = ~ ( n6006 ) ;
assign n9188 =  ( n9186 ) | ( n9187 )  ;
assign n9189 =  ( n9188 ) | ( n6020 )  ;
assign n9190 = ~ ( n6297 ) ;
assign n9191 =  ( n9189 ) | ( n9190 )  ;
assign n9192 =  ( n9191 ) | ( n6314 )  ;
assign n9193 = ~ ( n6473 ) ;
assign n9194 =  ( n9192 ) | ( n9193 )  ;
assign n9195 =  ( n9194 ) | ( n6815 )  ;
assign n9196 = ~ ( n7117 ) ;
assign n9197 =  ( n9195 ) | ( n9196 )  ;
assign n9198 =  ( n9197 ) | ( n7445 )  ;
assign n9199 = ~ ( n7765 ) ;
assign n9200 =  ( n9198 ) | ( n9199 )  ;
assign n9201 =  ( n9200 ) | ( n8121 )  ;
assign n9202 = ~ ( n8413 ) ;
assign n9203 =  ( n9201 ) | ( n9202 )  ;
assign n9204 = ~ ( n8717 ) ;
assign n9205 =  ( n9203 ) | ( n9204 )  ;
assign n9206 = ~ ( n9012 ) ;
assign n9207 =  ( n9205 ) | ( n9206 )  ;
assign n9208 = ~ ( n9088 ) ;
assign n9209 = ~ ( n9126 ) ;
assign n9210 =  ( n9208 ) | ( n9209 )  ;
assign n9211 = ~ ( n9210 ) ;
assign n9212 =  ( n9211 ) ^ ( n8880 )  ;
assign n9213 =  ( n9212 ) ^ ( n8490 )  ;
assign n9214 = ~ ( n7905 ) ;
assign n9215 =  ( n8179 ) | ( n8427 )  ;
assign n9216 = ~ ( n9215 ) ;
assign n9217 =  ( n9214 ) | ( n9216 )  ;
assign n9218 =  ( n9213 ) ^ ( n9217 )  ;
assign n9219 = ~ ( n7779 ) ;
assign n9220 =  ( n7784 ) | ( n6524 )  ;
assign n9221 = ~ ( n9220 ) ;
assign n9222 =  ( n9219 ) | ( n9221 )  ;
assign n9223 = ~ ( n7801 ) ;
assign n9224 =  ( n9222 ) | ( n9223 )  ;
assign n9225 =  ( n9218 ) ^ ( n9224 )  ;
assign n9226 = ~ ( n7809 ) ;
assign n9227 = ~ ( n6553 ) ;
assign n9228 =  ( n9226 ) | ( n9227 )  ;
assign n9229 =  ( n9225 ) ^ ( n9228 )  ;
assign n9230 =  ( n9229 ) ^ ( n8164 )  ;
assign n9231 =  ( n9230 ) ^ ( n7455 )  ;
assign n9232 =  ( n6825 ) | ( n6834 )  ;
assign n9233 =  ( n9232 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9234 =  ( n9231 ) ^ ( n9233 )  ;
assign n9235 =  ( n6483 ) | ( n6492 )  ;
assign n9236 =  ( n9235 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9237 =  ( n9234 ) ^ ( n9236 )  ;
assign n9238 =  ( n6030 ) | ( n6039 )  ;
assign n9239 =  ( n9238 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9240 =  ( n9237 ) ^ ( n9239 )  ;
assign n9241 =  ( n5802 ) | ( n5811 )  ;
assign n9242 =  ( n9241 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9243 =  ( n9240 ) ^ ( n9242 )  ;
assign n9244 =  ( n5832 ) | ( n5841 )  ;
assign n9245 =  ( n9244 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9246 =  ( n9243 ) ^ ( n9245 )  ;
assign n9247 =  ( n5682 ) | ( n5691 )  ;
assign n9248 =  ( n9247 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9249 =  ( n9246 ) ^ ( n9248 )  ;
assign n9250 =  ( n5713 ) | ( n5722 )  ;
assign n9251 =  ( n9250 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n9252 =  ( n9249 ) ^ ( n9251 )  ;
assign n9253 = ~ ( n9252 ) ;
assign n9254 =  ( n9207 ) | ( n9253 )  ;
assign n9255 = ~ ( n9018 ) ;
assign n9256 = ~ ( n7779 ) ;
assign n9257 =  ( n7784 ) | ( n6524 )  ;
assign n9258 = ~ ( n9257 ) ;
assign n9259 =  ( n9256 ) | ( n9258 )  ;
assign n9260 = ~ ( n7801 ) ;
assign n9261 =  ( n9259 ) | ( n9260 )  ;
assign n9262 = ~ ( n7809 ) ;
assign n9263 = ~ ( n6553 ) ;
assign n9264 =  ( n9262 ) | ( n9263 )  ;
assign n9265 =  ( n9261 ) ^ ( n9264 )  ;
assign n9266 =  ( n9265 ) ^ ( n7455 )  ;
assign n9267 =  ( n6825 ) | ( n6834 )  ;
assign n9268 =  ( n9267 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9269 =  ( n9266 ) ^ ( n9268 )  ;
assign n9270 =  ( n6483 ) | ( n6492 )  ;
assign n9271 =  ( n9270 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9272 =  ( n9269 ) ^ ( n9271 )  ;
assign n9273 =  ( n6030 ) | ( n6039 )  ;
assign n9274 =  ( n9273 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9275 =  ( n9272 ) ^ ( n9274 )  ;
assign n9276 =  ( n5802 ) | ( n5811 )  ;
assign n9277 =  ( n9276 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9278 =  ( n9275 ) ^ ( n9277 )  ;
assign n9279 = ~ ( n9278 ) ;
assign n9280 =  ( n9255 ) | ( n9279 )  ;
assign n9281 = ~ ( n9280 ) ;
assign n9282 = ~ ( n7779 ) ;
assign n9283 =  ( n7784 ) | ( n6524 )  ;
assign n9284 = ~ ( n9283 ) ;
assign n9285 =  ( n9282 ) | ( n9284 )  ;
assign n9286 = ~ ( n7801 ) ;
assign n9287 =  ( n9285 ) | ( n9286 )  ;
assign n9288 =  ( n9018 ) ^ ( n9287 )  ;
assign n9289 = ~ ( n7809 ) ;
assign n9290 = ~ ( n6553 ) ;
assign n9291 =  ( n9289 ) | ( n9290 )  ;
assign n9292 =  ( n9288 ) ^ ( n9291 )  ;
assign n9293 =  ( n9292 ) ^ ( n7455 )  ;
assign n9294 =  ( n6825 ) | ( n6834 )  ;
assign n9295 =  ( n9294 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9296 =  ( n9293 ) ^ ( n9295 )  ;
assign n9297 =  ( n6483 ) | ( n6492 )  ;
assign n9298 =  ( n9297 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9299 =  ( n9296 ) ^ ( n9298 )  ;
assign n9300 =  ( n6030 ) | ( n6039 )  ;
assign n9301 =  ( n9300 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9302 =  ( n9299 ) ^ ( n9301 )  ;
assign n9303 =  ( n5802 ) | ( n5811 )  ;
assign n9304 =  ( n9303 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9305 =  ( n9302 ) ^ ( n9304 )  ;
assign n9306 = ~ ( n9305 ) ;
assign n9307 =  ( n5832 ) | ( n5841 )  ;
assign n9308 =  ( n9307 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9309 =  ( n9308 ) ^ ( n8759 )  ;
assign n9310 =  ( n9309 ) ^ ( n8756 )  ;
assign n9311 = ~ ( n9310 ) ;
assign n9312 =  ( n9306 ) | ( n9311 )  ;
assign n9313 = ~ ( n9312 ) ;
assign n9314 =  ( n9281 ) | ( n9313 )  ;
assign n9315 = ~ ( n9314 ) ;
assign n9316 = ~ ( n7779 ) ;
assign n9317 =  ( n7784 ) | ( n6524 )  ;
assign n9318 = ~ ( n9317 ) ;
assign n9319 =  ( n9316 ) | ( n9318 )  ;
assign n9320 = ~ ( n7801 ) ;
assign n9321 =  ( n9319 ) | ( n9320 )  ;
assign n9322 =  ( n9018 ) ^ ( n9321 )  ;
assign n9323 = ~ ( n7809 ) ;
assign n9324 = ~ ( n6553 ) ;
assign n9325 =  ( n9323 ) | ( n9324 )  ;
assign n9326 =  ( n9322 ) ^ ( n9325 )  ;
assign n9327 = ~ ( n8761 ) ;
assign n9328 =  ( n9327 ) | ( n8771 )  ;
assign n9329 =  ( n9326 ) ^ ( n9328 )  ;
assign n9330 =  ( n9329 ) ^ ( n7455 )  ;
assign n9331 =  ( n6825 ) | ( n6834 )  ;
assign n9332 =  ( n9331 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9333 =  ( n9330 ) ^ ( n9332 )  ;
assign n9334 =  ( n6483 ) | ( n6492 )  ;
assign n9335 =  ( n9334 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9336 =  ( n9333 ) ^ ( n9335 )  ;
assign n9337 =  ( n6030 ) | ( n6039 )  ;
assign n9338 =  ( n9337 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9339 =  ( n9336 ) ^ ( n9338 )  ;
assign n9340 =  ( n5802 ) | ( n5811 )  ;
assign n9341 =  ( n9340 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9342 =  ( n9339 ) ^ ( n9341 )  ;
assign n9343 =  ( n5832 ) | ( n5841 )  ;
assign n9344 =  ( n9343 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9345 =  ( n9342 ) ^ ( n9344 )  ;
assign n9346 =  ( n5682 ) | ( n5691 )  ;
assign n9347 =  ( n9346 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9348 =  ( n9345 ) ^ ( n9347 )  ;
assign n9349 = ~ ( n9348 ) ;
assign n9350 =  ( n9315 ) | ( n9349 )  ;
assign n9351 =  ( n9088 ) ^ ( n8829 )  ;
assign n9352 = ~ ( n7905 ) ;
assign n9353 = ~ ( n8835 ) ;
assign n9354 =  ( n9352 ) | ( n9353 )  ;
assign n9355 =  ( n9351 ) ^ ( n9354 )  ;
assign n9356 = ~ ( n7779 ) ;
assign n9357 =  ( n7784 ) | ( n6524 )  ;
assign n9358 = ~ ( n9357 ) ;
assign n9359 =  ( n9356 ) | ( n9358 )  ;
assign n9360 = ~ ( n7801 ) ;
assign n9361 =  ( n9359 ) | ( n9360 )  ;
assign n9362 =  ( n9355 ) ^ ( n9361 )  ;
assign n9363 = ~ ( n7809 ) ;
assign n9364 = ~ ( n6553 ) ;
assign n9365 =  ( n9363 ) | ( n9364 )  ;
assign n9366 =  ( n9362 ) ^ ( n9365 )  ;
assign n9367 =  ( n9366 ) ^ ( n7455 )  ;
assign n9368 =  ( n6825 ) | ( n6834 )  ;
assign n9369 =  ( n9368 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9370 =  ( n9367 ) ^ ( n9369 )  ;
assign n9371 =  ( n6483 ) | ( n6492 )  ;
assign n9372 =  ( n9371 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9373 =  ( n9370 ) ^ ( n9372 )  ;
assign n9374 =  ( n6030 ) | ( n6039 )  ;
assign n9375 =  ( n9374 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9376 =  ( n9373 ) ^ ( n9375 )  ;
assign n9377 =  ( n5802 ) | ( n5811 )  ;
assign n9378 =  ( n9377 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9379 =  ( n9376 ) ^ ( n9378 )  ;
assign n9380 =  ( n5832 ) | ( n5841 )  ;
assign n9381 =  ( n9380 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9382 =  ( n9379 ) ^ ( n9381 )  ;
assign n9383 =  ( n5682 ) | ( n5691 )  ;
assign n9384 =  ( n9383 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9385 =  ( n9382 ) ^ ( n9384 )  ;
assign n9386 =  ( n9385 ) ^ ( n8160 )  ;
assign n9387 =  ( n9386 ) ^ ( n8157 )  ;
assign n9388 = ~ ( n9387 ) ;
assign n9389 =  ( n9350 ) | ( n9388 )  ;
assign n9390 = ~ ( n9389 ) ;
assign n9391 = ~ ( n9314 ) ;
assign n9392 = ~ ( n9348 ) ;
assign n9393 =  ( n9391 ) | ( n9392 )  ;
assign n9394 = ~ ( n9393 ) ;
assign n9395 =  ( n9394 ) ^ ( n9088 )  ;
assign n9396 =  ( n9395 ) ^ ( n8829 )  ;
assign n9397 = ~ ( n7905 ) ;
assign n9398 = ~ ( n8835 ) ;
assign n9399 =  ( n9397 ) | ( n9398 )  ;
assign n9400 =  ( n9396 ) ^ ( n9399 )  ;
assign n9401 = ~ ( n7779 ) ;
assign n9402 =  ( n7784 ) | ( n6524 )  ;
assign n9403 = ~ ( n9402 ) ;
assign n9404 =  ( n9401 ) | ( n9403 )  ;
assign n9405 = ~ ( n7801 ) ;
assign n9406 =  ( n9404 ) | ( n9405 )  ;
assign n9407 =  ( n9400 ) ^ ( n9406 )  ;
assign n9408 = ~ ( n7809 ) ;
assign n9409 = ~ ( n6553 ) ;
assign n9410 =  ( n9408 ) | ( n9409 )  ;
assign n9411 =  ( n9407 ) ^ ( n9410 )  ;
assign n9412 =  ( n9411 ) ^ ( n7455 )  ;
assign n9413 =  ( n6825 ) | ( n6834 )  ;
assign n9414 =  ( n9413 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9415 =  ( n9412 ) ^ ( n9414 )  ;
assign n9416 =  ( n6483 ) | ( n6492 )  ;
assign n9417 =  ( n9416 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9418 =  ( n9415 ) ^ ( n9417 )  ;
assign n9419 =  ( n6030 ) | ( n6039 )  ;
assign n9420 =  ( n9419 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9421 =  ( n9418 ) ^ ( n9420 )  ;
assign n9422 =  ( n5802 ) | ( n5811 )  ;
assign n9423 =  ( n9422 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9424 =  ( n9421 ) ^ ( n9423 )  ;
assign n9425 =  ( n5832 ) | ( n5841 )  ;
assign n9426 =  ( n9425 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9427 =  ( n9424 ) ^ ( n9426 )  ;
assign n9428 =  ( n5682 ) | ( n5691 )  ;
assign n9429 =  ( n9428 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9430 =  ( n9427 ) ^ ( n9429 )  ;
assign n9431 =  ( n9430 ) ^ ( n8160 )  ;
assign n9432 =  ( n9431 ) ^ ( n8157 )  ;
assign n9433 = ~ ( n9432 ) ;
assign n9434 = ~ ( n7809 ) ;
assign n9435 = ~ ( n6553 ) ;
assign n9436 =  ( n9434 ) | ( n9435 )  ;
assign n9437 = ~ ( n9436 ) ;
assign n9438 =  ( n7804 ) | ( n9437 )  ;
assign n9439 =  ( n9438 ) | ( n8179 )  ;
assign n9440 = kd[11:11] ;
assign n9441 =  ( n9440 ) == ( bv_1_0_n2 )  ;
assign n9442 = kd[10:10] ;
assign n9443 =  ( n9442 ) == ( bv_1_1_n5 )  ;
assign n9444 =  ( n9441 ) | ( n9443 )  ;
assign n9445 = kd[9:9] ;
assign n9446 =  ( n9445 ) == ( bv_1_1_n5 )  ;
assign n9447 =  ( n9444 ) | ( n9446 )  ;
assign n9448 = ~ ( n9447 )  ;
assign n9449 = kd[11:11] ;
assign n9450 =  ( n9449 ) == ( bv_1_1_n5 )  ;
assign n9451 = kd[10:10] ;
assign n9452 =  ( n9451 ) == ( bv_1_0_n2 )  ;
assign n9453 =  ( n9450 ) | ( n9452 )  ;
assign n9454 = kd[9:9] ;
assign n9455 =  ( n9454 ) == ( bv_1_0_n2 )  ;
assign n9456 =  ( n9453 ) | ( n9455 )  ;
assign n9457 = ~ ( n9456 )  ;
assign n9458 =  ( n9448 ) | ( n9457 )  ;
assign n9459 = kd[11:11] ;
assign n9460 = ~ ( n9459 ) ;
assign n9461 = kd[10:10] ;
assign n9462 = ~ ( n9461 ) ;
assign n9463 = kd[9:9] ;
assign n9464 = ~ ( n9463 ) ;
assign n9465 =  ( n9462 ) | ( n9464 )  ;
assign n9466 = ~ ( n9465 ) ;
assign n9467 =  ( n9460 ) | ( n9466 )  ;
assign n9468 = ~ ( n9467 ) ;
assign n9469 =  ( n5832 ) | ( n5841 )  ;
assign n9470 =  ( n9469 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9471 =  ( n9458 ) ? ( n9468 ) : ( n9470 ) ;
assign n9472 = ~ ( n9471 ) ;
assign n9473 =  ( n9439 ) | ( n9472 )  ;
assign n9474 = ~ ( n9473 ) ;
assign n9475 = ~ ( n7845 ) ;
assign n9476 =  ( n6825 ) | ( n6834 )  ;
assign n9477 =  ( n9476 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9478 =  ( n7455 ) ^ ( n9477 )  ;
assign n9479 =  ( n6483 ) | ( n6492 )  ;
assign n9480 =  ( n9479 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9481 =  ( n9478 ) ^ ( n9480 )  ;
assign n9482 =  ( n6030 ) | ( n6039 )  ;
assign n9483 =  ( n9482 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9484 =  ( n9481 ) ^ ( n9483 )  ;
assign n9485 =  ( n5802 ) | ( n5811 )  ;
assign n9486 =  ( n9485 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9487 =  ( n9484 ) ^ ( n9486 )  ;
assign n9488 =  ( n9487 ) ^ ( n9471 )  ;
assign n9489 = ~ ( n9488 ) ;
assign n9490 =  ( n9475 ) | ( n9489 )  ;
assign n9491 = ~ ( n9490 ) ;
assign n9492 =  ( n9474 ) | ( n9491 )  ;
assign n9493 = ~ ( n7779 ) ;
assign n9494 =  ( n7784 ) | ( n6524 )  ;
assign n9495 = ~ ( n9494 ) ;
assign n9496 =  ( n9493 ) | ( n9495 )  ;
assign n9497 = ~ ( n7801 ) ;
assign n9498 =  ( n9496 ) | ( n9497 )  ;
assign n9499 = ~ ( n7809 ) ;
assign n9500 = ~ ( n6553 ) ;
assign n9501 =  ( n9499 ) | ( n9500 )  ;
assign n9502 =  ( n9498 ) ^ ( n9501 )  ;
assign n9503 =  ( n9502 ) ^ ( n7455 )  ;
assign n9504 =  ( n6825 ) | ( n6834 )  ;
assign n9505 =  ( n9504 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9506 =  ( n9503 ) ^ ( n9505 )  ;
assign n9507 =  ( n6483 ) | ( n6492 )  ;
assign n9508 =  ( n9507 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9509 =  ( n9506 ) ^ ( n9508 )  ;
assign n9510 =  ( n6030 ) | ( n6039 )  ;
assign n9511 =  ( n9510 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9512 =  ( n9509 ) ^ ( n9511 )  ;
assign n9513 =  ( n5802 ) | ( n5811 )  ;
assign n9514 =  ( n9513 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9515 =  ( n9512 ) ^ ( n9514 )  ;
assign n9516 =  ( n9515 ) ^ ( n9471 )  ;
assign n9517 = ~ ( n9516 ) ;
assign n9518 = kd[11:11] ;
assign n9519 = ~ ( n9518 ) ;
assign n9520 =  ( n9517 ) | ( n9519 )  ;
assign n9521 =  ( n9520 ) | ( n9466 )  ;
assign n9522 = ~ ( n9521 ) ;
assign n9523 =  ( n9492 ) | ( n9522 )  ;
assign n9524 = ~ ( n9523 ) ;
assign n9525 = ~ ( n7905 ) ;
assign n9526 = ~ ( n9471 ) ;
assign n9527 =  ( n8179 ) | ( n9526 )  ;
assign n9528 = ~ ( n9527 ) ;
assign n9529 =  ( n9525 ) | ( n9528 )  ;
assign n9530 = ~ ( n9529 ) ;
assign n9531 =  ( n9524 ) | ( n9530 )  ;
assign n9532 = ~ ( n9531 ) ;
assign n9533 =  ( n9523 ) ^ ( n9529 )  ;
assign n9534 = ~ ( n9533 ) ;
assign n9535 = ~ ( n9278 ) ;
assign n9536 =  ( n9534 ) | ( n9535 )  ;
assign n9537 = ~ ( n9536 ) ;
assign n9538 =  ( n9532 ) | ( n9537 )  ;
assign n9539 = ~ ( n9538 ) ;
assign n9540 =  ( n9433 ) | ( n9539 )  ;
assign n9541 = ~ ( n7779 ) ;
assign n9542 =  ( n7784 ) | ( n6524 )  ;
assign n9543 = ~ ( n9542 ) ;
assign n9544 =  ( n9541 ) | ( n9543 )  ;
assign n9545 = ~ ( n7801 ) ;
assign n9546 =  ( n9544 ) | ( n9545 )  ;
assign n9547 =  ( n9018 ) ^ ( n9546 )  ;
assign n9548 = ~ ( n7809 ) ;
assign n9549 = ~ ( n6553 ) ;
assign n9550 =  ( n9548 ) | ( n9549 )  ;
assign n9551 =  ( n9547 ) ^ ( n9550 )  ;
assign n9552 =  ( n9551 ) ^ ( n7455 )  ;
assign n9553 =  ( n6825 ) | ( n6834 )  ;
assign n9554 =  ( n9553 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9555 =  ( n9552 ) ^ ( n9554 )  ;
assign n9556 =  ( n6483 ) | ( n6492 )  ;
assign n9557 =  ( n9556 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9558 =  ( n9555 ) ^ ( n9557 )  ;
assign n9559 =  ( n6030 ) | ( n6039 )  ;
assign n9560 =  ( n9559 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9561 =  ( n9558 ) ^ ( n9560 )  ;
assign n9562 =  ( n5802 ) | ( n5811 )  ;
assign n9563 =  ( n9562 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9564 =  ( n9561 ) ^ ( n9563 )  ;
assign n9565 =  ( n5832 ) | ( n5841 )  ;
assign n9566 =  ( n9565 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9567 =  ( n9564 ) ^ ( n9566 )  ;
assign n9568 =  ( n9567 ) ^ ( n8759 )  ;
assign n9569 =  ( n9568 ) ^ ( n8756 )  ;
assign n9570 = ~ ( n9569 ) ;
assign n9571 =  ( n9540 ) | ( n9570 )  ;
assign n9572 =  ( n9314 ) ^ ( n9018 )  ;
assign n9573 = ~ ( n7779 ) ;
assign n9574 =  ( n7784 ) | ( n6524 )  ;
assign n9575 = ~ ( n9574 ) ;
assign n9576 =  ( n9573 ) | ( n9575 )  ;
assign n9577 = ~ ( n7801 ) ;
assign n9578 =  ( n9576 ) | ( n9577 )  ;
assign n9579 =  ( n9572 ) ^ ( n9578 )  ;
assign n9580 = ~ ( n7809 ) ;
assign n9581 = ~ ( n6553 ) ;
assign n9582 =  ( n9580 ) | ( n9581 )  ;
assign n9583 =  ( n9579 ) ^ ( n9582 )  ;
assign n9584 = ~ ( n8761 ) ;
assign n9585 =  ( n9584 ) | ( n8771 )  ;
assign n9586 =  ( n9583 ) ^ ( n9585 )  ;
assign n9587 =  ( n9586 ) ^ ( n7455 )  ;
assign n9588 =  ( n6825 ) | ( n6834 )  ;
assign n9589 =  ( n9588 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9590 =  ( n9587 ) ^ ( n9589 )  ;
assign n9591 =  ( n6483 ) | ( n6492 )  ;
assign n9592 =  ( n9591 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9593 =  ( n9590 ) ^ ( n9592 )  ;
assign n9594 =  ( n6030 ) | ( n6039 )  ;
assign n9595 =  ( n9594 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9596 =  ( n9593 ) ^ ( n9595 )  ;
assign n9597 =  ( n5802 ) | ( n5811 )  ;
assign n9598 =  ( n9597 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9599 =  ( n9596 ) ^ ( n9598 )  ;
assign n9600 =  ( n5832 ) | ( n5841 )  ;
assign n9601 =  ( n9600 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9602 =  ( n9599 ) ^ ( n9601 )  ;
assign n9603 =  ( n5682 ) | ( n5691 )  ;
assign n9604 =  ( n9603 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9605 =  ( n9602 ) ^ ( n9604 )  ;
assign n9606 = ~ ( n9605 ) ;
assign n9607 =  ( n9571 ) | ( n9606 )  ;
assign n9608 = ~ ( n9607 ) ;
assign n9609 =  ( n9390 ) | ( n9608 )  ;
assign n9610 = ~ ( n9432 ) ;
assign n9611 = ~ ( n9538 ) ;
assign n9612 = ~ ( n9569 ) ;
assign n9613 =  ( n9611 ) | ( n9612 )  ;
assign n9614 = ~ ( n9613 ) ;
assign n9615 =  ( n9614 ) ^ ( n9314 )  ;
assign n9616 =  ( n9615 ) ^ ( n9018 )  ;
assign n9617 = ~ ( n7779 ) ;
assign n9618 =  ( n7784 ) | ( n6524 )  ;
assign n9619 = ~ ( n9618 ) ;
assign n9620 =  ( n9617 ) | ( n9619 )  ;
assign n9621 = ~ ( n7801 ) ;
assign n9622 =  ( n9620 ) | ( n9621 )  ;
assign n9623 =  ( n9616 ) ^ ( n9622 )  ;
assign n9624 = ~ ( n7809 ) ;
assign n9625 = ~ ( n6553 ) ;
assign n9626 =  ( n9624 ) | ( n9625 )  ;
assign n9627 =  ( n9623 ) ^ ( n9626 )  ;
assign n9628 = ~ ( n8761 ) ;
assign n9629 =  ( n9628 ) | ( n8771 )  ;
assign n9630 =  ( n9627 ) ^ ( n9629 )  ;
assign n9631 =  ( n9630 ) ^ ( n7455 )  ;
assign n9632 =  ( n6825 ) | ( n6834 )  ;
assign n9633 =  ( n9632 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9634 =  ( n9631 ) ^ ( n9633 )  ;
assign n9635 =  ( n6483 ) | ( n6492 )  ;
assign n9636 =  ( n9635 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9637 =  ( n9634 ) ^ ( n9636 )  ;
assign n9638 =  ( n6030 ) | ( n6039 )  ;
assign n9639 =  ( n9638 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9640 =  ( n9637 ) ^ ( n9639 )  ;
assign n9641 =  ( n5802 ) | ( n5811 )  ;
assign n9642 =  ( n9641 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9643 =  ( n9640 ) ^ ( n9642 )  ;
assign n9644 =  ( n5832 ) | ( n5841 )  ;
assign n9645 =  ( n9644 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9646 =  ( n9643 ) ^ ( n9645 )  ;
assign n9647 =  ( n5682 ) | ( n5691 )  ;
assign n9648 =  ( n9647 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n9649 =  ( n9646 ) ^ ( n9648 )  ;
assign n9650 = ~ ( n9649 ) ;
assign n9651 =  ( n9610 ) | ( n9650 )  ;
assign n9652 =  ( n9523 ) ^ ( n9529 )  ;
assign n9653 = ~ ( n7779 ) ;
assign n9654 =  ( n7784 ) | ( n6524 )  ;
assign n9655 = ~ ( n9654 ) ;
assign n9656 =  ( n9653 ) | ( n9655 )  ;
assign n9657 = ~ ( n7801 ) ;
assign n9658 =  ( n9656 ) | ( n9657 )  ;
assign n9659 =  ( n9652 ) ^ ( n9658 )  ;
assign n9660 = ~ ( n7809 ) ;
assign n9661 = ~ ( n6553 ) ;
assign n9662 =  ( n9660 ) | ( n9661 )  ;
assign n9663 =  ( n9659 ) ^ ( n9662 )  ;
assign n9664 =  ( n9663 ) ^ ( n7455 )  ;
assign n9665 =  ( n6825 ) | ( n6834 )  ;
assign n9666 =  ( n9665 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9667 =  ( n9664 ) ^ ( n9666 )  ;
assign n9668 =  ( n6483 ) | ( n6492 )  ;
assign n9669 =  ( n9668 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9670 =  ( n9667 ) ^ ( n9669 )  ;
assign n9671 =  ( n6030 ) | ( n6039 )  ;
assign n9672 =  ( n9671 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9673 =  ( n9670 ) ^ ( n9672 )  ;
assign n9674 =  ( n5802 ) | ( n5811 )  ;
assign n9675 =  ( n9674 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9676 =  ( n9673 ) ^ ( n9675 )  ;
assign n9677 = ~ ( n9676 ) ;
assign n9678 =  ( n5832 ) | ( n5841 )  ;
assign n9679 =  ( n9678 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9680 = ~ ( n9679 ) ;
assign n9681 =  ( n9677 ) | ( n9680 )  ;
assign n9682 =  ( n9538 ) ^ ( n9018 )  ;
assign n9683 = ~ ( n7779 ) ;
assign n9684 =  ( n7784 ) | ( n6524 )  ;
assign n9685 = ~ ( n9684 ) ;
assign n9686 =  ( n9683 ) | ( n9685 )  ;
assign n9687 = ~ ( n7801 ) ;
assign n9688 =  ( n9686 ) | ( n9687 )  ;
assign n9689 =  ( n9682 ) ^ ( n9688 )  ;
assign n9690 = ~ ( n7809 ) ;
assign n9691 = ~ ( n6553 ) ;
assign n9692 =  ( n9690 ) | ( n9691 )  ;
assign n9693 =  ( n9689 ) ^ ( n9692 )  ;
assign n9694 =  ( n9693 ) ^ ( n7455 )  ;
assign n9695 =  ( n6825 ) | ( n6834 )  ;
assign n9696 =  ( n9695 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9697 =  ( n9694 ) ^ ( n9696 )  ;
assign n9698 =  ( n6483 ) | ( n6492 )  ;
assign n9699 =  ( n9698 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9700 =  ( n9697 ) ^ ( n9699 )  ;
assign n9701 =  ( n6030 ) | ( n6039 )  ;
assign n9702 =  ( n9701 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9703 =  ( n9700 ) ^ ( n9702 )  ;
assign n9704 =  ( n5802 ) | ( n5811 )  ;
assign n9705 =  ( n9704 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9706 =  ( n9703 ) ^ ( n9705 )  ;
assign n9707 =  ( n5832 ) | ( n5841 )  ;
assign n9708 =  ( n9707 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9709 =  ( n9706 ) ^ ( n9708 )  ;
assign n9710 =  ( n9709 ) ^ ( n8759 )  ;
assign n9711 =  ( n9710 ) ^ ( n8756 )  ;
assign n9712 = ~ ( n9711 ) ;
assign n9713 =  ( n9681 ) | ( n9712 )  ;
assign n9714 = ~ ( n9713 ) ;
assign n9715 = ~ ( n9676 ) ;
assign n9716 =  ( n5832 ) | ( n5841 )  ;
assign n9717 =  ( n9716 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9718 = ~ ( n9717 ) ;
assign n9719 =  ( n9715 ) | ( n9718 )  ;
assign n9720 = ~ ( n9719 ) ;
assign n9721 =  ( n9720 ) ^ ( n9538 )  ;
assign n9722 =  ( n9721 ) ^ ( n9018 )  ;
assign n9723 = ~ ( n7779 ) ;
assign n9724 =  ( n7784 ) | ( n6524 )  ;
assign n9725 = ~ ( n9724 ) ;
assign n9726 =  ( n9723 ) | ( n9725 )  ;
assign n9727 = ~ ( n7801 ) ;
assign n9728 =  ( n9726 ) | ( n9727 )  ;
assign n9729 =  ( n9722 ) ^ ( n9728 )  ;
assign n9730 = ~ ( n7809 ) ;
assign n9731 = ~ ( n6553 ) ;
assign n9732 =  ( n9730 ) | ( n9731 )  ;
assign n9733 =  ( n9729 ) ^ ( n9732 )  ;
assign n9734 =  ( n9733 ) ^ ( n7455 )  ;
assign n9735 =  ( n6825 ) | ( n6834 )  ;
assign n9736 =  ( n9735 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9737 =  ( n9734 ) ^ ( n9736 )  ;
assign n9738 =  ( n6483 ) | ( n6492 )  ;
assign n9739 =  ( n9738 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9740 =  ( n9737 ) ^ ( n9739 )  ;
assign n9741 =  ( n6030 ) | ( n6039 )  ;
assign n9742 =  ( n9741 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9743 =  ( n9740 ) ^ ( n9742 )  ;
assign n9744 =  ( n5802 ) | ( n5811 )  ;
assign n9745 =  ( n9744 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9746 =  ( n9743 ) ^ ( n9745 )  ;
assign n9747 =  ( n5832 ) | ( n5841 )  ;
assign n9748 =  ( n9747 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9749 =  ( n9746 ) ^ ( n9748 )  ;
assign n9750 =  ( n9749 ) ^ ( n8759 )  ;
assign n9751 =  ( n9750 ) ^ ( n8756 )  ;
assign n9752 = ~ ( n9751 ) ;
assign n9753 = ~ ( n7779 ) ;
assign n9754 =  ( n7784 ) | ( n6524 )  ;
assign n9755 = ~ ( n9754 ) ;
assign n9756 =  ( n9753 ) | ( n9755 )  ;
assign n9757 = kd[9:9] ;
assign n9758 =  ( n9757 ) == ( bv_1_0_n2 )  ;
assign n9759 = kd[8:8] ;
assign n9760 =  ( n9759 ) == ( bv_1_1_n5 )  ;
assign n9761 =  ( n9758 ) | ( n9760 )  ;
assign n9762 = kd[7:7] ;
assign n9763 =  ( n9762 ) == ( bv_1_1_n5 )  ;
assign n9764 =  ( n9761 ) | ( n9763 )  ;
assign n9765 = ~ ( n9764 )  ;
assign n9766 = kd[9:9] ;
assign n9767 =  ( n9766 ) == ( bv_1_1_n5 )  ;
assign n9768 = kd[8:8] ;
assign n9769 =  ( n9768 ) == ( bv_1_0_n2 )  ;
assign n9770 =  ( n9767 ) | ( n9769 )  ;
assign n9771 = kd[7:7] ;
assign n9772 =  ( n9771 ) == ( bv_1_0_n2 )  ;
assign n9773 =  ( n9770 ) | ( n9772 )  ;
assign n9774 = ~ ( n9773 )  ;
assign n9775 =  ( n9765 ) | ( n9774 )  ;
assign n9776 = kd[9:9] ;
assign n9777 = ~ ( n9776 ) ;
assign n9778 = kd[8:8] ;
assign n9779 = ~ ( n9778 ) ;
assign n9780 = kd[7:7] ;
assign n9781 = ~ ( n9780 ) ;
assign n9782 =  ( n9779 ) | ( n9781 )  ;
assign n9783 = ~ ( n9782 ) ;
assign n9784 =  ( n9777 ) | ( n9783 )  ;
assign n9785 = ~ ( n9784 ) ;
assign n9786 =  ( n5802 ) | ( n5811 )  ;
assign n9787 =  ( n9786 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9788 =  ( n9775 ) ? ( n9785 ) : ( n9787 ) ;
assign n9789 = ~ ( n9788 ) ;
assign n9790 =  ( n7797 ) | ( n9789 )  ;
assign n9791 = ~ ( n9790 ) ;
assign n9792 =  ( n9756 ) | ( n9791 )  ;
assign n9793 = ~ ( n9792 ) ;
assign n9794 = ~ ( n7809 ) ;
assign n9795 = ~ ( n6553 ) ;
assign n9796 =  ( n9794 ) | ( n9795 )  ;
assign n9797 = ~ ( n9796 ) ;
assign n9798 =  ( n9793 ) | ( n9797 )  ;
assign n9799 = ~ ( n9798 ) ;
assign n9800 = ~ ( n7809 ) ;
assign n9801 = ~ ( n6553 ) ;
assign n9802 =  ( n9800 ) | ( n9801 )  ;
assign n9803 =  ( n9792 ) ^ ( n9802 )  ;
assign n9804 = ~ ( n9803 ) ;
assign n9805 =  ( n9804 ) | ( n8179 )  ;
assign n9806 = ~ ( n9805 ) ;
assign n9807 =  ( n9799 ) | ( n9806 )  ;
assign n9808 = ~ ( n9807 ) ;
assign n9809 =  ( n9752 ) | ( n9808 )  ;
assign n9810 = ~ ( n7779 ) ;
assign n9811 =  ( n7784 ) | ( n6524 )  ;
assign n9812 = ~ ( n9811 ) ;
assign n9813 =  ( n9810 ) | ( n9812 )  ;
assign n9814 = ~ ( n7801 ) ;
assign n9815 =  ( n9813 ) | ( n9814 )  ;
assign n9816 = ~ ( n7809 ) ;
assign n9817 = ~ ( n6553 ) ;
assign n9818 =  ( n9816 ) | ( n9817 )  ;
assign n9819 =  ( n9815 ) ^ ( n9818 )  ;
assign n9820 =  ( n9819 ) ^ ( n7455 )  ;
assign n9821 =  ( n6825 ) | ( n6834 )  ;
assign n9822 =  ( n9821 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9823 =  ( n9820 ) ^ ( n9822 )  ;
assign n9824 =  ( n6483 ) | ( n6492 )  ;
assign n9825 =  ( n9824 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9826 =  ( n9823 ) ^ ( n9825 )  ;
assign n9827 =  ( n6030 ) | ( n6039 )  ;
assign n9828 =  ( n9827 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9829 =  ( n9826 ) ^ ( n9828 )  ;
assign n9830 =  ( n5802 ) | ( n5811 )  ;
assign n9831 =  ( n9830 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9832 =  ( n9829 ) ^ ( n9831 )  ;
assign n9833 =  ( n9832 ) ^ ( n9471 )  ;
assign n9834 =  ( n9833 ) ^ ( n9468 )  ;
assign n9835 = ~ ( n9834 ) ;
assign n9836 =  ( n9809 ) | ( n9835 )  ;
assign n9837 =  ( n9523 ) ^ ( n9529 )  ;
assign n9838 = ~ ( n7779 ) ;
assign n9839 =  ( n7784 ) | ( n6524 )  ;
assign n9840 = ~ ( n9839 ) ;
assign n9841 =  ( n9838 ) | ( n9840 )  ;
assign n9842 = ~ ( n7801 ) ;
assign n9843 =  ( n9841 ) | ( n9842 )  ;
assign n9844 =  ( n9837 ) ^ ( n9843 )  ;
assign n9845 = ~ ( n7809 ) ;
assign n9846 = ~ ( n6553 ) ;
assign n9847 =  ( n9845 ) | ( n9846 )  ;
assign n9848 =  ( n9844 ) ^ ( n9847 )  ;
assign n9849 =  ( n9848 ) ^ ( n7455 )  ;
assign n9850 =  ( n6825 ) | ( n6834 )  ;
assign n9851 =  ( n9850 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9852 =  ( n9849 ) ^ ( n9851 )  ;
assign n9853 =  ( n6483 ) | ( n6492 )  ;
assign n9854 =  ( n9853 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9855 =  ( n9852 ) ^ ( n9854 )  ;
assign n9856 =  ( n6030 ) | ( n6039 )  ;
assign n9857 =  ( n9856 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9858 =  ( n9855 ) ^ ( n9857 )  ;
assign n9859 =  ( n5802 ) | ( n5811 )  ;
assign n9860 =  ( n9859 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9861 =  ( n9858 ) ^ ( n9860 )  ;
assign n9862 =  ( n5832 ) | ( n5841 )  ;
assign n9863 =  ( n9862 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9864 =  ( n9861 ) ^ ( n9863 )  ;
assign n9865 = ~ ( n9864 ) ;
assign n9866 =  ( n9836 ) | ( n9865 )  ;
assign n9867 = ~ ( n9866 ) ;
assign n9868 =  ( n9714 ) | ( n9867 )  ;
assign n9869 = ~ ( n9868 ) ;
assign n9870 =  ( n9651 ) | ( n9869 )  ;
assign n9871 = ~ ( n9870 ) ;
assign n9872 =  ( n9609 ) | ( n9871 )  ;
assign n9873 = ~ ( n9432 ) ;
assign n9874 = ~ ( n9649 ) ;
assign n9875 =  ( n9873 ) | ( n9874 )  ;
assign n9876 = ~ ( n9751 ) ;
assign n9877 =  ( n9875 ) | ( n9876 )  ;
assign n9878 = ~ ( n9834 ) ;
assign n9879 =  ( n9808 ) | ( n9878 )  ;
assign n9880 = ~ ( n9879 ) ;
assign n9881 =  ( n9880 ) ^ ( n9523 )  ;
assign n9882 =  ( n9881 ) ^ ( n9529 )  ;
assign n9883 = ~ ( n7779 ) ;
assign n9884 =  ( n7784 ) | ( n6524 )  ;
assign n9885 = ~ ( n9884 ) ;
assign n9886 =  ( n9883 ) | ( n9885 )  ;
assign n9887 = ~ ( n7801 ) ;
assign n9888 =  ( n9886 ) | ( n9887 )  ;
assign n9889 =  ( n9882 ) ^ ( n9888 )  ;
assign n9890 = ~ ( n7809 ) ;
assign n9891 = ~ ( n6553 ) ;
assign n9892 =  ( n9890 ) | ( n9891 )  ;
assign n9893 =  ( n9889 ) ^ ( n9892 )  ;
assign n9894 =  ( n9893 ) ^ ( n7455 )  ;
assign n9895 =  ( n6825 ) | ( n6834 )  ;
assign n9896 =  ( n9895 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9897 =  ( n9894 ) ^ ( n9896 )  ;
assign n9898 =  ( n6483 ) | ( n6492 )  ;
assign n9899 =  ( n9898 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9900 =  ( n9897 ) ^ ( n9899 )  ;
assign n9901 =  ( n6030 ) | ( n6039 )  ;
assign n9902 =  ( n9901 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9903 =  ( n9900 ) ^ ( n9902 )  ;
assign n9904 =  ( n5802 ) | ( n5811 )  ;
assign n9905 =  ( n9904 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9906 =  ( n9903 ) ^ ( n9905 )  ;
assign n9907 =  ( n5832 ) | ( n5841 )  ;
assign n9908 =  ( n9907 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n9909 =  ( n9906 ) ^ ( n9908 )  ;
assign n9910 = ~ ( n9909 ) ;
assign n9911 =  ( n9877 ) | ( n9910 )  ;
assign n9912 = ~ ( n7809 ) ;
assign n9913 =  ( n6483 ) | ( n6492 )  ;
assign n9914 =  ( n9913 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9915 = ~ ( n9914 ) ;
assign n9916 =  ( n7784 ) | ( n9915 )  ;
assign n9917 = ~ ( n9916 ) ;
assign n9918 =  ( n9912 ) | ( n9917 )  ;
assign n9919 = ~ ( n9918 ) ;
assign n9920 =  ( n6825 ) | ( n6834 )  ;
assign n9921 =  ( n9920 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9922 =  ( n7455 ) ^ ( n9921 )  ;
assign n9923 =  ( n6483 ) | ( n6492 )  ;
assign n9924 =  ( n9923 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9925 =  ( n9922 ) ^ ( n9924 )  ;
assign n9926 =  ( n6030 ) | ( n6039 )  ;
assign n9927 =  ( n9926 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9928 =  ( n9925 ) ^ ( n9927 )  ;
assign n9929 =  ( n9928 ) ^ ( n9788 )  ;
assign n9930 = ~ ( n9929 ) ;
assign n9931 =  ( n9919 ) | ( n9930 )  ;
assign n9932 = ~ ( n9931 ) ;
assign n9933 = ~ ( n7809 ) ;
assign n9934 = ~ ( n9916 ) ;
assign n9935 =  ( n9933 ) | ( n9934 )  ;
assign n9936 =  ( n9935 ) ^ ( n7455 )  ;
assign n9937 =  ( n6825 ) | ( n6834 )  ;
assign n9938 =  ( n9937 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9939 =  ( n9936 ) ^ ( n9938 )  ;
assign n9940 =  ( n6483 ) | ( n6492 )  ;
assign n9941 =  ( n9940 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9942 =  ( n9939 ) ^ ( n9941 )  ;
assign n9943 =  ( n6030 ) | ( n6039 )  ;
assign n9944 =  ( n9943 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9945 =  ( n9942 ) ^ ( n9944 )  ;
assign n9946 =  ( n9945 ) ^ ( n9788 )  ;
assign n9947 = ~ ( n9946 ) ;
assign n9948 = kd[9:9] ;
assign n9949 = ~ ( n9948 ) ;
assign n9950 =  ( n9947 ) | ( n9949 )  ;
assign n9951 =  ( n9950 ) | ( n9783 )  ;
assign n9952 = ~ ( n9951 ) ;
assign n9953 =  ( n9932 ) | ( n9952 )  ;
assign n9954 = ~ ( n9953 ) ;
assign n9955 = ~ ( n7809 ) ;
assign n9956 = ~ ( n6553 ) ;
assign n9957 =  ( n9955 ) | ( n9956 )  ;
assign n9958 =  ( n9792 ) ^ ( n9957 )  ;
assign n9959 =  ( n9958 ) ^ ( n7455 )  ;
assign n9960 =  ( n6825 ) | ( n6834 )  ;
assign n9961 =  ( n9960 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9962 =  ( n9959 ) ^ ( n9961 )  ;
assign n9963 =  ( n6483 ) | ( n6492 )  ;
assign n9964 =  ( n9963 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9965 =  ( n9962 ) ^ ( n9964 )  ;
assign n9966 =  ( n6030 ) | ( n6039 )  ;
assign n9967 =  ( n9966 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9968 =  ( n9965 ) ^ ( n9967 )  ;
assign n9969 =  ( n5802 ) | ( n5811 )  ;
assign n9970 =  ( n9969 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n9971 =  ( n9968 ) ^ ( n9970 )  ;
assign n9972 = ~ ( n9971 ) ;
assign n9973 =  ( n9954 ) | ( n9972 )  ;
assign n9974 = ~ ( n9798 ) ;
assign n9975 =  ( n9804 ) | ( n8179 )  ;
assign n9976 = ~ ( n9975 ) ;
assign n9977 =  ( n9974 ) | ( n9976 )  ;
assign n9978 = ~ ( n7779 ) ;
assign n9979 =  ( n7784 ) | ( n6524 )  ;
assign n9980 = ~ ( n9979 ) ;
assign n9981 =  ( n9978 ) | ( n9980 )  ;
assign n9982 = ~ ( n7801 ) ;
assign n9983 =  ( n9981 ) | ( n9982 )  ;
assign n9984 =  ( n9977 ) ^ ( n9983 )  ;
assign n9985 = ~ ( n7809 ) ;
assign n9986 = ~ ( n6553 ) ;
assign n9987 =  ( n9985 ) | ( n9986 )  ;
assign n9988 =  ( n9984 ) ^ ( n9987 )  ;
assign n9989 =  ( n9988 ) ^ ( n7455 )  ;
assign n9990 =  ( n6825 ) | ( n6834 )  ;
assign n9991 =  ( n9990 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n9992 =  ( n9989 ) ^ ( n9991 )  ;
assign n9993 =  ( n6483 ) | ( n6492 )  ;
assign n9994 =  ( n9993 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n9995 =  ( n9992 ) ^ ( n9994 )  ;
assign n9996 =  ( n6030 ) | ( n6039 )  ;
assign n9997 =  ( n9996 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n9998 =  ( n9995 ) ^ ( n9997 )  ;
assign n9999 =  ( n5802 ) | ( n5811 )  ;
assign n10000 =  ( n9999 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n10001 =  ( n9998 ) ^ ( n10000 )  ;
assign n10002 =  ( n10001 ) ^ ( n9471 )  ;
assign n10003 =  ( n10002 ) ^ ( n9468 )  ;
assign n10004 = ~ ( n10003 ) ;
assign n10005 =  ( n9973 ) | ( n10004 )  ;
assign n10006 = ~ ( n10005 ) ;
assign n10007 = ~ ( n9931 ) ;
assign n10008 =  ( n10007 ) | ( n9952 )  ;
assign n10009 = ~ ( n10008 ) ;
assign n10010 =  ( n10009 ) | ( n9972 )  ;
assign n10011 = ~ ( n10010 ) ;
assign n10012 = ~ ( n9798 ) ;
assign n10013 =  ( n9804 ) | ( n8179 )  ;
assign n10014 = ~ ( n10013 ) ;
assign n10015 =  ( n10012 ) | ( n10014 )  ;
assign n10016 =  ( n10011 ) ^ ( n10015 )  ;
assign n10017 = ~ ( n7779 ) ;
assign n10018 =  ( n7784 ) | ( n6524 )  ;
assign n10019 = ~ ( n10018 ) ;
assign n10020 =  ( n10017 ) | ( n10019 )  ;
assign n10021 = ~ ( n7801 ) ;
assign n10022 =  ( n10020 ) | ( n10021 )  ;
assign n10023 =  ( n10016 ) ^ ( n10022 )  ;
assign n10024 = ~ ( n7809 ) ;
assign n10025 = ~ ( n6553 ) ;
assign n10026 =  ( n10024 ) | ( n10025 )  ;
assign n10027 =  ( n10023 ) ^ ( n10026 )  ;
assign n10028 =  ( n10027 ) ^ ( n7455 )  ;
assign n10029 =  ( n6825 ) | ( n6834 )  ;
assign n10030 =  ( n10029 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10031 =  ( n10028 ) ^ ( n10030 )  ;
assign n10032 =  ( n6483 ) | ( n6492 )  ;
assign n10033 =  ( n10032 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10034 =  ( n10031 ) ^ ( n10033 )  ;
assign n10035 =  ( n6030 ) | ( n6039 )  ;
assign n10036 =  ( n10035 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10037 =  ( n10034 ) ^ ( n10036 )  ;
assign n10038 =  ( n5802 ) | ( n5811 )  ;
assign n10039 =  ( n10038 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n10040 =  ( n10037 ) ^ ( n10039 )  ;
assign n10041 =  ( n10040 ) ^ ( n9471 )  ;
assign n10042 =  ( n10041 ) ^ ( n9468 )  ;
assign n10043 = ~ ( n10042 ) ;
assign n10044 = ~ ( n7455 ) ;
assign n10045 =  ( n6825 ) | ( n6834 )  ;
assign n10046 =  ( n10045 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10047 = ~ ( n10046 ) ;
assign n10048 =  ( n10044 ) | ( n10047 )  ;
assign n10049 =  ( n6483 ) | ( n6492 )  ;
assign n10050 =  ( n10049 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10051 = ~ ( n10050 ) ;
assign n10052 =  ( n10048 ) | ( n10051 )  ;
assign n10053 = kd[7:7] ;
assign n10054 =  ( n10053 ) == ( bv_1_0_n2 )  ;
assign n10055 = kd[6:6] ;
assign n10056 =  ( n10055 ) == ( bv_1_1_n5 )  ;
assign n10057 =  ( n10054 ) | ( n10056 )  ;
assign n10058 = kd[5:5] ;
assign n10059 =  ( n10058 ) == ( bv_1_1_n5 )  ;
assign n10060 =  ( n10057 ) | ( n10059 )  ;
assign n10061 = ~ ( n10060 )  ;
assign n10062 = kd[7:7] ;
assign n10063 =  ( n10062 ) == ( bv_1_1_n5 )  ;
assign n10064 = kd[6:6] ;
assign n10065 =  ( n10064 ) == ( bv_1_0_n2 )  ;
assign n10066 =  ( n10063 ) | ( n10065 )  ;
assign n10067 = kd[5:5] ;
assign n10068 =  ( n10067 ) == ( bv_1_0_n2 )  ;
assign n10069 =  ( n10066 ) | ( n10068 )  ;
assign n10070 = ~ ( n10069 )  ;
assign n10071 =  ( n10061 ) | ( n10070 )  ;
assign n10072 = kd[7:7] ;
assign n10073 = ~ ( n10072 ) ;
assign n10074 = kd[6:6] ;
assign n10075 = ~ ( n10074 ) ;
assign n10076 = kd[5:5] ;
assign n10077 = ~ ( n10076 ) ;
assign n10078 =  ( n10075 ) | ( n10077 )  ;
assign n10079 = ~ ( n10078 ) ;
assign n10080 =  ( n10073 ) | ( n10079 )  ;
assign n10081 = ~ ( n10080 ) ;
assign n10082 =  ( n6030 ) | ( n6039 )  ;
assign n10083 =  ( n10082 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10084 =  ( n10071 ) ? ( n10081 ) : ( n10083 ) ;
assign n10085 = ~ ( n10084 ) ;
assign n10086 =  ( n10052 ) | ( n10085 )  ;
assign n10087 = ~ ( n10086 ) ;
assign n10088 =  ( n6483 ) | ( n6492 )  ;
assign n10089 =  ( n10088 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10090 =  ( n10089 ) ^ ( n10084 )  ;
assign n10091 = ~ ( n10090 ) ;
assign n10092 =  ( n7784 ) | ( n10091 )  ;
assign n10093 = ~ ( n10092 ) ;
assign n10094 =  ( n10087 ) | ( n10093 )  ;
assign n10095 =  ( n6825 ) | ( n6834 )  ;
assign n10096 =  ( n10095 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10097 =  ( n7455 ) ^ ( n10096 )  ;
assign n10098 =  ( n6483 ) | ( n6492 )  ;
assign n10099 =  ( n10098 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10100 =  ( n10097 ) ^ ( n10099 )  ;
assign n10101 =  ( n10100 ) ^ ( n10084 )  ;
assign n10102 = ~ ( n10101 ) ;
assign n10103 = kd[7:7] ;
assign n10104 = ~ ( n10103 ) ;
assign n10105 =  ( n10102 ) | ( n10104 )  ;
assign n10106 =  ( n10105 ) | ( n10079 )  ;
assign n10107 = ~ ( n10106 ) ;
assign n10108 =  ( n10094 ) | ( n10107 )  ;
assign n10109 = ~ ( n10108 ) ;
assign n10110 = ~ ( n7809 ) ;
assign n10111 =  ( n6483 ) | ( n6492 )  ;
assign n10112 =  ( n10111 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10113 = ~ ( n10112 ) ;
assign n10114 = ~ ( n10084 ) ;
assign n10115 =  ( n10113 ) | ( n10114 )  ;
assign n10116 = ~ ( n10115 ) ;
assign n10117 =  ( n10110 ) | ( n10116 )  ;
assign n10118 = ~ ( n10117 ) ;
assign n10119 =  ( n10109 ) | ( n10118 )  ;
assign n10120 = ~ ( n10119 ) ;
assign n10121 = ~ ( n10086 ) ;
assign n10122 =  ( n7784 ) | ( n10091 )  ;
assign n10123 = ~ ( n10122 ) ;
assign n10124 =  ( n10121 ) | ( n10123 )  ;
assign n10125 =  ( n10124 ) | ( n10107 )  ;
assign n10126 = ~ ( n7809 ) ;
assign n10127 = ~ ( n10115 ) ;
assign n10128 =  ( n10126 ) | ( n10127 )  ;
assign n10129 =  ( n10125 ) ^ ( n10128 )  ;
assign n10130 = ~ ( n10129 ) ;
assign n10131 =  ( n6825 ) | ( n6834 )  ;
assign n10132 =  ( n10131 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10133 =  ( n7455 ) ^ ( n10132 )  ;
assign n10134 =  ( n6483 ) | ( n6492 )  ;
assign n10135 =  ( n10134 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10136 =  ( n10133 ) ^ ( n10135 )  ;
assign n10137 = ~ ( n10136 ) ;
assign n10138 =  ( n10130 ) | ( n10137 )  ;
assign n10139 = ~ ( n10138 ) ;
assign n10140 =  ( n10120 ) | ( n10139 )  ;
assign n10141 = ~ ( n10140 ) ;
assign n10142 =  ( n10043 ) | ( n10141 )  ;
assign n10143 = ~ ( n7809 ) ;
assign n10144 = ~ ( n9916 ) ;
assign n10145 =  ( n10143 ) | ( n10144 )  ;
assign n10146 =  ( n10145 ) ^ ( n7455 )  ;
assign n10147 =  ( n6825 ) | ( n6834 )  ;
assign n10148 =  ( n10147 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10149 =  ( n10146 ) ^ ( n10148 )  ;
assign n10150 =  ( n6483 ) | ( n6492 )  ;
assign n10151 =  ( n10150 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10152 =  ( n10149 ) ^ ( n10151 )  ;
assign n10153 =  ( n6030 ) | ( n6039 )  ;
assign n10154 =  ( n10153 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10155 =  ( n10152 ) ^ ( n10154 )  ;
assign n10156 =  ( n10155 ) ^ ( n9788 )  ;
assign n10157 =  ( n10156 ) ^ ( n9785 )  ;
assign n10158 = ~ ( n10157 ) ;
assign n10159 =  ( n10142 ) | ( n10158 )  ;
assign n10160 = ~ ( n9931 ) ;
assign n10161 =  ( n10160 ) | ( n9952 )  ;
assign n10162 =  ( n10161 ) ^ ( n9792 )  ;
assign n10163 = ~ ( n7809 ) ;
assign n10164 = ~ ( n6553 ) ;
assign n10165 =  ( n10163 ) | ( n10164 )  ;
assign n10166 =  ( n10162 ) ^ ( n10165 )  ;
assign n10167 =  ( n10166 ) ^ ( n7455 )  ;
assign n10168 =  ( n6825 ) | ( n6834 )  ;
assign n10169 =  ( n10168 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10170 =  ( n10167 ) ^ ( n10169 )  ;
assign n10171 =  ( n6483 ) | ( n6492 )  ;
assign n10172 =  ( n10171 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10173 =  ( n10170 ) ^ ( n10172 )  ;
assign n10174 =  ( n6030 ) | ( n6039 )  ;
assign n10175 =  ( n10174 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10176 =  ( n10173 ) ^ ( n10175 )  ;
assign n10177 =  ( n5802 ) | ( n5811 )  ;
assign n10178 =  ( n10177 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n10179 =  ( n10176 ) ^ ( n10178 )  ;
assign n10180 = ~ ( n10179 ) ;
assign n10181 =  ( n10159 ) | ( n10180 )  ;
assign n10182 = ~ ( n10181 ) ;
assign n10183 =  ( n10006 ) | ( n10182 )  ;
assign n10184 = ~ ( n10042 ) ;
assign n10185 = ~ ( n10140 ) ;
assign n10186 =  ( n10185 ) | ( n10158 )  ;
assign n10187 = ~ ( n10186 ) ;
assign n10188 = ~ ( n9931 ) ;
assign n10189 =  ( n10188 ) | ( n9952 )  ;
assign n10190 =  ( n10187 ) ^ ( n10189 )  ;
assign n10191 =  ( n10190 ) ^ ( n9792 )  ;
assign n10192 = ~ ( n7809 ) ;
assign n10193 = ~ ( n6553 ) ;
assign n10194 =  ( n10192 ) | ( n10193 )  ;
assign n10195 =  ( n10191 ) ^ ( n10194 )  ;
assign n10196 =  ( n10195 ) ^ ( n7455 )  ;
assign n10197 =  ( n6825 ) | ( n6834 )  ;
assign n10198 =  ( n10197 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10199 =  ( n10196 ) ^ ( n10198 )  ;
assign n10200 =  ( n6483 ) | ( n6492 )  ;
assign n10201 =  ( n10200 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10202 =  ( n10199 ) ^ ( n10201 )  ;
assign n10203 =  ( n6030 ) | ( n6039 )  ;
assign n10204 =  ( n10203 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10205 =  ( n10202 ) ^ ( n10204 )  ;
assign n10206 =  ( n5802 ) | ( n5811 )  ;
assign n10207 =  ( n10206 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n10208 =  ( n10205 ) ^ ( n10207 )  ;
assign n10209 = ~ ( n10208 ) ;
assign n10210 =  ( n10184 ) | ( n10209 )  ;
assign n10211 = ~ ( n10086 ) ;
assign n10212 =  ( n7784 ) | ( n10091 )  ;
assign n10213 = ~ ( n10212 ) ;
assign n10214 =  ( n10211 ) | ( n10213 )  ;
assign n10215 =  ( n10214 ) | ( n10107 )  ;
assign n10216 = ~ ( n7809 ) ;
assign n10217 = ~ ( n10115 ) ;
assign n10218 =  ( n10216 ) | ( n10217 )  ;
assign n10219 =  ( n10215 ) ^ ( n10218 )  ;
assign n10220 =  ( n10219 ) ^ ( n7455 )  ;
assign n10221 =  ( n6825 ) | ( n6834 )  ;
assign n10222 =  ( n10221 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10223 =  ( n10220 ) ^ ( n10222 )  ;
assign n10224 =  ( n6483 ) | ( n6492 )  ;
assign n10225 =  ( n10224 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10226 =  ( n10223 ) ^ ( n10225 )  ;
assign n10227 = ~ ( n10226 ) ;
assign n10228 =  ( n6030 ) | ( n6039 )  ;
assign n10229 =  ( n10228 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10230 = ~ ( n10229 ) ;
assign n10231 =  ( n10227 ) | ( n10230 )  ;
assign n10232 = ~ ( n7809 ) ;
assign n10233 = ~ ( n9916 ) ;
assign n10234 =  ( n10232 ) | ( n10233 )  ;
assign n10235 =  ( n10140 ) ^ ( n10234 )  ;
assign n10236 =  ( n10235 ) ^ ( n7455 )  ;
assign n10237 =  ( n6825 ) | ( n6834 )  ;
assign n10238 =  ( n10237 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10239 =  ( n10236 ) ^ ( n10238 )  ;
assign n10240 =  ( n6483 ) | ( n6492 )  ;
assign n10241 =  ( n10240 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10242 =  ( n10239 ) ^ ( n10241 )  ;
assign n10243 =  ( n6030 ) | ( n6039 )  ;
assign n10244 =  ( n10243 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10245 =  ( n10242 ) ^ ( n10244 )  ;
assign n10246 =  ( n10245 ) ^ ( n9788 )  ;
assign n10247 =  ( n10246 ) ^ ( n9785 )  ;
assign n10248 = ~ ( n10247 ) ;
assign n10249 =  ( n10231 ) | ( n10248 )  ;
assign n10250 = ~ ( n10249 ) ;
assign n10251 = ~ ( n10226 ) ;
assign n10252 =  ( n6030 ) | ( n6039 )  ;
assign n10253 =  ( n10252 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10254 = ~ ( n10253 ) ;
assign n10255 =  ( n10251 ) | ( n10254 )  ;
assign n10256 = ~ ( n10255 ) ;
assign n10257 =  ( n10256 ) ^ ( n10140 )  ;
assign n10258 = ~ ( n7809 ) ;
assign n10259 = ~ ( n9916 ) ;
assign n10260 =  ( n10258 ) | ( n10259 )  ;
assign n10261 =  ( n10257 ) ^ ( n10260 )  ;
assign n10262 =  ( n10261 ) ^ ( n7455 )  ;
assign n10263 =  ( n6825 ) | ( n6834 )  ;
assign n10264 =  ( n10263 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10265 =  ( n10262 ) ^ ( n10264 )  ;
assign n10266 =  ( n6483 ) | ( n6492 )  ;
assign n10267 =  ( n10266 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10268 =  ( n10265 ) ^ ( n10267 )  ;
assign n10269 =  ( n6030 ) | ( n6039 )  ;
assign n10270 =  ( n10269 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10271 =  ( n10268 ) ^ ( n10270 )  ;
assign n10272 =  ( n10271 ) ^ ( n9788 )  ;
assign n10273 =  ( n10272 ) ^ ( n9785 )  ;
assign n10274 = ~ ( n10273 ) ;
assign n10275 = ~ ( n7809 ) ;
assign n10276 = ~ ( n9916 ) ;
assign n10277 =  ( n10275 ) | ( n10276 )  ;
assign n10278 = ~ ( n10277 ) ;
assign n10279 =  ( n10274 ) | ( n10278 )  ;
assign n10280 =  ( n6825 ) | ( n6834 )  ;
assign n10281 =  ( n10280 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10282 =  ( n7455 ) ^ ( n10281 )  ;
assign n10283 =  ( n6483 ) | ( n6492 )  ;
assign n10284 =  ( n10283 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10285 =  ( n10282 ) ^ ( n10284 )  ;
assign n10286 =  ( n10285 ) ^ ( n10084 )  ;
assign n10287 =  ( n10286 ) ^ ( n10081 )  ;
assign n10288 = ~ ( n10287 ) ;
assign n10289 =  ( n10279 ) | ( n10288 )  ;
assign n10290 = ~ ( n10086 ) ;
assign n10291 =  ( n7784 ) | ( n10091 )  ;
assign n10292 = ~ ( n10291 ) ;
assign n10293 =  ( n10290 ) | ( n10292 )  ;
assign n10294 =  ( n10293 ) | ( n10107 )  ;
assign n10295 = ~ ( n7809 ) ;
assign n10296 = ~ ( n10115 ) ;
assign n10297 =  ( n10295 ) | ( n10296 )  ;
assign n10298 =  ( n10294 ) ^ ( n10297 )  ;
assign n10299 =  ( n10298 ) ^ ( n7455 )  ;
assign n10300 =  ( n6825 ) | ( n6834 )  ;
assign n10301 =  ( n10300 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10302 =  ( n10299 ) ^ ( n10301 )  ;
assign n10303 =  ( n6483 ) | ( n6492 )  ;
assign n10304 =  ( n10303 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10305 =  ( n10302 ) ^ ( n10304 )  ;
assign n10306 =  ( n6030 ) | ( n6039 )  ;
assign n10307 =  ( n10306 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10308 =  ( n10305 ) ^ ( n10307 )  ;
assign n10309 = ~ ( n10308 ) ;
assign n10310 =  ( n10289 ) | ( n10309 )  ;
assign n10311 = ~ ( n10310 ) ;
assign n10312 =  ( n10250 ) | ( n10311 )  ;
assign n10313 = ~ ( n10312 ) ;
assign n10314 =  ( n10210 ) | ( n10313 )  ;
assign n10315 = ~ ( n10314 ) ;
assign n10316 =  ( n10183 ) | ( n10315 )  ;
assign n10317 = ~ ( n10316 ) ;
assign n10318 =  ( n9911 ) | ( n10317 )  ;
assign n10319 = ~ ( n10318 ) ;
assign n10320 =  ( n9872 ) | ( n10319 )  ;
assign n10321 = ~ ( n9432 ) ;
assign n10322 = ~ ( n9649 ) ;
assign n10323 =  ( n10321 ) | ( n10322 )  ;
assign n10324 = ~ ( n9751 ) ;
assign n10325 =  ( n10323 ) | ( n10324 )  ;
assign n10326 = ~ ( n9909 ) ;
assign n10327 =  ( n10325 ) | ( n10326 )  ;
assign n10328 = ~ ( n10042 ) ;
assign n10329 =  ( n10327 ) | ( n10328 )  ;
assign n10330 = ~ ( n10208 ) ;
assign n10331 =  ( n10329 ) | ( n10330 )  ;
assign n10332 =  ( n10331 ) | ( n10274 )  ;
assign n10333 = ~ ( n7809 ) ;
assign n10334 = ~ ( n9916 ) ;
assign n10335 =  ( n10333 ) | ( n10334 )  ;
assign n10336 = ~ ( n10335 ) ;
assign n10337 =  ( n10336 ) | ( n10288 )  ;
assign n10338 = ~ ( n10337 ) ;
assign n10339 = ~ ( n10086 ) ;
assign n10340 =  ( n7784 ) | ( n10091 )  ;
assign n10341 = ~ ( n10340 ) ;
assign n10342 =  ( n10339 ) | ( n10341 )  ;
assign n10343 =  ( n10342 ) | ( n10107 )  ;
assign n10344 =  ( n10338 ) ^ ( n10343 )  ;
assign n10345 = ~ ( n7809 ) ;
assign n10346 = ~ ( n10115 ) ;
assign n10347 =  ( n10345 ) | ( n10346 )  ;
assign n10348 =  ( n10344 ) ^ ( n10347 )  ;
assign n10349 =  ( n10348 ) ^ ( n7455 )  ;
assign n10350 =  ( n6825 ) | ( n6834 )  ;
assign n10351 =  ( n10350 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10352 =  ( n10349 ) ^ ( n10351 )  ;
assign n10353 =  ( n6483 ) | ( n6492 )  ;
assign n10354 =  ( n10353 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10355 =  ( n10352 ) ^ ( n10354 )  ;
assign n10356 =  ( n6030 ) | ( n6039 )  ;
assign n10357 =  ( n10356 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n10358 =  ( n10355 ) ^ ( n10357 )  ;
assign n10359 = ~ ( n10358 ) ;
assign n10360 =  ( n10332 ) | ( n10359 )  ;
assign n10361 = ~ ( n7809 ) ;
assign n10362 = kd[5:5] ;
assign n10363 =  ( n10362 ) == ( bv_1_0_n2 )  ;
assign n10364 = kd[4:4] ;
assign n10365 =  ( n10364 ) == ( bv_1_1_n5 )  ;
assign n10366 =  ( n10363 ) | ( n10365 )  ;
assign n10367 = kd[3:3] ;
assign n10368 =  ( n10367 ) == ( bv_1_1_n5 )  ;
assign n10369 =  ( n10366 ) | ( n10368 )  ;
assign n10370 = ~ ( n10369 )  ;
assign n10371 = kd[5:5] ;
assign n10372 =  ( n10371 ) == ( bv_1_1_n5 )  ;
assign n10373 = kd[4:4] ;
assign n10374 =  ( n10373 ) == ( bv_1_0_n2 )  ;
assign n10375 =  ( n10372 ) | ( n10374 )  ;
assign n10376 = kd[3:3] ;
assign n10377 =  ( n10376 ) == ( bv_1_0_n2 )  ;
assign n10378 =  ( n10375 ) | ( n10377 )  ;
assign n10379 = ~ ( n10378 )  ;
assign n10380 =  ( n10370 ) | ( n10379 )  ;
assign n10381 = kd[5:5] ;
assign n10382 = ~ ( n10381 ) ;
assign n10383 = kd[4:4] ;
assign n10384 = ~ ( n10383 ) ;
assign n10385 = kd[3:3] ;
assign n10386 = ~ ( n10385 ) ;
assign n10387 =  ( n10384 ) | ( n10386 )  ;
assign n10388 = ~ ( n10387 ) ;
assign n10389 =  ( n10382 ) | ( n10388 )  ;
assign n10390 = ~ ( n10389 ) ;
assign n10391 =  ( n6483 ) | ( n6492 )  ;
assign n10392 =  ( n10391 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10393 =  ( n10380 ) ? ( n10390 ) : ( n10392 ) ;
assign n10394 = ~ ( n10393 ) ;
assign n10395 =  ( n7784 ) | ( n10394 )  ;
assign n10396 = ~ ( n10395 ) ;
assign n10397 =  ( n10361 ) | ( n10396 )  ;
assign n10398 = ~ ( n10397 ) ;
assign n10399 =  ( n10398 ) | ( n10137 )  ;
assign n10400 = ~ ( n7809 ) ;
assign n10401 = ~ ( n9916 ) ;
assign n10402 =  ( n10400 ) | ( n10401 )  ;
assign n10403 =  ( n10402 ) ^ ( n7455 )  ;
assign n10404 =  ( n6825 ) | ( n6834 )  ;
assign n10405 =  ( n10404 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10406 =  ( n10403 ) ^ ( n10405 )  ;
assign n10407 =  ( n6483 ) | ( n6492 )  ;
assign n10408 =  ( n10407 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10409 =  ( n10406 ) ^ ( n10408 )  ;
assign n10410 =  ( n10409 ) ^ ( n10084 )  ;
assign n10411 =  ( n10410 ) ^ ( n10081 )  ;
assign n10412 = ~ ( n10411 ) ;
assign n10413 =  ( n10399 ) | ( n10412 )  ;
assign n10414 = ~ ( n10413 ) ;
assign n10415 = ~ ( n10397 ) ;
assign n10416 =  ( n10415 ) | ( n10137 )  ;
assign n10417 = ~ ( n10416 ) ;
assign n10418 = ~ ( n7809 ) ;
assign n10419 = ~ ( n9916 ) ;
assign n10420 =  ( n10418 ) | ( n10419 )  ;
assign n10421 =  ( n10417 ) ^ ( n10420 )  ;
assign n10422 =  ( n10421 ) ^ ( n7455 )  ;
assign n10423 =  ( n6825 ) | ( n6834 )  ;
assign n10424 =  ( n10423 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10425 =  ( n10422 ) ^ ( n10424 )  ;
assign n10426 =  ( n6483 ) | ( n6492 )  ;
assign n10427 =  ( n10426 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10428 =  ( n10425 ) ^ ( n10427 )  ;
assign n10429 =  ( n10428 ) ^ ( n10084 )  ;
assign n10430 =  ( n10429 ) ^ ( n10081 )  ;
assign n10431 = ~ ( n10430 ) ;
assign n10432 =  ( n6825 ) | ( n6834 )  ;
assign n10433 =  ( n10432 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10434 =  ( n7455 ) ^ ( n10433 )  ;
assign n10435 =  ( n10434 ) ^ ( n10393 )  ;
assign n10436 = ~ ( n10435 ) ;
assign n10437 =  ( n10431 ) | ( n10436 )  ;
assign n10438 = kd[5:5] ;
assign n10439 = ~ ( n10438 ) ;
assign n10440 =  ( n10437 ) | ( n10439 )  ;
assign n10441 =  ( n10440 ) | ( n10388 )  ;
assign n10442 =  ( n10397 ) ^ ( n7455 )  ;
assign n10443 =  ( n6825 ) | ( n6834 )  ;
assign n10444 =  ( n10443 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10445 =  ( n10442 ) ^ ( n10444 )  ;
assign n10446 =  ( n6483 ) | ( n6492 )  ;
assign n10447 =  ( n10446 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10448 =  ( n10445 ) ^ ( n10447 )  ;
assign n10449 = ~ ( n10448 ) ;
assign n10450 =  ( n10441 ) | ( n10449 )  ;
assign n10451 = ~ ( n10450 ) ;
assign n10452 =  ( n10414 ) | ( n10451 )  ;
assign n10453 = ~ ( n10430 ) ;
assign n10454 = kd[5:5] ;
assign n10455 = ~ ( n10454 ) ;
assign n10456 =  ( n10436 ) | ( n10455 )  ;
assign n10457 =  ( n10456 ) | ( n10388 )  ;
assign n10458 = ~ ( n10457 ) ;
assign n10459 =  ( n10458 ) ^ ( n10397 )  ;
assign n10460 =  ( n10459 ) ^ ( n7455 )  ;
assign n10461 =  ( n6825 ) | ( n6834 )  ;
assign n10462 =  ( n10461 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10463 =  ( n10460 ) ^ ( n10462 )  ;
assign n10464 =  ( n6483 ) | ( n6492 )  ;
assign n10465 =  ( n10464 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n10466 =  ( n10463 ) ^ ( n10465 )  ;
assign n10467 = ~ ( n10466 ) ;
assign n10468 =  ( n10453 ) | ( n10467 )  ;
assign n10469 = ~ ( n7455 ) ;
assign n10470 =  ( n6825 ) | ( n6834 )  ;
assign n10471 =  ( n10470 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10472 = ~ ( n10471 ) ;
assign n10473 =  ( n10469 ) | ( n10472 )  ;
assign n10474 =  ( n6825 ) | ( n6834 )  ;
assign n10475 =  ( n10474 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10476 =  ( n7455 ) ^ ( n10475 )  ;
assign n10477 =  ( n10476 ) ^ ( n10393 )  ;
assign n10478 =  ( n10477 ) ^ ( n10390 )  ;
assign n10479 = ~ ( n10478 ) ;
assign n10480 =  ( n10473 ) | ( n10479 )  ;
assign n10481 = ~ ( n10480 ) ;
assign n10482 = ~ ( n7809 ) ;
assign n10483 =  ( n10482 ) ^ ( n7455 )  ;
assign n10484 =  ( n6825 ) | ( n6834 )  ;
assign n10485 =  ( n10484 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10486 =  ( n10483 ) ^ ( n10485 )  ;
assign n10487 =  ( n10486 ) ^ ( n10393 )  ;
assign n10488 =  ( n10487 ) ^ ( n10390 )  ;
assign n10489 = ~ ( n10488 ) ;
assign n10490 = ~ ( n7455 ) ;
assign n10491 = kd[3:3] ;
assign n10492 =  ( n10491 ) == ( bv_1_0_n2 )  ;
assign n10493 = kd[2:2] ;
assign n10494 =  ( n10493 ) == ( bv_1_1_n5 )  ;
assign n10495 =  ( n10492 ) | ( n10494 )  ;
assign n10496 = kd[1:1] ;
assign n10497 =  ( n10496 ) == ( bv_1_1_n5 )  ;
assign n10498 =  ( n10495 ) | ( n10497 )  ;
assign n10499 = ~ ( n10498 )  ;
assign n10500 = kd[3:3] ;
assign n10501 =  ( n10500 ) == ( bv_1_1_n5 )  ;
assign n10502 = kd[2:2] ;
assign n10503 =  ( n10502 ) == ( bv_1_0_n2 )  ;
assign n10504 =  ( n10501 ) | ( n10503 )  ;
assign n10505 = kd[1:1] ;
assign n10506 =  ( n10505 ) == ( bv_1_0_n2 )  ;
assign n10507 =  ( n10504 ) | ( n10506 )  ;
assign n10508 = ~ ( n10507 )  ;
assign n10509 =  ( n10499 ) | ( n10508 )  ;
assign n10510 = kd[3:3] ;
assign n10511 = ~ ( n10510 ) ;
assign n10512 = kd[2:2] ;
assign n10513 = ~ ( n10512 ) ;
assign n10514 = kd[1:1] ;
assign n10515 = ~ ( n10514 ) ;
assign n10516 =  ( n10513 ) | ( n10515 )  ;
assign n10517 = ~ ( n10516 ) ;
assign n10518 =  ( n10511 ) | ( n10517 )  ;
assign n10519 = ~ ( n10518 ) ;
assign n10520 =  ( n6825 ) | ( n6834 )  ;
assign n10521 =  ( n10520 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10522 =  ( n10509 ) ? ( n10519 ) : ( n10521 ) ;
assign n10523 = ~ ( n10522 ) ;
assign n10524 =  ( n10490 ) | ( n10523 )  ;
assign n10525 = ~ ( n10524 ) ;
assign n10526 =  ( n7455 ) ^ ( n10522 )  ;
assign n10527 = ~ ( n10526 ) ;
assign n10528 = kd[3:3] ;
assign n10529 = ~ ( n10528 ) ;
assign n10530 =  ( n10527 ) | ( n10529 )  ;
assign n10531 =  ( n10530 ) | ( n10517 )  ;
assign n10532 = ~ ( n10531 ) ;
assign n10533 =  ( n10525 ) | ( n10532 )  ;
assign n10534 = ~ ( n10533 ) ;
assign n10535 =  ( n10489 ) | ( n10534 )  ;
assign n10536 =  ( n10535 ) | ( n7784 )  ;
assign n10537 = ~ ( n10536 ) ;
assign n10538 =  ( n10481 ) | ( n10537 )  ;
assign n10539 = ~ ( n10538 ) ;
assign n10540 =  ( n10468 ) | ( n10539 )  ;
assign n10541 = ~ ( n10540 ) ;
assign n10542 =  ( n10452 ) | ( n10541 )  ;
assign n10543 = ~ ( n10430 ) ;
assign n10544 =  ( n10543 ) | ( n10467 )  ;
assign n10545 =  ( n10544 ) | ( n10489 )  ;
assign n10546 =  ( n10533 ) ^ ( n7455 )  ;
assign n10547 =  ( n6825 ) | ( n6834 )  ;
assign n10548 =  ( n10547 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n10549 =  ( n10546 ) ^ ( n10548 )  ;
assign n10550 = ~ ( n10549 ) ;
assign n10551 =  ( n10545 ) | ( n10550 )  ;
assign n10552 =  ( n7455 ) ^ ( n10522 )  ;
assign n10553 =  ( n10552 ) ^ ( n10519 )  ;
assign n10554 = ~ ( n10553 ) ;
assign n10555 =  ( n10551 ) | ( n10554 )  ;
assign n10556 = ~ ( n7455 ) ;
assign n10557 =  ( n10555 ) | ( n10556 )  ;
assign n10558 = kd[0:0] ;
assign n10559 =  ( n10558 ) == ( bv_1_1_n5 )  ;
assign n10560 = kd[1:1] ;
assign n10561 =  ( n10560 ) == ( bv_1_0_n2 )  ;
assign n10562 =  ( n10559 ) | ( n10561 )  ;
assign n10563 = kd[1:1] ;
assign n10564 =  ( n10562 ) ? ( n7455 ) : ( n10563 ) ;
assign n10565 = ~ ( n10564 ) ;
assign n10566 =  ( n10557 ) | ( n10565 )  ;
assign n10567 = kd[1:1] ;
assign n10568 = ~ ( n10567 ) ;
assign n10569 =  ( n10566 ) | ( n10568 )  ;
assign n10570 = ~ ( n10569 ) ;
assign n10571 =  ( n10542 ) | ( n10570 )  ;
assign n10572 = ~ ( n10571 ) ;
assign n10573 =  ( n10360 ) | ( n10572 )  ;
assign n10574 = ~ ( n10573 ) ;
assign n10575 =  ( n10320 ) | ( n10574 )  ;
assign n10576 = ~ ( n10575 ) ;
assign n10577 =  ( n9254 ) | ( n10576 )  ;
assign n10578 = ~ ( n10577 ) ;
assign n10579 =  ( n9184 ) | ( n10578 )  ;
assign n10580 = ~ ( n10579 ) ;
assign n10581 =  ( n5673 ) ^ ( n10580 )  ;
assign n10582 =  ( n373 ) | ( n382 )  ;
assign n10583 =  ( n10582 ) ? ( bv_1_0_n2 ) : ( n502 ) ;
assign n10584 = ~ ( n10583 ) ;
assign n10585 =  ( n509 ) ^ ( n10584 )  ;
assign n10586 =  ( bv_1_1_n5 ) ^ ( n488 )  ;
assign n10587 =  ( n10586 ) ^ ( n504 )  ;
assign n10588 = ~ ( n10587 ) ;
assign n10589 = ~ ( n834 ) ;
assign n10590 = ~ ( n841 ) ;
assign n10591 =  ( n10589 ) | ( n10590 )  ;
assign n10592 = ~ ( n10591 ) ;
assign n10593 = ~ ( n856 ) ;
assign n10594 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n10595 =  ( n10594 ) ^ ( n823 )  ;
assign n10596 =  ( n10595 ) ^ ( n344 )  ;
assign n10597 =  ( n10596 ) ^ ( n454 )  ;
assign n10598 = ~ ( n10597 ) ;
assign n10599 =  ( n10593 ) | ( n10598 )  ;
assign n10600 = ~ ( n1212 ) ;
assign n10601 =  ( n10599 ) | ( n10600 )  ;
assign n10602 = ~ ( n1224 ) ;
assign n10603 =  ( n10601 ) | ( n10602 )  ;
assign n10604 = ~ ( n10603 ) ;
assign n10605 =  ( n10592 ) | ( n10604 )  ;
assign n10606 = ~ ( n856 ) ;
assign n10607 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n10608 =  ( n10607 ) ^ ( n823 )  ;
assign n10609 =  ( n10608 ) ^ ( n344 )  ;
assign n10610 =  ( n10609 ) ^ ( n454 )  ;
assign n10611 = ~ ( n10610 ) ;
assign n10612 =  ( n10606 ) | ( n10611 )  ;
assign n10613 = ~ ( n1239 ) ;
assign n10614 =  ( n10612 ) | ( n10613 )  ;
assign n10615 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n10616 =  ( n10615 ) ^ ( n1199 )  ;
assign n10617 =  ( n10616 ) ^ ( n666 )  ;
assign n10618 =  ( n10617 ) ^ ( n682 )  ;
assign n10619 =  ( n10618 ) ^ ( n697 )  ;
assign n10620 =  ( n10619 ) ^ ( n759 )  ;
assign n10621 = ~ ( n10620 ) ;
assign n10622 =  ( n10614 ) | ( n10621 )  ;
assign n10623 = ~ ( n1446 ) ;
assign n10624 = ~ ( n1773 ) ;
assign n10625 =  ( n10623 ) | ( n10624 )  ;
assign n10626 =  ( n10625 ) | ( n1783 )  ;
assign n10627 = ~ ( n10626 ) ;
assign n10628 =  ( n1426 ) | ( n10627 )  ;
assign n10629 = ~ ( n1446 ) ;
assign n10630 =  ( n10629 ) | ( n1828 )  ;
assign n10631 = ~ ( n2070 ) ;
assign n10632 =  ( n10631 ) | ( n2080 )  ;
assign n10633 = ~ ( n2092 ) ;
assign n10634 =  ( n10632 ) | ( n10633 )  ;
assign n10635 = ~ ( n10634 ) ;
assign n10636 = ~ ( n2110 ) ;
assign n10637 = ~ ( n2426 ) ;
assign n10638 =  ( n10636 ) | ( n10637 )  ;
assign n10639 =  ( n10638 ) | ( n2438 )  ;
assign n10640 = ~ ( n10639 ) ;
assign n10641 =  ( n10635 ) | ( n10640 )  ;
assign n10642 = ~ ( n10641 ) ;
assign n10643 =  ( n10630 ) | ( n10642 )  ;
assign n10644 = ~ ( n10643 ) ;
assign n10645 =  ( n10628 ) | ( n10644 )  ;
assign n10646 = ~ ( n10645 ) ;
assign n10647 =  ( n10622 ) | ( n10646 )  ;
assign n10648 = ~ ( n10647 ) ;
assign n10649 =  ( n10605 ) | ( n10648 )  ;
assign n10650 = ~ ( n856 ) ;
assign n10651 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n10652 =  ( n10651 ) ^ ( n823 )  ;
assign n10653 =  ( n10652 ) ^ ( n344 )  ;
assign n10654 =  ( n10653 ) ^ ( n454 )  ;
assign n10655 = ~ ( n10654 ) ;
assign n10656 =  ( n10650 ) | ( n10655 )  ;
assign n10657 = ~ ( n1239 ) ;
assign n10658 =  ( n10656 ) | ( n10657 )  ;
assign n10659 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n10660 =  ( n10659 ) ^ ( n1199 )  ;
assign n10661 =  ( n10660 ) ^ ( n666 )  ;
assign n10662 =  ( n10661 ) ^ ( n682 )  ;
assign n10663 =  ( n10662 ) ^ ( n697 )  ;
assign n10664 =  ( n10663 ) ^ ( n759 )  ;
assign n10665 = ~ ( n10664 ) ;
assign n10666 =  ( n10658 ) | ( n10665 )  ;
assign n10667 = ~ ( n1446 ) ;
assign n10668 =  ( n10666 ) | ( n10667 )  ;
assign n10669 =  ( n10668 ) | ( n1828 )  ;
assign n10670 = ~ ( n2110 ) ;
assign n10671 =  ( n10669 ) | ( n10670 )  ;
assign n10672 =  ( n10671 ) | ( n2453 )  ;
assign n10673 = ~ ( n2722 ) ;
assign n10674 = ~ ( n2742 ) ;
assign n10675 = ~ ( n3043 ) ;
assign n10676 =  ( n10674 ) | ( n10675 )  ;
assign n10677 =  ( n10676 ) | ( n3059 )  ;
assign n10678 = ~ ( n10677 ) ;
assign n10679 =  ( n10673 ) | ( n10678 )  ;
assign n10680 = ~ ( n2742 ) ;
assign n10681 =  ( n10680 ) | ( n3085 )  ;
assign n10682 = ~ ( n3366 ) ;
assign n10683 = ~ ( n3392 ) ;
assign n10684 = ~ ( n3623 ) ;
assign n10685 =  ( n10683 ) | ( n10684 )  ;
assign n10686 =  ( n10685 ) | ( n3646 )  ;
assign n10687 = ~ ( n10686 ) ;
assign n10688 =  ( n10682 ) | ( n10687 )  ;
assign n10689 = ~ ( n10688 ) ;
assign n10690 =  ( n10681 ) | ( n10689 )  ;
assign n10691 = ~ ( n10690 ) ;
assign n10692 =  ( n10679 ) | ( n10691 )  ;
assign n10693 = ~ ( n2742 ) ;
assign n10694 =  ( n10693 ) | ( n3085 )  ;
assign n10695 = ~ ( n3392 ) ;
assign n10696 =  ( n10694 ) | ( n10695 )  ;
assign n10697 =  ( n10696 ) | ( n3672 )  ;
assign n10698 = ~ ( n3958 ) ;
assign n10699 =  ( n10698 ) | ( n4181 )  ;
assign n10700 =  ( n3985 ) | ( n4253 )  ;
assign n10701 = ~ ( n4435 ) ;
assign n10702 = ~ ( n4689 ) ;
assign n10703 =  ( n10701 ) | ( n10702 )  ;
assign n10704 = ~ ( n10703 ) ;
assign n10705 =  ( n10700 ) | ( n10704 )  ;
assign n10706 = ~ ( n10705 ) ;
assign n10707 =  ( n10699 ) | ( n10706 )  ;
assign n10708 = ~ ( n10707 ) ;
assign n10709 =  ( n10697 ) | ( n10708 )  ;
assign n10710 = ~ ( n10709 ) ;
assign n10711 =  ( n10692 ) | ( n10710 )  ;
assign n10712 = ~ ( n10711 ) ;
assign n10713 =  ( n10672 ) | ( n10712 )  ;
assign n10714 = ~ ( n10713 ) ;
assign n10715 =  ( n10649 ) | ( n10714 )  ;
assign n10716 = ~ ( n856 ) ;
assign n10717 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n10718 =  ( n10717 ) ^ ( n823 )  ;
assign n10719 =  ( n10718 ) ^ ( n344 )  ;
assign n10720 =  ( n10719 ) ^ ( n454 )  ;
assign n10721 = ~ ( n10720 ) ;
assign n10722 =  ( n10716 ) | ( n10721 )  ;
assign n10723 = ~ ( n1239 ) ;
assign n10724 =  ( n10722 ) | ( n10723 )  ;
assign n10725 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n10726 =  ( n10725 ) ^ ( n1199 )  ;
assign n10727 =  ( n10726 ) ^ ( n666 )  ;
assign n10728 =  ( n10727 ) ^ ( n682 )  ;
assign n10729 =  ( n10728 ) ^ ( n697 )  ;
assign n10730 =  ( n10729 ) ^ ( n759 )  ;
assign n10731 = ~ ( n10730 ) ;
assign n10732 =  ( n10724 ) | ( n10731 )  ;
assign n10733 = ~ ( n1446 ) ;
assign n10734 =  ( n10732 ) | ( n10733 )  ;
assign n10735 =  ( n10734 ) | ( n1828 )  ;
assign n10736 = ~ ( n2110 ) ;
assign n10737 =  ( n10735 ) | ( n10736 )  ;
assign n10738 =  ( n10737 ) | ( n2453 )  ;
assign n10739 = ~ ( n2742 ) ;
assign n10740 =  ( n10738 ) | ( n10739 )  ;
assign n10741 =  ( n10740 ) | ( n3085 )  ;
assign n10742 = ~ ( n3392 ) ;
assign n10743 =  ( n10741 ) | ( n10742 )  ;
assign n10744 =  ( n10743 ) | ( n3672 )  ;
assign n10745 =  ( n10744 ) | ( n3985 )  ;
assign n10746 =  ( n10745 ) | ( n4253 )  ;
assign n10747 =  ( n10746 ) | ( n4458 )  ;
assign n10748 =  ( n10747 ) | ( n4710 )  ;
assign n10749 = ~ ( n4728 ) ;
assign n10750 =  ( n4722 ) | ( n10749 )  ;
assign n10751 =  ( n10750 ) | ( n4744 )  ;
assign n10752 = ~ ( n10751 ) ;
assign n10753 = ~ ( n4763 ) ;
assign n10754 = ~ ( n4889 ) ;
assign n10755 =  ( n10753 ) | ( n10754 )  ;
assign n10756 =  ( n10755 ) | ( n4900 )  ;
assign n10757 =  ( n10756 ) | ( n4913 )  ;
assign n10758 = ~ ( n10757 ) ;
assign n10759 =  ( n10752 ) | ( n10758 )  ;
assign n10760 = ~ ( n4763 ) ;
assign n10761 = ~ ( n4938 ) ;
assign n10762 =  ( n10760 ) | ( n10761 )  ;
assign n10763 =  ( n5041 ) | ( n5203 )  ;
assign n10764 = ~ ( n10763 ) ;
assign n10765 =  ( n10762 ) | ( n10764 )  ;
assign n10766 = ~ ( n10765 ) ;
assign n10767 =  ( n10759 ) | ( n10766 )  ;
assign n10768 = ~ ( n4763 ) ;
assign n10769 = ~ ( n4938 ) ;
assign n10770 =  ( n10768 ) | ( n10769 )  ;
assign n10771 =  ( n10770 ) | ( n5063 )  ;
assign n10772 =  ( n10771 ) | ( n5224 )  ;
assign n10773 =  ( n5248 ) | ( n5341 )  ;
assign n10774 =  ( n5366 ) ^ ( n5161 )  ;
assign n10775 =  ( n10774 ) ^ ( n5171 )  ;
assign n10776 =  ( n10775 ) ^ ( n4960 )  ;
assign n10777 =  ( n10776 ) ^ ( n4976 )  ;
assign n10778 =  ( n10777 ) ^ ( n4996 )  ;
assign n10779 =  ( n10778 ) ^ ( n5236 )  ;
assign n10780 = ~ ( n10779 ) ;
assign n10781 =  ( n5265 ) | ( n10780 )  ;
assign n10782 =  ( n5446 ) | ( n5473 )  ;
assign n10783 = ~ ( n10782 ) ;
assign n10784 =  ( n10781 ) | ( n10783 )  ;
assign n10785 = ~ ( n10784 ) ;
assign n10786 =  ( n10773 ) | ( n10785 )  ;
assign n10787 = ~ ( n10786 ) ;
assign n10788 =  ( n10772 ) | ( n10787 )  ;
assign n10789 = ~ ( n10788 ) ;
assign n10790 =  ( n10767 ) | ( n10789 )  ;
assign n10791 = ~ ( n4763 ) ;
assign n10792 = ~ ( n4938 ) ;
assign n10793 =  ( n10791 ) | ( n10792 )  ;
assign n10794 =  ( n10793 ) | ( n5063 )  ;
assign n10795 =  ( n10794 ) | ( n5224 )  ;
assign n10796 =  ( n10795 ) | ( n5265 )  ;
assign n10797 =  ( n5366 ) ^ ( n5161 )  ;
assign n10798 =  ( n10797 ) ^ ( n5171 )  ;
assign n10799 =  ( n10798 ) ^ ( n4960 )  ;
assign n10800 =  ( n10799 ) ^ ( n4976 )  ;
assign n10801 =  ( n10800 ) ^ ( n4996 )  ;
assign n10802 =  ( n10801 ) ^ ( n5236 )  ;
assign n10803 = ~ ( n10802 ) ;
assign n10804 =  ( n10796 ) | ( n10803 )  ;
assign n10805 =  ( n5452 ) ^ ( n5325 )  ;
assign n10806 =  ( n10805 ) ^ ( n5083 )  ;
assign n10807 =  ( n10806 ) ^ ( n5099 )  ;
assign n10808 =  ( n10807 ) ^ ( n5116 )  ;
assign n10809 =  ( n10808 ) ^ ( n5141 )  ;
assign n10810 =  ( n10809 ) ^ ( n5129 )  ;
assign n10811 = ~ ( n10810 ) ;
assign n10812 =  ( n10804 ) | ( n10811 )  ;
assign n10813 =  ( n5489 ) ^ ( n5433 )  ;
assign n10814 =  ( n10813 ) ^ ( n5285 )  ;
assign n10815 =  ( n10814 ) ^ ( n5301 )  ;
assign n10816 =  ( n10815 ) ^ ( n5321 )  ;
assign n10817 = ~ ( n10816 ) ;
assign n10818 =  ( n10812 ) | ( n10817 )  ;
assign n10819 =  ( n5539 ) | ( n5600 )  ;
assign n10820 = ~ ( n5547 ) ;
assign n10821 =  ( n5594 ) ^ ( n5515 )  ;
assign n10822 =  ( n10821 ) ^ ( n5531 )  ;
assign n10823 = ~ ( n10822 ) ;
assign n10824 =  ( n10820 ) | ( n10823 )  ;
assign n10825 =  ( n5568 ) ^ ( n5583 )  ;
assign n10826 =  ( n10825 ) ^ ( n5580 )  ;
assign n10827 = ~ ( n10826 ) ;
assign n10828 =  ( n10824 ) | ( n10827 )  ;
assign n10829 = ~ ( n5648 ) ;
assign n10830 =  ( n10828 ) | ( n10829 )  ;
assign n10831 = ~ ( n5657 ) ;
assign n10832 =  ( n10830 ) | ( n10831 )  ;
assign n10833 = ki[1:1] ;
assign n10834 = ~ ( n10833 ) ;
assign n10835 =  ( n10832 ) | ( n10834 )  ;
assign n10836 = ~ ( n10835 ) ;
assign n10837 =  ( n10819 ) | ( n10836 )  ;
assign n10838 = ~ ( n10837 ) ;
assign n10839 =  ( n10818 ) | ( n10838 )  ;
assign n10840 = ~ ( n10839 ) ;
assign n10841 =  ( n10790 ) | ( n10840 )  ;
assign n10842 = ~ ( n10841 ) ;
assign n10843 =  ( n10748 ) | ( n10842 )  ;
assign n10844 = ~ ( n10843 ) ;
assign n10845 =  ( n10715 ) | ( n10844 )  ;
assign n10846 = ~ ( n10845 ) ;
assign n10847 =  ( n10588 ) | ( n10846 )  ;
assign n10848 = ~ ( n10847 ) ;
assign n10849 =  ( n10585 ) ^ ( n10848 )  ;
assign n10850 = ~ ( n10849 ) ;
assign n10851 =  ( n5713 ) | ( n5722 )  ;
assign n10852 =  ( n10851 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n10853 = ~ ( n10852 ) ;
assign n10854 =  ( n5774 ) ^ ( n10853 )  ;
assign n10855 = ~ ( n5986 ) ;
assign n10856 =  ( n5976 ) | ( n10855 )  ;
assign n10857 = ~ ( n10856 ) ;
assign n10858 = ~ ( n6006 ) ;
assign n10859 =  ( n10858 ) | ( n6020 )  ;
assign n10860 = ~ ( n6264 ) ;
assign n10861 =  ( n10859 ) | ( n10860 )  ;
assign n10862 = ~ ( n6279 ) ;
assign n10863 =  ( n10861 ) | ( n10862 )  ;
assign n10864 = ~ ( n10863 ) ;
assign n10865 =  ( n10857 ) | ( n10864 )  ;
assign n10866 = ~ ( n6006 ) ;
assign n10867 =  ( n10866 ) | ( n6020 )  ;
assign n10868 = ~ ( n6297 ) ;
assign n10869 =  ( n10867 ) | ( n10868 )  ;
assign n10870 =  ( n10869 ) | ( n6314 )  ;
assign n10871 = ~ ( n6402 ) ;
assign n10872 =  ( n10871 ) | ( n6421 )  ;
assign n10873 = ~ ( n6444 ) ;
assign n10874 =  ( n10872 ) | ( n10873 )  ;
assign n10875 = ~ ( n10874 ) ;
assign n10876 = ~ ( n6473 ) ;
assign n10877 = ~ ( n6753 ) ;
assign n10878 =  ( n10876 ) | ( n10877 )  ;
assign n10879 =  ( n10878 ) | ( n6774 )  ;
assign n10880 = ~ ( n10879 ) ;
assign n10881 =  ( n10875 ) | ( n10880 )  ;
assign n10882 = ~ ( n6473 ) ;
assign n10883 =  ( n10882 ) | ( n6815 )  ;
assign n10884 = ~ ( n7022 ) ;
assign n10885 =  ( n10884 ) | ( n7045 )  ;
assign n10886 = ~ ( n7078 ) ;
assign n10887 =  ( n10885 ) | ( n10886 )  ;
assign n10888 = ~ ( n10887 ) ;
assign n10889 = ~ ( n7117 ) ;
assign n10890 = ~ ( n7392 ) ;
assign n10891 =  ( n10889 ) | ( n10890 )  ;
assign n10892 =  ( n10891 ) | ( n7417 )  ;
assign n10893 = ~ ( n10892 ) ;
assign n10894 =  ( n10888 ) | ( n10893 )  ;
assign n10895 = ~ ( n10894 ) ;
assign n10896 =  ( n10883 ) | ( n10895 )  ;
assign n10897 = ~ ( n10896 ) ;
assign n10898 =  ( n10881 ) | ( n10897 )  ;
assign n10899 = ~ ( n10898 ) ;
assign n10900 =  ( n10870 ) | ( n10899 )  ;
assign n10901 = ~ ( n10900 ) ;
assign n10902 =  ( n10865 ) | ( n10901 )  ;
assign n10903 = ~ ( n6006 ) ;
assign n10904 =  ( n10903 ) | ( n6020 )  ;
assign n10905 = ~ ( n6297 ) ;
assign n10906 =  ( n10904 ) | ( n10905 )  ;
assign n10907 =  ( n10906 ) | ( n6314 )  ;
assign n10908 = ~ ( n6473 ) ;
assign n10909 =  ( n10907 ) | ( n10908 )  ;
assign n10910 =  ( n10909 ) | ( n6815 )  ;
assign n10911 = ~ ( n7117 ) ;
assign n10912 =  ( n10910 ) | ( n10911 )  ;
assign n10913 =  ( n10912 ) | ( n7445 )  ;
assign n10914 = ~ ( n7649 ) ;
assign n10915 =  ( n10914 ) | ( n7679 )  ;
assign n10916 = ~ ( n7719 ) ;
assign n10917 =  ( n10915 ) | ( n10916 )  ;
assign n10918 = ~ ( n10917 ) ;
assign n10919 = ~ ( n7765 ) ;
assign n10920 = ~ ( n8047 ) ;
assign n10921 =  ( n10919 ) | ( n10920 )  ;
assign n10922 =  ( n10921 ) | ( n8079 )  ;
assign n10923 = ~ ( n10922 ) ;
assign n10924 =  ( n10918 ) | ( n10923 )  ;
assign n10925 = ~ ( n7765 ) ;
assign n10926 =  ( n10925 ) | ( n8121 )  ;
assign n10927 = ~ ( n8279 ) ;
assign n10928 = ~ ( n8321 ) ;
assign n10929 =  ( n10927 ) | ( n10928 )  ;
assign n10930 = ~ ( n8364 ) ;
assign n10931 =  ( n10929 ) | ( n10930 )  ;
assign n10932 = ~ ( n10931 ) ;
assign n10933 = ~ ( n8413 ) ;
assign n10934 = ~ ( n8625 ) ;
assign n10935 =  ( n10933 ) | ( n10934 )  ;
assign n10936 = ~ ( n8669 ) ;
assign n10937 =  ( n10935 ) | ( n10936 )  ;
assign n10938 = ~ ( n10937 ) ;
assign n10939 =  ( n10932 ) | ( n10938 )  ;
assign n10940 = ~ ( n10939 ) ;
assign n10941 =  ( n10926 ) | ( n10940 )  ;
assign n10942 = ~ ( n10941 ) ;
assign n10943 =  ( n10924 ) | ( n10942 )  ;
assign n10944 = ~ ( n7765 ) ;
assign n10945 =  ( n10944 ) | ( n8121 )  ;
assign n10946 = ~ ( n8413 ) ;
assign n10947 =  ( n10945 ) | ( n10946 )  ;
assign n10948 = ~ ( n8717 ) ;
assign n10949 =  ( n10947 ) | ( n10948 )  ;
assign n10950 = ~ ( n8880 ) ;
assign n10951 = ~ ( n8920 ) ;
assign n10952 =  ( n10950 ) | ( n10951 )  ;
assign n10953 = ~ ( n8963 ) ;
assign n10954 =  ( n10952 ) | ( n10953 )  ;
assign n10955 = ~ ( n10954 ) ;
assign n10956 =  ( n10955 ) | ( n9171 )  ;
assign n10957 = ~ ( n9012 ) ;
assign n10958 = ~ ( n9252 ) ;
assign n10959 =  ( n10957 ) | ( n10958 )  ;
assign n10960 = ~ ( n9314 ) ;
assign n10961 = ~ ( n9348 ) ;
assign n10962 =  ( n10960 ) | ( n10961 )  ;
assign n10963 = ~ ( n9387 ) ;
assign n10964 =  ( n10962 ) | ( n10963 )  ;
assign n10965 = ~ ( n10964 ) ;
assign n10966 =  ( n10965 ) | ( n9608 )  ;
assign n10967 = ~ ( n10966 ) ;
assign n10968 =  ( n10959 ) | ( n10967 )  ;
assign n10969 = ~ ( n10968 ) ;
assign n10970 =  ( n10956 ) | ( n10969 )  ;
assign n10971 = ~ ( n10970 ) ;
assign n10972 =  ( n10949 ) | ( n10971 )  ;
assign n10973 = ~ ( n10972 ) ;
assign n10974 =  ( n10943 ) | ( n10973 )  ;
assign n10975 = ~ ( n10974 ) ;
assign n10976 =  ( n10913 ) | ( n10975 )  ;
assign n10977 = ~ ( n10976 ) ;
assign n10978 =  ( n10902 ) | ( n10977 )  ;
assign n10979 = ~ ( n6006 ) ;
assign n10980 =  ( n10979 ) | ( n6020 )  ;
assign n10981 = ~ ( n6297 ) ;
assign n10982 =  ( n10980 ) | ( n10981 )  ;
assign n10983 =  ( n10982 ) | ( n6314 )  ;
assign n10984 = ~ ( n6473 ) ;
assign n10985 =  ( n10983 ) | ( n10984 )  ;
assign n10986 =  ( n10985 ) | ( n6815 )  ;
assign n10987 = ~ ( n7117 ) ;
assign n10988 =  ( n10986 ) | ( n10987 )  ;
assign n10989 =  ( n10988 ) | ( n7445 )  ;
assign n10990 = ~ ( n7765 ) ;
assign n10991 =  ( n10989 ) | ( n10990 )  ;
assign n10992 =  ( n10991 ) | ( n8121 )  ;
assign n10993 = ~ ( n8413 ) ;
assign n10994 =  ( n10992 ) | ( n10993 )  ;
assign n10995 = ~ ( n8717 ) ;
assign n10996 =  ( n10994 ) | ( n10995 )  ;
assign n10997 = ~ ( n9012 ) ;
assign n10998 =  ( n10996 ) | ( n10997 )  ;
assign n10999 = ~ ( n9252 ) ;
assign n11000 =  ( n10998 ) | ( n10999 )  ;
assign n11001 = ~ ( n9432 ) ;
assign n11002 =  ( n11000 ) | ( n11001 )  ;
assign n11003 = ~ ( n9649 ) ;
assign n11004 =  ( n11002 ) | ( n11003 )  ;
assign n11005 = ~ ( n9713 ) ;
assign n11006 = ~ ( n9751 ) ;
assign n11007 =  ( n11006 ) | ( n9808 )  ;
assign n11008 = ~ ( n9834 ) ;
assign n11009 =  ( n11007 ) | ( n11008 )  ;
assign n11010 = ~ ( n9864 ) ;
assign n11011 =  ( n11009 ) | ( n11010 )  ;
assign n11012 = ~ ( n11011 ) ;
assign n11013 =  ( n11005 ) | ( n11012 )  ;
assign n11014 = ~ ( n9751 ) ;
assign n11015 = ~ ( n9909 ) ;
assign n11016 =  ( n11014 ) | ( n11015 )  ;
assign n11017 = ~ ( n10005 ) ;
assign n11018 = ~ ( n10042 ) ;
assign n11019 = ~ ( n10140 ) ;
assign n11020 =  ( n11018 ) | ( n11019 )  ;
assign n11021 =  ( n11020 ) | ( n10158 )  ;
assign n11022 =  ( n11021 ) | ( n10180 )  ;
assign n11023 = ~ ( n11022 ) ;
assign n11024 =  ( n11017 ) | ( n11023 )  ;
assign n11025 = ~ ( n11024 ) ;
assign n11026 =  ( n11016 ) | ( n11025 )  ;
assign n11027 = ~ ( n11026 ) ;
assign n11028 =  ( n11013 ) | ( n11027 )  ;
assign n11029 = ~ ( n9751 ) ;
assign n11030 = ~ ( n9909 ) ;
assign n11031 =  ( n11029 ) | ( n11030 )  ;
assign n11032 = ~ ( n10042 ) ;
assign n11033 =  ( n11031 ) | ( n11032 )  ;
assign n11034 = ~ ( n10208 ) ;
assign n11035 =  ( n11033 ) | ( n11034 )  ;
assign n11036 = ~ ( n10249 ) ;
assign n11037 = ~ ( n10310 ) ;
assign n11038 =  ( n11036 ) | ( n11037 )  ;
assign n11039 = ~ ( n10358 ) ;
assign n11040 =  ( n10274 ) | ( n11039 )  ;
assign n11041 = ~ ( n10397 ) ;
assign n11042 =  ( n11041 ) | ( n10137 )  ;
assign n11043 =  ( n11042 ) | ( n10412 )  ;
assign n11044 = ~ ( n11043 ) ;
assign n11045 =  ( n11044 ) | ( n10451 )  ;
assign n11046 = ~ ( n11045 ) ;
assign n11047 =  ( n11040 ) | ( n11046 )  ;
assign n11048 = ~ ( n11047 ) ;
assign n11049 =  ( n11038 ) | ( n11048 )  ;
assign n11050 = ~ ( n11049 ) ;
assign n11051 =  ( n11035 ) | ( n11050 )  ;
assign n11052 = ~ ( n11051 ) ;
assign n11053 =  ( n11028 ) | ( n11052 )  ;
assign n11054 = ~ ( n9751 ) ;
assign n11055 = ~ ( n9909 ) ;
assign n11056 =  ( n11054 ) | ( n11055 )  ;
assign n11057 = ~ ( n10042 ) ;
assign n11058 =  ( n11056 ) | ( n11057 )  ;
assign n11059 = ~ ( n10208 ) ;
assign n11060 =  ( n11058 ) | ( n11059 )  ;
assign n11061 =  ( n11060 ) | ( n10274 )  ;
assign n11062 = ~ ( n10358 ) ;
assign n11063 =  ( n11061 ) | ( n11062 )  ;
assign n11064 = ~ ( n10430 ) ;
assign n11065 =  ( n11063 ) | ( n11064 )  ;
assign n11066 =  ( n11065 ) | ( n10467 )  ;
assign n11067 = ~ ( n10480 ) ;
assign n11068 = ~ ( n10533 ) ;
assign n11069 =  ( n10489 ) | ( n11068 )  ;
assign n11070 =  ( n11069 ) | ( n7784 )  ;
assign n11071 = ~ ( n11070 ) ;
assign n11072 =  ( n11067 ) | ( n11071 )  ;
assign n11073 =  ( n10489 ) | ( n10550 )  ;
assign n11074 =  ( n7455 ) ^ ( n10522 )  ;
assign n11075 =  ( n11074 ) ^ ( n10519 )  ;
assign n11076 = ~ ( n11075 ) ;
assign n11077 =  ( n11073 ) | ( n11076 )  ;
assign n11078 = ~ ( n7455 ) ;
assign n11079 =  ( n11077 ) | ( n11078 )  ;
assign n11080 = ~ ( n10564 ) ;
assign n11081 =  ( n11079 ) | ( n11080 )  ;
assign n11082 = kd[1:1] ;
assign n11083 = ~ ( n11082 ) ;
assign n11084 =  ( n11081 ) | ( n11083 )  ;
assign n11085 = ~ ( n11084 ) ;
assign n11086 =  ( n11072 ) | ( n11085 )  ;
assign n11087 = ~ ( n11086 ) ;
assign n11088 =  ( n11066 ) | ( n11087 )  ;
assign n11089 = ~ ( n11088 ) ;
assign n11090 =  ( n11053 ) | ( n11089 )  ;
assign n11091 = ~ ( n11090 ) ;
assign n11092 =  ( n11004 ) | ( n11091 )  ;
assign n11093 = ~ ( n11092 ) ;
assign n11094 =  ( n10978 ) | ( n11093 )  ;
assign n11095 = ~ ( n11094 ) ;
assign n11096 =  ( n5792 ) | ( n11095 )  ;
assign n11097 = ~ ( n11096 ) ;
assign n11098 =  ( n10854 ) ^ ( n11097 )  ;
assign n11099 = ~ ( n11098 ) ;
assign n11100 =  ( n10850 ) | ( n11099 )  ;
assign n11101 = ~ ( n11100 ) ;
assign n11102 =  ( n373 ) | ( n382 )  ;
assign n11103 =  ( n11102 ) ? ( bv_1_0_n2 ) : ( n502 ) ;
assign n11104 = ~ ( n11103 ) ;
assign n11105 =  ( n509 ) ^ ( n11104 )  ;
assign n11106 =  ( n11105 ) ^ ( n10848 )  ;
assign n11107 =  ( n11106 ) ^ ( n5774 )  ;
assign n11108 =  ( n5713 ) | ( n5722 )  ;
assign n11109 =  ( n11108 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11110 = ~ ( n11109 ) ;
assign n11111 =  ( n11107 ) ^ ( n11110 )  ;
assign n11112 = ~ ( n11094 ) ;
assign n11113 =  ( n5792 ) | ( n11112 )  ;
assign n11114 = ~ ( n11113 ) ;
assign n11115 =  ( n11111 ) ^ ( n11114 )  ;
assign n11116 = ~ ( n11115 ) ;
assign n11117 =  ( bv_1_1_n5 ) ^ ( n488 )  ;
assign n11118 =  ( n11117 ) ^ ( n504 )  ;
assign n11119 =  ( n11118 ) ^ ( n10845 )  ;
assign n11120 = ~ ( n11119 ) ;
assign n11121 =  ( n11116 ) | ( n11120 )  ;
assign n11122 = ~ ( n5747 ) ;
assign n11123 = ~ ( n5759 ) ;
assign n11124 =  ( n11122 ) | ( n11123 )  ;
assign n11125 =  ( bv_1_1_n5 ) ^ ( n11124 )  ;
assign n11126 =  ( n5713 ) | ( n5722 )  ;
assign n11127 =  ( n11126 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11128 =  ( n11125 ) ^ ( n11127 )  ;
assign n11129 =  ( n11128 ) ^ ( n11094 )  ;
assign n11130 = ~ ( n11129 ) ;
assign n11131 =  ( n11121 ) | ( n11130 )  ;
assign n11132 = ~ ( n11131 ) ;
assign n11133 =  ( n11101 ) | ( n11132 )  ;
assign n11134 = ~ ( n11115 ) ;
assign n11135 =  ( n488 ) ^ ( n504 )  ;
assign n11136 =  ( n11135 ) ^ ( n10845 )  ;
assign n11137 = ~ ( n5747 ) ;
assign n11138 = ~ ( n5759 ) ;
assign n11139 =  ( n11137 ) | ( n11138 )  ;
assign n11140 =  ( n11136 ) ^ ( n11139 )  ;
assign n11141 =  ( n5713 ) | ( n5722 )  ;
assign n11142 =  ( n11141 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11143 =  ( n11140 ) ^ ( n11142 )  ;
assign n11144 =  ( n11143 ) ^ ( n11094 )  ;
assign n11145 = ~ ( n11144 ) ;
assign n11146 =  ( n11134 ) | ( n11145 )  ;
assign n11147 =  ( n834 ) ^ ( n459 )  ;
assign n11148 =  ( n30 ) | ( n39 )  ;
assign n11149 =  ( n11148 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n11150 = ~ ( n11149 ) ;
assign n11151 =  ( n11147 ) ^ ( n11150 )  ;
assign n11152 =  ( n11151 ) ^ ( n484 )  ;
assign n11153 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n11154 =  ( n11153 ) ^ ( n823 )  ;
assign n11155 =  ( n11154 ) ^ ( n344 )  ;
assign n11156 =  ( n11155 ) ^ ( n454 )  ;
assign n11157 = ~ ( n11156 ) ;
assign n11158 = ~ ( n1212 ) ;
assign n11159 = ~ ( n1224 ) ;
assign n11160 =  ( n11158 ) | ( n11159 )  ;
assign n11161 = ~ ( n11160 ) ;
assign n11162 =  ( n11161 ) | ( n1789 )  ;
assign n11163 = ~ ( n1239 ) ;
assign n11164 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n11165 =  ( n11164 ) ^ ( n1199 )  ;
assign n11166 =  ( n11165 ) ^ ( n666 )  ;
assign n11167 =  ( n11166 ) ^ ( n682 )  ;
assign n11168 =  ( n11167 ) ^ ( n697 )  ;
assign n11169 =  ( n11168 ) ^ ( n759 )  ;
assign n11170 = ~ ( n11169 ) ;
assign n11171 =  ( n11163 ) | ( n11170 )  ;
assign n11172 = ~ ( n1446 ) ;
assign n11173 =  ( n11171 ) | ( n11172 )  ;
assign n11174 =  ( n11173 ) | ( n1828 )  ;
assign n11175 = ~ ( n2070 ) ;
assign n11176 =  ( n11175 ) | ( n2080 )  ;
assign n11177 = ~ ( n2092 ) ;
assign n11178 =  ( n11176 ) | ( n11177 )  ;
assign n11179 = ~ ( n11178 ) ;
assign n11180 = ~ ( n2110 ) ;
assign n11181 = ~ ( n2426 ) ;
assign n11182 =  ( n11180 ) | ( n11181 )  ;
assign n11183 =  ( n11182 ) | ( n2438 )  ;
assign n11184 = ~ ( n11183 ) ;
assign n11185 =  ( n11179 ) | ( n11184 )  ;
assign n11186 = ~ ( n2110 ) ;
assign n11187 =  ( n11186 ) | ( n2453 )  ;
assign n11188 = ~ ( n3062 ) ;
assign n11189 =  ( n11187 ) | ( n11188 )  ;
assign n11190 = ~ ( n11189 ) ;
assign n11191 =  ( n11185 ) | ( n11190 )  ;
assign n11192 = ~ ( n11191 ) ;
assign n11193 =  ( n11174 ) | ( n11192 )  ;
assign n11194 = ~ ( n11193 ) ;
assign n11195 =  ( n11162 ) | ( n11194 )  ;
assign n11196 = ~ ( n1239 ) ;
assign n11197 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n11198 =  ( n11197 ) ^ ( n1199 )  ;
assign n11199 =  ( n11198 ) ^ ( n666 )  ;
assign n11200 =  ( n11199 ) ^ ( n682 )  ;
assign n11201 =  ( n11200 ) ^ ( n697 )  ;
assign n11202 =  ( n11201 ) ^ ( n759 )  ;
assign n11203 = ~ ( n11202 ) ;
assign n11204 =  ( n11196 ) | ( n11203 )  ;
assign n11205 = ~ ( n1446 ) ;
assign n11206 =  ( n11204 ) | ( n11205 )  ;
assign n11207 =  ( n11206 ) | ( n1828 )  ;
assign n11208 = ~ ( n2110 ) ;
assign n11209 =  ( n11207 ) | ( n11208 )  ;
assign n11210 =  ( n11209 ) | ( n2453 )  ;
assign n11211 = ~ ( n2742 ) ;
assign n11212 =  ( n11210 ) | ( n11211 )  ;
assign n11213 =  ( n11212 ) | ( n3085 )  ;
assign n11214 = ~ ( n3366 ) ;
assign n11215 = ~ ( n3392 ) ;
assign n11216 = ~ ( n3623 ) ;
assign n11217 =  ( n11215 ) | ( n11216 )  ;
assign n11218 =  ( n11217 ) | ( n3646 )  ;
assign n11219 = ~ ( n11218 ) ;
assign n11220 =  ( n11214 ) | ( n11219 )  ;
assign n11221 = ~ ( n4184 ) ;
assign n11222 =  ( n11220 ) | ( n11221 )  ;
assign n11223 = ~ ( n3392 ) ;
assign n11224 =  ( n11223 ) | ( n3672 )  ;
assign n11225 =  ( n11224 ) | ( n3985 )  ;
assign n11226 =  ( n11225 ) | ( n4253 )  ;
assign n11227 = ~ ( n4435 ) ;
assign n11228 = ~ ( n4689 ) ;
assign n11229 =  ( n11227 ) | ( n11228 )  ;
assign n11230 =  ( n4458 ) | ( n4710 )  ;
assign n11231 = ~ ( n4916 ) ;
assign n11232 =  ( n11230 ) | ( n11231 )  ;
assign n11233 = ~ ( n11232 ) ;
assign n11234 =  ( n11229 ) | ( n11233 )  ;
assign n11235 = ~ ( n11234 ) ;
assign n11236 =  ( n11226 ) | ( n11235 )  ;
assign n11237 = ~ ( n11236 ) ;
assign n11238 =  ( n11222 ) | ( n11237 )  ;
assign n11239 = ~ ( n11238 ) ;
assign n11240 =  ( n11213 ) | ( n11239 )  ;
assign n11241 = ~ ( n11240 ) ;
assign n11242 =  ( n11195 ) | ( n11241 )  ;
assign n11243 = ~ ( n1239 ) ;
assign n11244 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n11245 =  ( n11244 ) ^ ( n1199 )  ;
assign n11246 =  ( n11245 ) ^ ( n666 )  ;
assign n11247 =  ( n11246 ) ^ ( n682 )  ;
assign n11248 =  ( n11247 ) ^ ( n697 )  ;
assign n11249 =  ( n11248 ) ^ ( n759 )  ;
assign n11250 = ~ ( n11249 ) ;
assign n11251 =  ( n11243 ) | ( n11250 )  ;
assign n11252 = ~ ( n1446 ) ;
assign n11253 =  ( n11251 ) | ( n11252 )  ;
assign n11254 =  ( n11253 ) | ( n1828 )  ;
assign n11255 = ~ ( n2110 ) ;
assign n11256 =  ( n11254 ) | ( n11255 )  ;
assign n11257 =  ( n11256 ) | ( n2453 )  ;
assign n11258 = ~ ( n2742 ) ;
assign n11259 =  ( n11257 ) | ( n11258 )  ;
assign n11260 =  ( n11259 ) | ( n3085 )  ;
assign n11261 = ~ ( n3392 ) ;
assign n11262 =  ( n11260 ) | ( n11261 )  ;
assign n11263 =  ( n11262 ) | ( n3672 )  ;
assign n11264 =  ( n11263 ) | ( n3985 )  ;
assign n11265 =  ( n11264 ) | ( n4253 )  ;
assign n11266 =  ( n11265 ) | ( n4458 )  ;
assign n11267 =  ( n11266 ) | ( n4710 )  ;
assign n11268 = ~ ( n4763 ) ;
assign n11269 =  ( n11267 ) | ( n11268 )  ;
assign n11270 = ~ ( n4938 ) ;
assign n11271 =  ( n11269 ) | ( n11270 )  ;
assign n11272 =  ( n5041 ) | ( n5203 )  ;
assign n11273 =  ( n11272 ) | ( n5345 )  ;
assign n11274 =  ( n5063 ) | ( n5224 )  ;
assign n11275 =  ( n11274 ) | ( n5265 )  ;
assign n11276 =  ( n5366 ) ^ ( n5161 )  ;
assign n11277 =  ( n11276 ) ^ ( n5171 )  ;
assign n11278 =  ( n11277 ) ^ ( n4960 )  ;
assign n11279 =  ( n11278 ) ^ ( n4976 )  ;
assign n11280 =  ( n11279 ) ^ ( n4996 )  ;
assign n11281 =  ( n11280 ) ^ ( n5236 )  ;
assign n11282 = ~ ( n11281 ) ;
assign n11283 =  ( n11275 ) | ( n11282 )  ;
assign n11284 =  ( n5446 ) | ( n5473 )  ;
assign n11285 =  ( n11284 ) | ( n5604 )  ;
assign n11286 = ~ ( n11285 ) ;
assign n11287 =  ( n11283 ) | ( n11286 )  ;
assign n11288 = ~ ( n11287 ) ;
assign n11289 =  ( n11273 ) | ( n11288 )  ;
assign n11290 =  ( n5063 ) | ( n5224 )  ;
assign n11291 =  ( n11290 ) | ( n5265 )  ;
assign n11292 =  ( n5366 ) ^ ( n5161 )  ;
assign n11293 =  ( n11292 ) ^ ( n5171 )  ;
assign n11294 =  ( n11293 ) ^ ( n4960 )  ;
assign n11295 =  ( n11294 ) ^ ( n4976 )  ;
assign n11296 =  ( n11295 ) ^ ( n4996 )  ;
assign n11297 =  ( n11296 ) ^ ( n5236 )  ;
assign n11298 = ~ ( n11297 ) ;
assign n11299 =  ( n11291 ) | ( n11298 )  ;
assign n11300 =  ( n5452 ) ^ ( n5325 )  ;
assign n11301 =  ( n11300 ) ^ ( n5083 )  ;
assign n11302 =  ( n11301 ) ^ ( n5099 )  ;
assign n11303 =  ( n11302 ) ^ ( n5116 )  ;
assign n11304 =  ( n11303 ) ^ ( n5141 )  ;
assign n11305 =  ( n11304 ) ^ ( n5129 )  ;
assign n11306 = ~ ( n11305 ) ;
assign n11307 =  ( n11299 ) | ( n11306 )  ;
assign n11308 =  ( n5489 ) ^ ( n5433 )  ;
assign n11309 =  ( n11308 ) ^ ( n5285 )  ;
assign n11310 =  ( n11309 ) ^ ( n5301 )  ;
assign n11311 =  ( n11310 ) ^ ( n5321 )  ;
assign n11312 = ~ ( n11311 ) ;
assign n11313 =  ( n11307 ) | ( n11312 )  ;
assign n11314 = ~ ( n5547 ) ;
assign n11315 =  ( n11313 ) | ( n11314 )  ;
assign n11316 =  ( n5594 ) ^ ( n5515 )  ;
assign n11317 =  ( n11316 ) ^ ( n5531 )  ;
assign n11318 = ~ ( n11317 ) ;
assign n11319 =  ( n11315 ) | ( n11318 )  ;
assign n11320 =  ( n5568 ) ^ ( n5583 )  ;
assign n11321 =  ( n11320 ) ^ ( n5580 )  ;
assign n11322 = ~ ( n11321 ) ;
assign n11323 =  ( n11319 ) | ( n11322 )  ;
assign n11324 = ~ ( n5648 ) ;
assign n11325 =  ( n11323 ) | ( n11324 )  ;
assign n11326 = ~ ( n5657 ) ;
assign n11327 =  ( n11325 ) | ( n11326 )  ;
assign n11328 = ki[1:1] ;
assign n11329 = ~ ( n11328 ) ;
assign n11330 =  ( n11327 ) | ( n11329 )  ;
assign n11331 = ~ ( n11330 ) ;
assign n11332 =  ( n11289 ) | ( n11331 )  ;
assign n11333 = ~ ( n11332 ) ;
assign n11334 =  ( n11271 ) | ( n11333 )  ;
assign n11335 = ~ ( n11334 ) ;
assign n11336 =  ( n11242 ) | ( n11335 )  ;
assign n11337 = ~ ( n11336 ) ;
assign n11338 =  ( n11157 ) | ( n11337 )  ;
assign n11339 = ~ ( n11338 ) ;
assign n11340 =  ( n11152 ) ^ ( n11339 )  ;
assign n11341 = ~ ( n11340 ) ;
assign n11342 = ~ ( n5959 ) ;
assign n11343 =  ( n5965 ) | ( n5972 )  ;
assign n11344 = ~ ( n11343 ) ;
assign n11345 =  ( n11342 ) | ( n11344 )  ;
assign n11346 = ~ ( n5736 ) ;
assign n11347 =  ( n11346 ) | ( n5742 )  ;
assign n11348 =  ( n11345 ) ^ ( n11347 )  ;
assign n11349 =  ( n5682 ) | ( n5691 )  ;
assign n11350 =  ( n11349 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n11351 = ~ ( n11350 ) ;
assign n11352 =  ( n11348 ) ^ ( n11351 )  ;
assign n11353 =  ( n5713 ) | ( n5722 )  ;
assign n11354 =  ( n11353 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11355 =  ( n11352 ) ^ ( n11354 )  ;
assign n11356 = ~ ( n6264 ) ;
assign n11357 = ~ ( n6279 ) ;
assign n11358 =  ( n11356 ) | ( n11357 )  ;
assign n11359 = ~ ( n11358 ) ;
assign n11360 = ~ ( n6297 ) ;
assign n11361 =  ( n11360 ) | ( n6314 )  ;
assign n11362 = ~ ( n6777 ) ;
assign n11363 =  ( n11361 ) | ( n11362 )  ;
assign n11364 = ~ ( n11363 ) ;
assign n11365 =  ( n11359 ) | ( n11364 )  ;
assign n11366 = ~ ( n6297 ) ;
assign n11367 =  ( n11366 ) | ( n6314 )  ;
assign n11368 = ~ ( n6473 ) ;
assign n11369 =  ( n11367 ) | ( n11368 )  ;
assign n11370 =  ( n11369 ) | ( n6815 )  ;
assign n11371 = ~ ( n7022 ) ;
assign n11372 =  ( n11371 ) | ( n7045 )  ;
assign n11373 = ~ ( n7078 ) ;
assign n11374 =  ( n11372 ) | ( n11373 )  ;
assign n11375 = ~ ( n11374 ) ;
assign n11376 = ~ ( n7117 ) ;
assign n11377 = ~ ( n7392 ) ;
assign n11378 =  ( n11376 ) | ( n11377 )  ;
assign n11379 =  ( n11378 ) | ( n7417 )  ;
assign n11380 = ~ ( n11379 ) ;
assign n11381 =  ( n11375 ) | ( n11380 )  ;
assign n11382 = ~ ( n7117 ) ;
assign n11383 =  ( n11382 ) | ( n7445 )  ;
assign n11384 = ~ ( n8082 ) ;
assign n11385 =  ( n11383 ) | ( n11384 )  ;
assign n11386 = ~ ( n11385 ) ;
assign n11387 =  ( n11381 ) | ( n11386 )  ;
assign n11388 = ~ ( n11387 ) ;
assign n11389 =  ( n11370 ) | ( n11388 )  ;
assign n11390 = ~ ( n11389 ) ;
assign n11391 =  ( n11365 ) | ( n11390 )  ;
assign n11392 = ~ ( n6297 ) ;
assign n11393 =  ( n11392 ) | ( n6314 )  ;
assign n11394 = ~ ( n6473 ) ;
assign n11395 =  ( n11393 ) | ( n11394 )  ;
assign n11396 =  ( n11395 ) | ( n6815 )  ;
assign n11397 = ~ ( n7117 ) ;
assign n11398 =  ( n11396 ) | ( n11397 )  ;
assign n11399 =  ( n11398 ) | ( n7445 )  ;
assign n11400 = ~ ( n7765 ) ;
assign n11401 =  ( n11399 ) | ( n11400 )  ;
assign n11402 =  ( n11401 ) | ( n8121 )  ;
assign n11403 = ~ ( n8279 ) ;
assign n11404 = ~ ( n8321 ) ;
assign n11405 =  ( n11403 ) | ( n11404 )  ;
assign n11406 = ~ ( n8364 ) ;
assign n11407 =  ( n11405 ) | ( n11406 )  ;
assign n11408 = ~ ( n11407 ) ;
assign n11409 = ~ ( n8413 ) ;
assign n11410 = ~ ( n8625 ) ;
assign n11411 =  ( n11409 ) | ( n11410 )  ;
assign n11412 = ~ ( n8669 ) ;
assign n11413 =  ( n11411 ) | ( n11412 )  ;
assign n11414 = ~ ( n11413 ) ;
assign n11415 =  ( n11408 ) | ( n11414 )  ;
assign n11416 = ~ ( n8413 ) ;
assign n11417 = ~ ( n8717 ) ;
assign n11418 =  ( n11416 ) | ( n11417 )  ;
assign n11419 = ~ ( n9172 ) ;
assign n11420 =  ( n11418 ) | ( n11419 )  ;
assign n11421 = ~ ( n11420 ) ;
assign n11422 =  ( n11415 ) | ( n11421 )  ;
assign n11423 = ~ ( n8413 ) ;
assign n11424 = ~ ( n8717 ) ;
assign n11425 =  ( n11423 ) | ( n11424 )  ;
assign n11426 = ~ ( n9012 ) ;
assign n11427 =  ( n11425 ) | ( n11426 )  ;
assign n11428 = ~ ( n9252 ) ;
assign n11429 =  ( n11427 ) | ( n11428 )  ;
assign n11430 = ~ ( n9314 ) ;
assign n11431 = ~ ( n9348 ) ;
assign n11432 =  ( n11430 ) | ( n11431 )  ;
assign n11433 = ~ ( n9387 ) ;
assign n11434 =  ( n11432 ) | ( n11433 )  ;
assign n11435 = ~ ( n11434 ) ;
assign n11436 =  ( n11435 ) | ( n9608 )  ;
assign n11437 = ~ ( n9432 ) ;
assign n11438 = ~ ( n9649 ) ;
assign n11439 =  ( n11437 ) | ( n11438 )  ;
assign n11440 = ~ ( n9868 ) ;
assign n11441 =  ( n11439 ) | ( n11440 )  ;
assign n11442 = ~ ( n11441 ) ;
assign n11443 =  ( n11436 ) | ( n11442 )  ;
assign n11444 = ~ ( n11443 ) ;
assign n11445 =  ( n11429 ) | ( n11444 )  ;
assign n11446 = ~ ( n11445 ) ;
assign n11447 =  ( n11422 ) | ( n11446 )  ;
assign n11448 = ~ ( n11447 ) ;
assign n11449 =  ( n11402 ) | ( n11448 )  ;
assign n11450 = ~ ( n11449 ) ;
assign n11451 =  ( n11391 ) | ( n11450 )  ;
assign n11452 = ~ ( n6297 ) ;
assign n11453 =  ( n11452 ) | ( n6314 )  ;
assign n11454 = ~ ( n6473 ) ;
assign n11455 =  ( n11453 ) | ( n11454 )  ;
assign n11456 =  ( n11455 ) | ( n6815 )  ;
assign n11457 = ~ ( n7117 ) ;
assign n11458 =  ( n11456 ) | ( n11457 )  ;
assign n11459 =  ( n11458 ) | ( n7445 )  ;
assign n11460 = ~ ( n7765 ) ;
assign n11461 =  ( n11459 ) | ( n11460 )  ;
assign n11462 =  ( n11461 ) | ( n8121 )  ;
assign n11463 = ~ ( n8413 ) ;
assign n11464 =  ( n11462 ) | ( n11463 )  ;
assign n11465 = ~ ( n8717 ) ;
assign n11466 =  ( n11464 ) | ( n11465 )  ;
assign n11467 = ~ ( n9012 ) ;
assign n11468 =  ( n11466 ) | ( n11467 )  ;
assign n11469 = ~ ( n9252 ) ;
assign n11470 =  ( n11468 ) | ( n11469 )  ;
assign n11471 = ~ ( n9432 ) ;
assign n11472 =  ( n11470 ) | ( n11471 )  ;
assign n11473 = ~ ( n9649 ) ;
assign n11474 =  ( n11472 ) | ( n11473 )  ;
assign n11475 = ~ ( n9751 ) ;
assign n11476 =  ( n11474 ) | ( n11475 )  ;
assign n11477 = ~ ( n9909 ) ;
assign n11478 =  ( n11476 ) | ( n11477 )  ;
assign n11479 = ~ ( n10005 ) ;
assign n11480 = ~ ( n10042 ) ;
assign n11481 = ~ ( n10140 ) ;
assign n11482 =  ( n11480 ) | ( n11481 )  ;
assign n11483 =  ( n11482 ) | ( n10158 )  ;
assign n11484 =  ( n11483 ) | ( n10180 )  ;
assign n11485 = ~ ( n11484 ) ;
assign n11486 =  ( n11479 ) | ( n11485 )  ;
assign n11487 = ~ ( n10314 ) ;
assign n11488 =  ( n11486 ) | ( n11487 )  ;
assign n11489 = ~ ( n10042 ) ;
assign n11490 = ~ ( n10208 ) ;
assign n11491 =  ( n11489 ) | ( n11490 )  ;
assign n11492 =  ( n11491 ) | ( n10274 )  ;
assign n11493 = ~ ( n10358 ) ;
assign n11494 =  ( n11492 ) | ( n11493 )  ;
assign n11495 = ~ ( n10397 ) ;
assign n11496 =  ( n11495 ) | ( n10137 )  ;
assign n11497 =  ( n11496 ) | ( n10412 )  ;
assign n11498 = ~ ( n11497 ) ;
assign n11499 =  ( n11498 ) | ( n10451 )  ;
assign n11500 = ~ ( n10430 ) ;
assign n11501 =  ( n11500 ) | ( n10467 )  ;
assign n11502 = ~ ( n10538 ) ;
assign n11503 =  ( n11501 ) | ( n11502 )  ;
assign n11504 = ~ ( n11503 ) ;
assign n11505 =  ( n11499 ) | ( n11504 )  ;
assign n11506 = ~ ( n11505 ) ;
assign n11507 =  ( n11494 ) | ( n11506 )  ;
assign n11508 = ~ ( n11507 ) ;
assign n11509 =  ( n11488 ) | ( n11508 )  ;
assign n11510 = ~ ( n10042 ) ;
assign n11511 = ~ ( n10208 ) ;
assign n11512 =  ( n11510 ) | ( n11511 )  ;
assign n11513 =  ( n11512 ) | ( n10274 )  ;
assign n11514 = ~ ( n10358 ) ;
assign n11515 =  ( n11513 ) | ( n11514 )  ;
assign n11516 = ~ ( n10430 ) ;
assign n11517 =  ( n11515 ) | ( n11516 )  ;
assign n11518 =  ( n11517 ) | ( n10467 )  ;
assign n11519 =  ( n11518 ) | ( n10489 )  ;
assign n11520 =  ( n11519 ) | ( n10550 )  ;
assign n11521 =  ( n7455 ) ^ ( n10522 )  ;
assign n11522 =  ( n11521 ) ^ ( n10519 )  ;
assign n11523 = ~ ( n11522 ) ;
assign n11524 =  ( n11520 ) | ( n11523 )  ;
assign n11525 = ~ ( n7455 ) ;
assign n11526 =  ( n11524 ) | ( n11525 )  ;
assign n11527 = ~ ( n10564 ) ;
assign n11528 =  ( n11526 ) | ( n11527 )  ;
assign n11529 = kd[1:1] ;
assign n11530 = ~ ( n11529 ) ;
assign n11531 =  ( n11528 ) | ( n11530 )  ;
assign n11532 = ~ ( n11531 ) ;
assign n11533 =  ( n11509 ) | ( n11532 )  ;
assign n11534 = ~ ( n11533 ) ;
assign n11535 =  ( n11478 ) | ( n11534 )  ;
assign n11536 = ~ ( n11535 ) ;
assign n11537 =  ( n11451 ) | ( n11536 )  ;
assign n11538 = ~ ( n11537 ) ;
assign n11539 =  ( n6020 ) | ( n11538 )  ;
assign n11540 = ~ ( n11539 ) ;
assign n11541 =  ( n11355 ) ^ ( n11540 )  ;
assign n11542 = ~ ( n11541 ) ;
assign n11543 =  ( n11341 ) | ( n11542 )  ;
assign n11544 = ~ ( n11543 ) ;
assign n11545 =  ( n834 ) ^ ( n459 )  ;
assign n11546 =  ( n30 ) | ( n39 )  ;
assign n11547 =  ( n11546 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n11548 = ~ ( n11547 ) ;
assign n11549 =  ( n11545 ) ^ ( n11548 )  ;
assign n11550 =  ( n11549 ) ^ ( n484 )  ;
assign n11551 =  ( n11550 ) ^ ( n11339 )  ;
assign n11552 = ~ ( n5959 ) ;
assign n11553 =  ( n5965 ) | ( n5972 )  ;
assign n11554 = ~ ( n11553 ) ;
assign n11555 =  ( n11552 ) | ( n11554 )  ;
assign n11556 =  ( n11551 ) ^ ( n11555 )  ;
assign n11557 = ~ ( n5736 ) ;
assign n11558 =  ( n11557 ) | ( n5742 )  ;
assign n11559 =  ( n11556 ) ^ ( n11558 )  ;
assign n11560 =  ( n5682 ) | ( n5691 )  ;
assign n11561 =  ( n11560 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n11562 = ~ ( n11561 ) ;
assign n11563 =  ( n11559 ) ^ ( n11562 )  ;
assign n11564 =  ( n5713 ) | ( n5722 )  ;
assign n11565 =  ( n11564 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11566 =  ( n11563 ) ^ ( n11565 )  ;
assign n11567 = ~ ( n11537 ) ;
assign n11568 =  ( n6020 ) | ( n11567 )  ;
assign n11569 = ~ ( n11568 ) ;
assign n11570 =  ( n11566 ) ^ ( n11569 )  ;
assign n11571 = ~ ( n11570 ) ;
assign n11572 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n11573 =  ( n11572 ) ^ ( n823 )  ;
assign n11574 =  ( n11573 ) ^ ( n344 )  ;
assign n11575 =  ( n11574 ) ^ ( n454 )  ;
assign n11576 =  ( n11575 ) ^ ( n11336 )  ;
assign n11577 = ~ ( n11576 ) ;
assign n11578 =  ( n11571 ) | ( n11577 )  ;
assign n11579 =  ( bv_1_1_n5 ) ^ ( n5936 )  ;
assign n11580 = ~ ( n5943 ) ;
assign n11581 = ~ ( n5955 ) ;
assign n11582 =  ( n11580 ) | ( n11581 )  ;
assign n11583 =  ( n11579 ) ^ ( n11582 )  ;
assign n11584 =  ( n5682 ) | ( n5691 )  ;
assign n11585 =  ( n11584 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n11586 =  ( n11583 ) ^ ( n11585 )  ;
assign n11587 =  ( n5713 ) | ( n5722 )  ;
assign n11588 =  ( n11587 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11589 =  ( n11586 ) ^ ( n11588 )  ;
assign n11590 =  ( n11589 ) ^ ( n11537 )  ;
assign n11591 = ~ ( n11590 ) ;
assign n11592 =  ( n11578 ) | ( n11591 )  ;
assign n11593 = ~ ( n11592 ) ;
assign n11594 =  ( n11544 ) | ( n11593 )  ;
assign n11595 = ~ ( n11594 ) ;
assign n11596 =  ( n11146 ) | ( n11595 )  ;
assign n11597 = ~ ( n11596 ) ;
assign n11598 =  ( n11133 ) | ( n11597 )  ;
assign n11599 = ~ ( n11115 ) ;
assign n11600 =  ( n11599 ) | ( n11145 )  ;
assign n11601 = ~ ( n11570 ) ;
assign n11602 =  ( n11600 ) | ( n11601 )  ;
assign n11603 =  ( n808 ) ^ ( n823 )  ;
assign n11604 =  ( n11603 ) ^ ( n344 )  ;
assign n11605 =  ( n11604 ) ^ ( n454 )  ;
assign n11606 =  ( n11605 ) ^ ( n11336 )  ;
assign n11607 =  ( n11606 ) ^ ( n5936 )  ;
assign n11608 = ~ ( n5943 ) ;
assign n11609 = ~ ( n5955 ) ;
assign n11610 =  ( n11608 ) | ( n11609 )  ;
assign n11611 =  ( n11607 ) ^ ( n11610 )  ;
assign n11612 =  ( n5682 ) | ( n5691 )  ;
assign n11613 =  ( n11612 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n11614 =  ( n11611 ) ^ ( n11613 )  ;
assign n11615 =  ( n5713 ) | ( n5722 )  ;
assign n11616 =  ( n11615 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11617 =  ( n11614 ) ^ ( n11616 )  ;
assign n11618 =  ( n11617 ) ^ ( n11537 )  ;
assign n11619 = ~ ( n11618 ) ;
assign n11620 =  ( n11602 ) | ( n11619 )  ;
assign n11621 =  ( n666 ) ^ ( n682 )  ;
assign n11622 =  ( n11621 ) ^ ( n697 )  ;
assign n11623 =  ( n11622 ) ^ ( n759 )  ;
assign n11624 =  ( n763 ) | ( n11623 )  ;
assign n11625 =  ( n1212 ) ^ ( n11624 )  ;
assign n11626 =  ( n11625 ) ^ ( n778 )  ;
assign n11627 =  ( n586 ) | ( n595 )  ;
assign n11628 =  ( n11627 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n11629 = ~ ( n11628 ) ;
assign n11630 =  ( n11626 ) ^ ( n11629 )  ;
assign n11631 =  ( n11630 ) ^ ( n796 )  ;
assign n11632 =  ( n11631 ) ^ ( n803 )  ;
assign n11633 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n11634 =  ( n11633 ) ^ ( n1199 )  ;
assign n11635 =  ( n11634 ) ^ ( n666 )  ;
assign n11636 =  ( n11635 ) ^ ( n682 )  ;
assign n11637 =  ( n11636 ) ^ ( n697 )  ;
assign n11638 =  ( n11637 ) ^ ( n759 )  ;
assign n11639 = ~ ( n11638 ) ;
assign n11640 = ~ ( n1446 ) ;
assign n11641 = ~ ( n1773 ) ;
assign n11642 =  ( n11640 ) | ( n11641 )  ;
assign n11643 =  ( n11642 ) | ( n1783 )  ;
assign n11644 = ~ ( n11643 ) ;
assign n11645 =  ( n1426 ) | ( n11644 )  ;
assign n11646 = ~ ( n1446 ) ;
assign n11647 =  ( n11646 ) | ( n1828 )  ;
assign n11648 = ~ ( n10641 ) ;
assign n11649 =  ( n11647 ) | ( n11648 )  ;
assign n11650 = ~ ( n11649 ) ;
assign n11651 =  ( n11645 ) | ( n11650 )  ;
assign n11652 = ~ ( n1446 ) ;
assign n11653 =  ( n11652 ) | ( n1828 )  ;
assign n11654 = ~ ( n2110 ) ;
assign n11655 =  ( n11653 ) | ( n11654 )  ;
assign n11656 =  ( n11655 ) | ( n2453 )  ;
assign n11657 = ~ ( n2722 ) ;
assign n11658 = ~ ( n2742 ) ;
assign n11659 = ~ ( n3043 ) ;
assign n11660 =  ( n11658 ) | ( n11659 )  ;
assign n11661 =  ( n11660 ) | ( n3059 )  ;
assign n11662 = ~ ( n11661 ) ;
assign n11663 =  ( n11657 ) | ( n11662 )  ;
assign n11664 = ~ ( n2742 ) ;
assign n11665 =  ( n11664 ) | ( n3085 )  ;
assign n11666 = ~ ( n10688 ) ;
assign n11667 =  ( n11665 ) | ( n11666 )  ;
assign n11668 = ~ ( n11667 ) ;
assign n11669 =  ( n11663 ) | ( n11668 )  ;
assign n11670 = ~ ( n11669 ) ;
assign n11671 =  ( n11656 ) | ( n11670 )  ;
assign n11672 = ~ ( n11671 ) ;
assign n11673 =  ( n11651 ) | ( n11672 )  ;
assign n11674 = ~ ( n1446 ) ;
assign n11675 =  ( n11674 ) | ( n1828 )  ;
assign n11676 = ~ ( n2110 ) ;
assign n11677 =  ( n11675 ) | ( n11676 )  ;
assign n11678 =  ( n11677 ) | ( n2453 )  ;
assign n11679 = ~ ( n2742 ) ;
assign n11680 =  ( n11678 ) | ( n11679 )  ;
assign n11681 =  ( n11680 ) | ( n3085 )  ;
assign n11682 = ~ ( n3392 ) ;
assign n11683 =  ( n11681 ) | ( n11682 )  ;
assign n11684 =  ( n11683 ) | ( n3672 )  ;
assign n11685 = ~ ( n3958 ) ;
assign n11686 =  ( n11685 ) | ( n4181 )  ;
assign n11687 = ~ ( n10705 ) ;
assign n11688 =  ( n11686 ) | ( n11687 )  ;
assign n11689 =  ( n3985 ) | ( n4253 )  ;
assign n11690 =  ( n11689 ) | ( n4458 )  ;
assign n11691 =  ( n11690 ) | ( n4710 )  ;
assign n11692 = ~ ( n4728 ) ;
assign n11693 =  ( n4722 ) | ( n11692 )  ;
assign n11694 =  ( n11693 ) | ( n4744 )  ;
assign n11695 = ~ ( n11694 ) ;
assign n11696 = ~ ( n4763 ) ;
assign n11697 = ~ ( n4889 ) ;
assign n11698 =  ( n11696 ) | ( n11697 )  ;
assign n11699 =  ( n11698 ) | ( n4900 )  ;
assign n11700 =  ( n11699 ) | ( n4913 )  ;
assign n11701 = ~ ( n11700 ) ;
assign n11702 =  ( n11695 ) | ( n11701 )  ;
assign n11703 =  ( n11702 ) | ( n10766 )  ;
assign n11704 = ~ ( n11703 ) ;
assign n11705 =  ( n11691 ) | ( n11704 )  ;
assign n11706 = ~ ( n11705 ) ;
assign n11707 =  ( n11688 ) | ( n11706 )  ;
assign n11708 = ~ ( n11707 ) ;
assign n11709 =  ( n11684 ) | ( n11708 )  ;
assign n11710 = ~ ( n11709 ) ;
assign n11711 =  ( n11673 ) | ( n11710 )  ;
assign n11712 = ~ ( n1446 ) ;
assign n11713 =  ( n11712 ) | ( n1828 )  ;
assign n11714 = ~ ( n2110 ) ;
assign n11715 =  ( n11713 ) | ( n11714 )  ;
assign n11716 =  ( n11715 ) | ( n2453 )  ;
assign n11717 = ~ ( n2742 ) ;
assign n11718 =  ( n11716 ) | ( n11717 )  ;
assign n11719 =  ( n11718 ) | ( n3085 )  ;
assign n11720 = ~ ( n3392 ) ;
assign n11721 =  ( n11719 ) | ( n11720 )  ;
assign n11722 =  ( n11721 ) | ( n3672 )  ;
assign n11723 =  ( n11722 ) | ( n3985 )  ;
assign n11724 =  ( n11723 ) | ( n4253 )  ;
assign n11725 =  ( n11724 ) | ( n4458 )  ;
assign n11726 =  ( n11725 ) | ( n4710 )  ;
assign n11727 = ~ ( n4763 ) ;
assign n11728 =  ( n11726 ) | ( n11727 )  ;
assign n11729 = ~ ( n4938 ) ;
assign n11730 =  ( n11728 ) | ( n11729 )  ;
assign n11731 =  ( n11730 ) | ( n5063 )  ;
assign n11732 =  ( n11731 ) | ( n5224 )  ;
assign n11733 =  ( n5248 ) | ( n5341 )  ;
assign n11734 =  ( n11733 ) | ( n10785 )  ;
assign n11735 =  ( n5366 ) ^ ( n5161 )  ;
assign n11736 =  ( n11735 ) ^ ( n5171 )  ;
assign n11737 =  ( n11736 ) ^ ( n4960 )  ;
assign n11738 =  ( n11737 ) ^ ( n4976 )  ;
assign n11739 =  ( n11738 ) ^ ( n4996 )  ;
assign n11740 =  ( n11739 ) ^ ( n5236 )  ;
assign n11741 = ~ ( n11740 ) ;
assign n11742 =  ( n5265 ) | ( n11741 )  ;
assign n11743 =  ( n5452 ) ^ ( n5325 )  ;
assign n11744 =  ( n11743 ) ^ ( n5083 )  ;
assign n11745 =  ( n11744 ) ^ ( n5099 )  ;
assign n11746 =  ( n11745 ) ^ ( n5116 )  ;
assign n11747 =  ( n11746 ) ^ ( n5141 )  ;
assign n11748 =  ( n11747 ) ^ ( n5129 )  ;
assign n11749 = ~ ( n11748 ) ;
assign n11750 =  ( n11742 ) | ( n11749 )  ;
assign n11751 =  ( n5489 ) ^ ( n5433 )  ;
assign n11752 =  ( n11751 ) ^ ( n5285 )  ;
assign n11753 =  ( n11752 ) ^ ( n5301 )  ;
assign n11754 =  ( n11753 ) ^ ( n5321 )  ;
assign n11755 = ~ ( n11754 ) ;
assign n11756 =  ( n11750 ) | ( n11755 )  ;
assign n11757 =  ( n5539 ) | ( n5600 )  ;
assign n11758 = ~ ( n11757 ) ;
assign n11759 =  ( n11756 ) | ( n11758 )  ;
assign n11760 = ~ ( n11759 ) ;
assign n11761 =  ( n11734 ) | ( n11760 )  ;
assign n11762 =  ( n5366 ) ^ ( n5161 )  ;
assign n11763 =  ( n11762 ) ^ ( n5171 )  ;
assign n11764 =  ( n11763 ) ^ ( n4960 )  ;
assign n11765 =  ( n11764 ) ^ ( n4976 )  ;
assign n11766 =  ( n11765 ) ^ ( n4996 )  ;
assign n11767 =  ( n11766 ) ^ ( n5236 )  ;
assign n11768 = ~ ( n11767 ) ;
assign n11769 =  ( n5265 ) | ( n11768 )  ;
assign n11770 =  ( n5452 ) ^ ( n5325 )  ;
assign n11771 =  ( n11770 ) ^ ( n5083 )  ;
assign n11772 =  ( n11771 ) ^ ( n5099 )  ;
assign n11773 =  ( n11772 ) ^ ( n5116 )  ;
assign n11774 =  ( n11773 ) ^ ( n5141 )  ;
assign n11775 =  ( n11774 ) ^ ( n5129 )  ;
assign n11776 = ~ ( n11775 ) ;
assign n11777 =  ( n11769 ) | ( n11776 )  ;
assign n11778 =  ( n5489 ) ^ ( n5433 )  ;
assign n11779 =  ( n11778 ) ^ ( n5285 )  ;
assign n11780 =  ( n11779 ) ^ ( n5301 )  ;
assign n11781 =  ( n11780 ) ^ ( n5321 )  ;
assign n11782 = ~ ( n11781 ) ;
assign n11783 =  ( n11777 ) | ( n11782 )  ;
assign n11784 = ~ ( n5547 ) ;
assign n11785 =  ( n11783 ) | ( n11784 )  ;
assign n11786 =  ( n5594 ) ^ ( n5515 )  ;
assign n11787 =  ( n11786 ) ^ ( n5531 )  ;
assign n11788 = ~ ( n11787 ) ;
assign n11789 =  ( n11785 ) | ( n11788 )  ;
assign n11790 =  ( n5568 ) ^ ( n5583 )  ;
assign n11791 =  ( n11790 ) ^ ( n5580 )  ;
assign n11792 = ~ ( n11791 ) ;
assign n11793 =  ( n11789 ) | ( n11792 )  ;
assign n11794 = ~ ( n5648 ) ;
assign n11795 =  ( n11793 ) | ( n11794 )  ;
assign n11796 = ~ ( n5657 ) ;
assign n11797 =  ( n11795 ) | ( n11796 )  ;
assign n11798 = ki[1:1] ;
assign n11799 = ~ ( n11798 ) ;
assign n11800 =  ( n11797 ) | ( n11799 )  ;
assign n11801 = ~ ( n11800 ) ;
assign n11802 =  ( n11761 ) | ( n11801 )  ;
assign n11803 = ~ ( n11802 ) ;
assign n11804 =  ( n11732 ) | ( n11803 )  ;
assign n11805 = ~ ( n11804 ) ;
assign n11806 =  ( n11711 ) | ( n11805 )  ;
assign n11807 = ~ ( n11806 ) ;
assign n11808 =  ( n11639 ) | ( n11807 )  ;
assign n11809 = ~ ( n11808 ) ;
assign n11810 =  ( n11632 ) ^ ( n11809 )  ;
assign n11811 = ~ ( n11810 ) ;
assign n11812 =  ( n6264 ) ^ ( n5894 )  ;
assign n11813 = ~ ( n5902 ) ;
assign n11814 = ~ ( n5913 ) ;
assign n11815 =  ( n11813 ) | ( n11814 )  ;
assign n11816 =  ( n11812 ) ^ ( n11815 )  ;
assign n11817 =  ( n5832 ) | ( n5841 )  ;
assign n11818 =  ( n11817 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n11819 = ~ ( n11818 ) ;
assign n11820 =  ( n11816 ) ^ ( n11819 )  ;
assign n11821 =  ( n5682 ) | ( n5691 )  ;
assign n11822 =  ( n11821 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n11823 =  ( n11820 ) ^ ( n11822 )  ;
assign n11824 =  ( n5713 ) | ( n5722 )  ;
assign n11825 =  ( n11824 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n11826 =  ( n11823 ) ^ ( n11825 )  ;
assign n11827 = ~ ( n6402 ) ;
assign n11828 =  ( n11827 ) | ( n6421 )  ;
assign n11829 = ~ ( n6444 ) ;
assign n11830 =  ( n11828 ) | ( n11829 )  ;
assign n11831 = ~ ( n11830 ) ;
assign n11832 = ~ ( n6473 ) ;
assign n11833 = ~ ( n6753 ) ;
assign n11834 =  ( n11832 ) | ( n11833 )  ;
assign n11835 =  ( n11834 ) | ( n6774 )  ;
assign n11836 = ~ ( n11835 ) ;
assign n11837 =  ( n11831 ) | ( n11836 )  ;
assign n11838 = ~ ( n6473 ) ;
assign n11839 =  ( n11838 ) | ( n6815 )  ;
assign n11840 = ~ ( n10894 ) ;
assign n11841 =  ( n11839 ) | ( n11840 )  ;
assign n11842 = ~ ( n11841 ) ;
assign n11843 =  ( n11837 ) | ( n11842 )  ;
assign n11844 = ~ ( n6473 ) ;
assign n11845 =  ( n11844 ) | ( n6815 )  ;
assign n11846 = ~ ( n7117 ) ;
assign n11847 =  ( n11845 ) | ( n11846 )  ;
assign n11848 =  ( n11847 ) | ( n7445 )  ;
assign n11849 = ~ ( n7649 ) ;
assign n11850 =  ( n11849 ) | ( n7679 )  ;
assign n11851 = ~ ( n7719 ) ;
assign n11852 =  ( n11850 ) | ( n11851 )  ;
assign n11853 = ~ ( n11852 ) ;
assign n11854 = ~ ( n7765 ) ;
assign n11855 = ~ ( n8047 ) ;
assign n11856 =  ( n11854 ) | ( n11855 )  ;
assign n11857 =  ( n11856 ) | ( n8079 )  ;
assign n11858 = ~ ( n11857 ) ;
assign n11859 =  ( n11853 ) | ( n11858 )  ;
assign n11860 = ~ ( n7765 ) ;
assign n11861 =  ( n11860 ) | ( n8121 )  ;
assign n11862 = ~ ( n10939 ) ;
assign n11863 =  ( n11861 ) | ( n11862 )  ;
assign n11864 = ~ ( n11863 ) ;
assign n11865 =  ( n11859 ) | ( n11864 )  ;
assign n11866 = ~ ( n11865 ) ;
assign n11867 =  ( n11848 ) | ( n11866 )  ;
assign n11868 = ~ ( n11867 ) ;
assign n11869 =  ( n11843 ) | ( n11868 )  ;
assign n11870 = ~ ( n6473 ) ;
assign n11871 =  ( n11870 ) | ( n6815 )  ;
assign n11872 = ~ ( n7117 ) ;
assign n11873 =  ( n11871 ) | ( n11872 )  ;
assign n11874 =  ( n11873 ) | ( n7445 )  ;
assign n11875 = ~ ( n7765 ) ;
assign n11876 =  ( n11874 ) | ( n11875 )  ;
assign n11877 =  ( n11876 ) | ( n8121 )  ;
assign n11878 = ~ ( n8413 ) ;
assign n11879 =  ( n11877 ) | ( n11878 )  ;
assign n11880 = ~ ( n8717 ) ;
assign n11881 =  ( n11879 ) | ( n11880 )  ;
assign n11882 = ~ ( n8880 ) ;
assign n11883 = ~ ( n8920 ) ;
assign n11884 =  ( n11882 ) | ( n11883 )  ;
assign n11885 = ~ ( n8963 ) ;
assign n11886 =  ( n11884 ) | ( n11885 )  ;
assign n11887 = ~ ( n11886 ) ;
assign n11888 =  ( n11887 ) | ( n9171 )  ;
assign n11889 = ~ ( n9012 ) ;
assign n11890 = ~ ( n9252 ) ;
assign n11891 =  ( n11889 ) | ( n11890 )  ;
assign n11892 = ~ ( n10966 ) ;
assign n11893 =  ( n11891 ) | ( n11892 )  ;
assign n11894 = ~ ( n11893 ) ;
assign n11895 =  ( n11888 ) | ( n11894 )  ;
assign n11896 = ~ ( n9012 ) ;
assign n11897 = ~ ( n9252 ) ;
assign n11898 =  ( n11896 ) | ( n11897 )  ;
assign n11899 = ~ ( n9432 ) ;
assign n11900 =  ( n11898 ) | ( n11899 )  ;
assign n11901 = ~ ( n9649 ) ;
assign n11902 =  ( n11900 ) | ( n11901 )  ;
assign n11903 = ~ ( n9713 ) ;
assign n11904 = ~ ( n9751 ) ;
assign n11905 =  ( n11904 ) | ( n9808 )  ;
assign n11906 = ~ ( n9834 ) ;
assign n11907 =  ( n11905 ) | ( n11906 )  ;
assign n11908 = ~ ( n9864 ) ;
assign n11909 =  ( n11907 ) | ( n11908 )  ;
assign n11910 = ~ ( n11909 ) ;
assign n11911 =  ( n11903 ) | ( n11910 )  ;
assign n11912 = ~ ( n9751 ) ;
assign n11913 = ~ ( n9909 ) ;
assign n11914 =  ( n11912 ) | ( n11913 )  ;
assign n11915 = ~ ( n11024 ) ;
assign n11916 =  ( n11914 ) | ( n11915 )  ;
assign n11917 = ~ ( n11916 ) ;
assign n11918 =  ( n11911 ) | ( n11917 )  ;
assign n11919 = ~ ( n11918 ) ;
assign n11920 =  ( n11902 ) | ( n11919 )  ;
assign n11921 = ~ ( n11920 ) ;
assign n11922 =  ( n11895 ) | ( n11921 )  ;
assign n11923 = ~ ( n11922 ) ;
assign n11924 =  ( n11881 ) | ( n11923 )  ;
assign n11925 = ~ ( n11924 ) ;
assign n11926 =  ( n11869 ) | ( n11925 )  ;
assign n11927 = ~ ( n6473 ) ;
assign n11928 =  ( n11927 ) | ( n6815 )  ;
assign n11929 = ~ ( n7117 ) ;
assign n11930 =  ( n11928 ) | ( n11929 )  ;
assign n11931 =  ( n11930 ) | ( n7445 )  ;
assign n11932 = ~ ( n7765 ) ;
assign n11933 =  ( n11931 ) | ( n11932 )  ;
assign n11934 =  ( n11933 ) | ( n8121 )  ;
assign n11935 = ~ ( n8413 ) ;
assign n11936 =  ( n11934 ) | ( n11935 )  ;
assign n11937 = ~ ( n8717 ) ;
assign n11938 =  ( n11936 ) | ( n11937 )  ;
assign n11939 = ~ ( n9012 ) ;
assign n11940 =  ( n11938 ) | ( n11939 )  ;
assign n11941 = ~ ( n9252 ) ;
assign n11942 =  ( n11940 ) | ( n11941 )  ;
assign n11943 = ~ ( n9432 ) ;
assign n11944 =  ( n11942 ) | ( n11943 )  ;
assign n11945 = ~ ( n9649 ) ;
assign n11946 =  ( n11944 ) | ( n11945 )  ;
assign n11947 = ~ ( n9751 ) ;
assign n11948 =  ( n11946 ) | ( n11947 )  ;
assign n11949 = ~ ( n9909 ) ;
assign n11950 =  ( n11948 ) | ( n11949 )  ;
assign n11951 = ~ ( n10042 ) ;
assign n11952 =  ( n11950 ) | ( n11951 )  ;
assign n11953 = ~ ( n10208 ) ;
assign n11954 =  ( n11952 ) | ( n11953 )  ;
assign n11955 = ~ ( n10249 ) ;
assign n11956 = ~ ( n10310 ) ;
assign n11957 =  ( n11955 ) | ( n11956 )  ;
assign n11958 = ~ ( n10358 ) ;
assign n11959 =  ( n10274 ) | ( n11958 )  ;
assign n11960 = ~ ( n11045 ) ;
assign n11961 =  ( n11959 ) | ( n11960 )  ;
assign n11962 = ~ ( n11961 ) ;
assign n11963 =  ( n11957 ) | ( n11962 )  ;
assign n11964 = ~ ( n10358 ) ;
assign n11965 =  ( n10274 ) | ( n11964 )  ;
assign n11966 = ~ ( n10430 ) ;
assign n11967 =  ( n11965 ) | ( n11966 )  ;
assign n11968 =  ( n11967 ) | ( n10467 )  ;
assign n11969 = ~ ( n10538 ) ;
assign n11970 =  ( n11968 ) | ( n11969 )  ;
assign n11971 = ~ ( n11970 ) ;
assign n11972 =  ( n11963 ) | ( n11971 )  ;
assign n11973 = ~ ( n10358 ) ;
assign n11974 =  ( n10274 ) | ( n11973 )  ;
assign n11975 = ~ ( n10430 ) ;
assign n11976 =  ( n11974 ) | ( n11975 )  ;
assign n11977 =  ( n11976 ) | ( n10467 )  ;
assign n11978 =  ( n11977 ) | ( n10489 )  ;
assign n11979 =  ( n11978 ) | ( n10550 )  ;
assign n11980 =  ( n7455 ) ^ ( n10522 )  ;
assign n11981 =  ( n11980 ) ^ ( n10519 )  ;
assign n11982 = ~ ( n11981 ) ;
assign n11983 =  ( n11979 ) | ( n11982 )  ;
assign n11984 = ~ ( n7455 ) ;
assign n11985 =  ( n11983 ) | ( n11984 )  ;
assign n11986 = ~ ( n10564 ) ;
assign n11987 =  ( n11985 ) | ( n11986 )  ;
assign n11988 = kd[1:1] ;
assign n11989 = ~ ( n11988 ) ;
assign n11990 =  ( n11987 ) | ( n11989 )  ;
assign n11991 = ~ ( n11990 ) ;
assign n11992 =  ( n11972 ) | ( n11991 )  ;
assign n11993 = ~ ( n11992 ) ;
assign n11994 =  ( n11954 ) | ( n11993 )  ;
assign n11995 = ~ ( n11994 ) ;
assign n11996 =  ( n11926 ) | ( n11995 )  ;
assign n11997 = ~ ( n11996 ) ;
assign n11998 =  ( n6314 ) | ( n11997 )  ;
assign n11999 = ~ ( n11998 ) ;
assign n12000 =  ( n11826 ) ^ ( n11999 )  ;
assign n12001 = ~ ( n12000 ) ;
assign n12002 =  ( n11811 ) | ( n12001 )  ;
assign n12003 = ~ ( n12002 ) ;
assign n12004 =  ( n666 ) ^ ( n682 )  ;
assign n12005 =  ( n12004 ) ^ ( n697 )  ;
assign n12006 =  ( n12005 ) ^ ( n759 )  ;
assign n12007 =  ( n763 ) | ( n12006 )  ;
assign n12008 =  ( n1212 ) ^ ( n12007 )  ;
assign n12009 =  ( n12008 ) ^ ( n778 )  ;
assign n12010 =  ( n586 ) | ( n595 )  ;
assign n12011 =  ( n12010 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n12012 = ~ ( n12011 ) ;
assign n12013 =  ( n12009 ) ^ ( n12012 )  ;
assign n12014 =  ( n12013 ) ^ ( n796 )  ;
assign n12015 =  ( n12014 ) ^ ( n803 )  ;
assign n12016 =  ( n12015 ) ^ ( n11809 )  ;
assign n12017 =  ( n12016 ) ^ ( n6264 )  ;
assign n12018 =  ( n12017 ) ^ ( n5894 )  ;
assign n12019 = ~ ( n5902 ) ;
assign n12020 = ~ ( n5913 ) ;
assign n12021 =  ( n12019 ) | ( n12020 )  ;
assign n12022 =  ( n12018 ) ^ ( n12021 )  ;
assign n12023 =  ( n5832 ) | ( n5841 )  ;
assign n12024 =  ( n12023 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12025 = ~ ( n12024 ) ;
assign n12026 =  ( n12022 ) ^ ( n12025 )  ;
assign n12027 =  ( n5682 ) | ( n5691 )  ;
assign n12028 =  ( n12027 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12029 =  ( n12026 ) ^ ( n12028 )  ;
assign n12030 =  ( n5713 ) | ( n5722 )  ;
assign n12031 =  ( n12030 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12032 =  ( n12029 ) ^ ( n12031 )  ;
assign n12033 = ~ ( n11996 ) ;
assign n12034 =  ( n6314 ) | ( n12033 )  ;
assign n12035 = ~ ( n12034 ) ;
assign n12036 =  ( n12032 ) ^ ( n12035 )  ;
assign n12037 = ~ ( n12036 ) ;
assign n12038 =  ( bv_1_1_n5 ) ^ ( n1183 )  ;
assign n12039 =  ( n12038 ) ^ ( n1199 )  ;
assign n12040 =  ( n12039 ) ^ ( n666 )  ;
assign n12041 =  ( n12040 ) ^ ( n682 )  ;
assign n12042 =  ( n12041 ) ^ ( n697 )  ;
assign n12043 =  ( n12042 ) ^ ( n759 )  ;
assign n12044 =  ( n12043 ) ^ ( n11806 )  ;
assign n12045 = ~ ( n12044 ) ;
assign n12046 =  ( n12037 ) | ( n12045 )  ;
assign n12047 =  ( bv_1_1_n5 ) ^ ( n6216 )  ;
assign n12048 =  ( n12047 ) ^ ( n6242 )  ;
assign n12049 = ~ ( n5855 ) ;
assign n12050 = ~ ( n5867 ) ;
assign n12051 =  ( n12049 ) | ( n12050 )  ;
assign n12052 =  ( n12048 ) ^ ( n12051 )  ;
assign n12053 =  ( n5832 ) | ( n5841 )  ;
assign n12054 =  ( n12053 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12055 =  ( n12052 ) ^ ( n12054 )  ;
assign n12056 =  ( n5682 ) | ( n5691 )  ;
assign n12057 =  ( n12056 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12058 =  ( n12055 ) ^ ( n12057 )  ;
assign n12059 =  ( n5713 ) | ( n5722 )  ;
assign n12060 =  ( n12059 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12061 =  ( n12058 ) ^ ( n12060 )  ;
assign n12062 =  ( n12061 ) ^ ( n11996 )  ;
assign n12063 = ~ ( n12062 ) ;
assign n12064 =  ( n12046 ) | ( n12063 )  ;
assign n12065 = ~ ( n12064 ) ;
assign n12066 =  ( n12003 ) | ( n12065 )  ;
assign n12067 = ~ ( n12036 ) ;
assign n12068 =  ( n1183 ) ^ ( n1199 )  ;
assign n12069 =  ( n12068 ) ^ ( n666 )  ;
assign n12070 =  ( n12069 ) ^ ( n682 )  ;
assign n12071 =  ( n12070 ) ^ ( n697 )  ;
assign n12072 =  ( n12071 ) ^ ( n759 )  ;
assign n12073 =  ( n12072 ) ^ ( n11806 )  ;
assign n12074 =  ( n12073 ) ^ ( n6216 )  ;
assign n12075 =  ( n12074 ) ^ ( n6242 )  ;
assign n12076 = ~ ( n5855 ) ;
assign n12077 = ~ ( n5867 ) ;
assign n12078 =  ( n12076 ) | ( n12077 )  ;
assign n12079 =  ( n12075 ) ^ ( n12078 )  ;
assign n12080 =  ( n5832 ) | ( n5841 )  ;
assign n12081 =  ( n12080 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12082 =  ( n12079 ) ^ ( n12081 )  ;
assign n12083 =  ( n5682 ) | ( n5691 )  ;
assign n12084 =  ( n12083 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12085 =  ( n12082 ) ^ ( n12084 )  ;
assign n12086 =  ( n5713 ) | ( n5722 )  ;
assign n12087 =  ( n12086 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12088 =  ( n12085 ) ^ ( n12087 )  ;
assign n12089 =  ( n12088 ) ^ ( n11996 )  ;
assign n12090 = ~ ( n12089 ) ;
assign n12091 =  ( n12067 ) | ( n12090 )  ;
assign n12092 =  ( n1436 ) ^ ( n1125 )  ;
assign n12093 =  ( n12092 ) ^ ( n1145 )  ;
assign n12094 =  ( n12093 ) ^ ( n1154 )  ;
assign n12095 =  ( n532 ) | ( n541 )  ;
assign n12096 =  ( n12095 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n12097 = ~ ( n12096 ) ;
assign n12098 =  ( n12094 ) ^ ( n12097 )  ;
assign n12099 =  ( n12098 ) ^ ( n624 )  ;
assign n12100 =  ( n12099 ) ^ ( n662 )  ;
assign n12101 =  ( n12100 ) ^ ( n1179 )  ;
assign n12102 = ~ ( n1773 ) ;
assign n12103 =  ( n12102 ) | ( n1783 )  ;
assign n12104 = ~ ( n12103 ) ;
assign n12105 = ~ ( n2070 ) ;
assign n12106 =  ( n12105 ) | ( n2080 )  ;
assign n12107 = ~ ( n2092 ) ;
assign n12108 =  ( n12106 ) | ( n12107 )  ;
assign n12109 = ~ ( n12108 ) ;
assign n12110 = ~ ( n2110 ) ;
assign n12111 = ~ ( n2426 ) ;
assign n12112 =  ( n12110 ) | ( n12111 )  ;
assign n12113 =  ( n12112 ) | ( n2438 )  ;
assign n12114 = ~ ( n12113 ) ;
assign n12115 =  ( n12109 ) | ( n12114 )  ;
assign n12116 = ~ ( n2110 ) ;
assign n12117 =  ( n12116 ) | ( n2453 )  ;
assign n12118 = ~ ( n3062 ) ;
assign n12119 =  ( n12117 ) | ( n12118 )  ;
assign n12120 = ~ ( n12119 ) ;
assign n12121 =  ( n12115 ) | ( n12120 )  ;
assign n12122 =  ( n12121 ) | ( n4189 )  ;
assign n12123 = ~ ( n2110 ) ;
assign n12124 =  ( n12123 ) | ( n2453 )  ;
assign n12125 = ~ ( n2742 ) ;
assign n12126 =  ( n12124 ) | ( n12125 )  ;
assign n12127 =  ( n12126 ) | ( n3085 )  ;
assign n12128 = ~ ( n3392 ) ;
assign n12129 =  ( n12127 ) | ( n12128 )  ;
assign n12130 =  ( n12129 ) | ( n3672 )  ;
assign n12131 =  ( n12130 ) | ( n3985 )  ;
assign n12132 =  ( n12131 ) | ( n4253 )  ;
assign n12133 = ~ ( n4435 ) ;
assign n12134 = ~ ( n4689 ) ;
assign n12135 =  ( n12133 ) | ( n12134 )  ;
assign n12136 =  ( n4458 ) | ( n4710 )  ;
assign n12137 = ~ ( n4916 ) ;
assign n12138 =  ( n12136 ) | ( n12137 )  ;
assign n12139 = ~ ( n12138 ) ;
assign n12140 =  ( n12135 ) | ( n12139 )  ;
assign n12141 =  ( n12140 ) | ( n5349 )  ;
assign n12142 = ~ ( n12141 ) ;
assign n12143 =  ( n12132 ) | ( n12142 )  ;
assign n12144 = ~ ( n12143 ) ;
assign n12145 =  ( n12122 ) | ( n12144 )  ;
assign n12146 = ~ ( n2110 ) ;
assign n12147 =  ( n12146 ) | ( n2453 )  ;
assign n12148 = ~ ( n2742 ) ;
assign n12149 =  ( n12147 ) | ( n12148 )  ;
assign n12150 =  ( n12149 ) | ( n3085 )  ;
assign n12151 = ~ ( n3392 ) ;
assign n12152 =  ( n12150 ) | ( n12151 )  ;
assign n12153 =  ( n12152 ) | ( n3672 )  ;
assign n12154 =  ( n12153 ) | ( n3985 )  ;
assign n12155 =  ( n12154 ) | ( n4253 )  ;
assign n12156 =  ( n12155 ) | ( n4458 )  ;
assign n12157 =  ( n12156 ) | ( n4710 )  ;
assign n12158 = ~ ( n4763 ) ;
assign n12159 =  ( n12157 ) | ( n12158 )  ;
assign n12160 = ~ ( n4938 ) ;
assign n12161 =  ( n12159 ) | ( n12160 )  ;
assign n12162 =  ( n12161 ) | ( n5063 )  ;
assign n12163 =  ( n12162 ) | ( n5224 )  ;
assign n12164 =  ( n12163 ) | ( n5265 )  ;
assign n12165 =  ( n5366 ) ^ ( n5161 )  ;
assign n12166 =  ( n12165 ) ^ ( n5171 )  ;
assign n12167 =  ( n12166 ) ^ ( n4960 )  ;
assign n12168 =  ( n12167 ) ^ ( n4976 )  ;
assign n12169 =  ( n12168 ) ^ ( n4996 )  ;
assign n12170 =  ( n12169 ) ^ ( n5236 )  ;
assign n12171 = ~ ( n12170 ) ;
assign n12172 =  ( n12164 ) | ( n12171 )  ;
assign n12173 =  ( n5446 ) | ( n5473 )  ;
assign n12174 =  ( n12173 ) | ( n5604 )  ;
assign n12175 =  ( n12174 ) | ( n5663 )  ;
assign n12176 = ~ ( n12175 ) ;
assign n12177 =  ( n12172 ) | ( n12176 )  ;
assign n12178 = ~ ( n12177 ) ;
assign n12179 =  ( n12145 ) | ( n12178 )  ;
assign n12180 = ~ ( n12179 ) ;
assign n12181 =  ( n1828 ) | ( n12180 )  ;
assign n12182 = ~ ( n12181 ) ;
assign n12183 =  ( n12104 ) | ( n12182 )  ;
assign n12184 =  ( n12101 ) ^ ( n12183 )  ;
assign n12185 = ~ ( n12184 ) ;
assign n12186 = ~ ( n6402 ) ;
assign n12187 =  ( n12186 ) | ( n6421 )  ;
assign n12188 = ~ ( n12187 ) ;
assign n12189 = ~ ( n6105 ) ;
assign n12190 =  ( n6111 ) | ( n6124 )  ;
assign n12191 = ~ ( n12190 ) ;
assign n12192 =  ( n12189 ) | ( n12191 )  ;
assign n12193 =  ( n12188 ) ^ ( n12192 )  ;
assign n12194 =  ( n12193 ) ^ ( n6166 )  ;
assign n12195 = ~ ( n6173 ) ;
assign n12196 = ~ ( n5736 ) ;
assign n12197 =  ( n12195 ) | ( n12196 )  ;
assign n12198 =  ( n12194 ) ^ ( n12197 )  ;
assign n12199 =  ( n5802 ) | ( n5811 )  ;
assign n12200 =  ( n12199 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12201 = ~ ( n12200 ) ;
assign n12202 =  ( n12198 ) ^ ( n12201 )  ;
assign n12203 =  ( n5832 ) | ( n5841 )  ;
assign n12204 =  ( n12203 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12205 =  ( n12202 ) ^ ( n12204 )  ;
assign n12206 =  ( n5682 ) | ( n5691 )  ;
assign n12207 =  ( n12206 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12208 =  ( n12205 ) ^ ( n12207 )  ;
assign n12209 =  ( n5713 ) | ( n5722 )  ;
assign n12210 =  ( n12209 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12211 =  ( n12208 ) ^ ( n12210 )  ;
assign n12212 = ~ ( n6753 ) ;
assign n12213 =  ( n12212 ) | ( n6774 )  ;
assign n12214 = ~ ( n12213 ) ;
assign n12215 = ~ ( n7022 ) ;
assign n12216 =  ( n12215 ) | ( n7045 )  ;
assign n12217 = ~ ( n7078 ) ;
assign n12218 =  ( n12216 ) | ( n12217 )  ;
assign n12219 = ~ ( n12218 ) ;
assign n12220 = ~ ( n7117 ) ;
assign n12221 = ~ ( n7392 ) ;
assign n12222 =  ( n12220 ) | ( n12221 )  ;
assign n12223 =  ( n12222 ) | ( n7417 )  ;
assign n12224 = ~ ( n12223 ) ;
assign n12225 =  ( n12219 ) | ( n12224 )  ;
assign n12226 = ~ ( n7117 ) ;
assign n12227 =  ( n12226 ) | ( n7445 )  ;
assign n12228 = ~ ( n8082 ) ;
assign n12229 =  ( n12227 ) | ( n12228 )  ;
assign n12230 = ~ ( n12229 ) ;
assign n12231 =  ( n12225 ) | ( n12230 )  ;
assign n12232 =  ( n12231 ) | ( n9179 )  ;
assign n12233 = ~ ( n7117 ) ;
assign n12234 =  ( n12233 ) | ( n7445 )  ;
assign n12235 = ~ ( n7765 ) ;
assign n12236 =  ( n12234 ) | ( n12235 )  ;
assign n12237 =  ( n12236 ) | ( n8121 )  ;
assign n12238 = ~ ( n8413 ) ;
assign n12239 =  ( n12237 ) | ( n12238 )  ;
assign n12240 = ~ ( n8717 ) ;
assign n12241 =  ( n12239 ) | ( n12240 )  ;
assign n12242 = ~ ( n9012 ) ;
assign n12243 =  ( n12241 ) | ( n12242 )  ;
assign n12244 = ~ ( n9252 ) ;
assign n12245 =  ( n12243 ) | ( n12244 )  ;
assign n12246 = ~ ( n9314 ) ;
assign n12247 = ~ ( n9348 ) ;
assign n12248 =  ( n12246 ) | ( n12247 )  ;
assign n12249 = ~ ( n9387 ) ;
assign n12250 =  ( n12248 ) | ( n12249 )  ;
assign n12251 = ~ ( n12250 ) ;
assign n12252 =  ( n12251 ) | ( n9608 )  ;
assign n12253 = ~ ( n9432 ) ;
assign n12254 = ~ ( n9649 ) ;
assign n12255 =  ( n12253 ) | ( n12254 )  ;
assign n12256 = ~ ( n9868 ) ;
assign n12257 =  ( n12255 ) | ( n12256 )  ;
assign n12258 = ~ ( n12257 ) ;
assign n12259 =  ( n12252 ) | ( n12258 )  ;
assign n12260 =  ( n12259 ) | ( n10319 )  ;
assign n12261 = ~ ( n12260 ) ;
assign n12262 =  ( n12245 ) | ( n12261 )  ;
assign n12263 = ~ ( n12262 ) ;
assign n12264 =  ( n12232 ) | ( n12263 )  ;
assign n12265 = ~ ( n7117 ) ;
assign n12266 =  ( n12265 ) | ( n7445 )  ;
assign n12267 = ~ ( n7765 ) ;
assign n12268 =  ( n12266 ) | ( n12267 )  ;
assign n12269 =  ( n12268 ) | ( n8121 )  ;
assign n12270 = ~ ( n8413 ) ;
assign n12271 =  ( n12269 ) | ( n12270 )  ;
assign n12272 = ~ ( n8717 ) ;
assign n12273 =  ( n12271 ) | ( n12272 )  ;
assign n12274 = ~ ( n9012 ) ;
assign n12275 =  ( n12273 ) | ( n12274 )  ;
assign n12276 = ~ ( n9252 ) ;
assign n12277 =  ( n12275 ) | ( n12276 )  ;
assign n12278 = ~ ( n9432 ) ;
assign n12279 =  ( n12277 ) | ( n12278 )  ;
assign n12280 = ~ ( n9649 ) ;
assign n12281 =  ( n12279 ) | ( n12280 )  ;
assign n12282 = ~ ( n9751 ) ;
assign n12283 =  ( n12281 ) | ( n12282 )  ;
assign n12284 = ~ ( n9909 ) ;
assign n12285 =  ( n12283 ) | ( n12284 )  ;
assign n12286 = ~ ( n10042 ) ;
assign n12287 =  ( n12285 ) | ( n12286 )  ;
assign n12288 = ~ ( n10208 ) ;
assign n12289 =  ( n12287 ) | ( n12288 )  ;
assign n12290 =  ( n12289 ) | ( n10274 )  ;
assign n12291 = ~ ( n10358 ) ;
assign n12292 =  ( n12290 ) | ( n12291 )  ;
assign n12293 = ~ ( n10571 ) ;
assign n12294 =  ( n12292 ) | ( n12293 )  ;
assign n12295 = ~ ( n12294 ) ;
assign n12296 =  ( n12264 ) | ( n12295 )  ;
assign n12297 = ~ ( n12296 ) ;
assign n12298 =  ( n6815 ) | ( n12297 )  ;
assign n12299 = ~ ( n12298 ) ;
assign n12300 =  ( n12214 ) | ( n12299 )  ;
assign n12301 =  ( n12211 ) ^ ( n12300 )  ;
assign n12302 = ~ ( n12301 ) ;
assign n12303 =  ( n12185 ) | ( n12302 )  ;
assign n12304 = ~ ( n12303 ) ;
assign n12305 =  ( n1436 ) ^ ( n1125 )  ;
assign n12306 =  ( n12305 ) ^ ( n1145 )  ;
assign n12307 =  ( n12306 ) ^ ( n1154 )  ;
assign n12308 =  ( n532 ) | ( n541 )  ;
assign n12309 =  ( n12308 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n12310 = ~ ( n12309 ) ;
assign n12311 =  ( n12307 ) ^ ( n12310 )  ;
assign n12312 =  ( n12311 ) ^ ( n624 )  ;
assign n12313 =  ( n12312 ) ^ ( n662 )  ;
assign n12314 =  ( n12313 ) ^ ( n1179 )  ;
assign n12315 =  ( n12314 ) ^ ( n12183 )  ;
assign n12316 = ~ ( n6402 ) ;
assign n12317 =  ( n12316 ) | ( n6421 )  ;
assign n12318 = ~ ( n12317 ) ;
assign n12319 =  ( n12315 ) ^ ( n12318 )  ;
assign n12320 = ~ ( n6105 ) ;
assign n12321 =  ( n6111 ) | ( n6124 )  ;
assign n12322 = ~ ( n12321 ) ;
assign n12323 =  ( n12320 ) | ( n12322 )  ;
assign n12324 =  ( n12319 ) ^ ( n12323 )  ;
assign n12325 =  ( n12324 ) ^ ( n6166 )  ;
assign n12326 = ~ ( n6173 ) ;
assign n12327 = ~ ( n5736 ) ;
assign n12328 =  ( n12326 ) | ( n12327 )  ;
assign n12329 =  ( n12325 ) ^ ( n12328 )  ;
assign n12330 =  ( n5802 ) | ( n5811 )  ;
assign n12331 =  ( n12330 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12332 = ~ ( n12331 ) ;
assign n12333 =  ( n12329 ) ^ ( n12332 )  ;
assign n12334 =  ( n5832 ) | ( n5841 )  ;
assign n12335 =  ( n12334 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12336 =  ( n12333 ) ^ ( n12335 )  ;
assign n12337 =  ( n5682 ) | ( n5691 )  ;
assign n12338 =  ( n12337 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12339 =  ( n12336 ) ^ ( n12338 )  ;
assign n12340 =  ( n5713 ) | ( n5722 )  ;
assign n12341 =  ( n12340 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12342 =  ( n12339 ) ^ ( n12341 )  ;
assign n12343 =  ( n12342 ) ^ ( n12300 )  ;
assign n12344 = ~ ( n12343 ) ;
assign n12345 =  ( bv_1_1_n5 ) ^ ( n1773 )  ;
assign n12346 =  ( n12345 ) ^ ( n1405 )  ;
assign n12347 =  ( n12346 ) ^ ( n1068 )  ;
assign n12348 =  ( n12347 ) ^ ( n1079 )  ;
assign n12349 =  ( n12348 ) ^ ( n1090 )  ;
assign n12350 =  ( n12349 ) ^ ( n1097 )  ;
assign n12351 =  ( n12350 ) ^ ( n1104 )  ;
assign n12352 =  ( n12351 ) ^ ( n1120 )  ;
assign n12353 =  ( n12352 ) ^ ( n12179 )  ;
assign n12354 = ~ ( n12353 ) ;
assign n12355 =  ( n12344 ) | ( n12354 )  ;
assign n12356 =  ( bv_1_1_n5 ) ^ ( n6753 )  ;
assign n12357 =  ( n12356 ) ^ ( n6402 )  ;
assign n12358 =  ( n12357 ) ^ ( n6093 )  ;
assign n12359 = ~ ( n6100 ) ;
assign n12360 = ~ ( n5902 ) ;
assign n12361 =  ( n12359 ) | ( n12360 )  ;
assign n12362 =  ( n12358 ) ^ ( n12361 )  ;
assign n12363 =  ( n5802 ) | ( n5811 )  ;
assign n12364 =  ( n12363 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12365 =  ( n12362 ) ^ ( n12364 )  ;
assign n12366 =  ( n5832 ) | ( n5841 )  ;
assign n12367 =  ( n12366 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12368 =  ( n12365 ) ^ ( n12367 )  ;
assign n12369 =  ( n5682 ) | ( n5691 )  ;
assign n12370 =  ( n12369 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12371 =  ( n12368 ) ^ ( n12370 )  ;
assign n12372 =  ( n5713 ) | ( n5722 )  ;
assign n12373 =  ( n12372 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12374 =  ( n12371 ) ^ ( n12373 )  ;
assign n12375 =  ( n12374 ) ^ ( n12296 )  ;
assign n12376 = ~ ( n12375 ) ;
assign n12377 =  ( n12355 ) | ( n12376 )  ;
assign n12378 = ~ ( n12377 ) ;
assign n12379 =  ( n12304 ) | ( n12378 )  ;
assign n12380 = ~ ( n12379 ) ;
assign n12381 =  ( n12091 ) | ( n12380 )  ;
assign n12382 = ~ ( n12381 ) ;
assign n12383 =  ( n12066 ) | ( n12382 )  ;
assign n12384 = ~ ( n12383 ) ;
assign n12385 =  ( n11620 ) | ( n12384 )  ;
assign n12386 = ~ ( n12385 ) ;
assign n12387 =  ( n11598 ) | ( n12386 )  ;
assign n12388 = ~ ( n11115 ) ;
assign n12389 =  ( n12388 ) | ( n11145 )  ;
assign n12390 = ~ ( n11570 ) ;
assign n12391 =  ( n12389 ) | ( n12390 )  ;
assign n12392 =  ( n12391 ) | ( n11619 )  ;
assign n12393 = ~ ( n12036 ) ;
assign n12394 =  ( n12392 ) | ( n12393 )  ;
assign n12395 =  ( n12394 ) | ( n12090 )  ;
assign n12396 = ~ ( n12343 ) ;
assign n12397 =  ( n12395 ) | ( n12396 )  ;
assign n12398 =  ( n1773 ) ^ ( n1405 )  ;
assign n12399 =  ( n12398 ) ^ ( n1068 )  ;
assign n12400 =  ( n12399 ) ^ ( n1079 )  ;
assign n12401 =  ( n12400 ) ^ ( n1090 )  ;
assign n12402 =  ( n12401 ) ^ ( n1097 )  ;
assign n12403 =  ( n12402 ) ^ ( n1104 )  ;
assign n12404 =  ( n12403 ) ^ ( n1120 )  ;
assign n12405 =  ( n12404 ) ^ ( n12179 )  ;
assign n12406 =  ( n12405 ) ^ ( n6753 )  ;
assign n12407 =  ( n12406 ) ^ ( n6402 )  ;
assign n12408 =  ( n12407 ) ^ ( n6093 )  ;
assign n12409 = ~ ( n6100 ) ;
assign n12410 = ~ ( n5902 ) ;
assign n12411 =  ( n12409 ) | ( n12410 )  ;
assign n12412 =  ( n12408 ) ^ ( n12411 )  ;
assign n12413 =  ( n5802 ) | ( n5811 )  ;
assign n12414 =  ( n12413 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12415 =  ( n12412 ) ^ ( n12414 )  ;
assign n12416 =  ( n5832 ) | ( n5841 )  ;
assign n12417 =  ( n12416 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12418 =  ( n12415 ) ^ ( n12417 )  ;
assign n12419 =  ( n5682 ) | ( n5691 )  ;
assign n12420 =  ( n12419 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12421 =  ( n12418 ) ^ ( n12420 )  ;
assign n12422 =  ( n5713 ) | ( n5722 )  ;
assign n12423 =  ( n12422 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12424 =  ( n12421 ) ^ ( n12423 )  ;
assign n12425 =  ( n12424 ) ^ ( n12296 )  ;
assign n12426 = ~ ( n12425 ) ;
assign n12427 =  ( n12397 ) | ( n12426 )  ;
assign n12428 = ~ ( n2070 ) ;
assign n12429 =  ( n12428 ) | ( n2080 )  ;
assign n12430 = ~ ( n12429 ) ;
assign n12431 =  ( n12430 ) ^ ( n1740 )  ;
assign n12432 =  ( n12431 ) ^ ( n1755 )  ;
assign n12433 =  ( n12432 ) ^ ( n1379 )  ;
assign n12434 =  ( n12433 ) ^ ( n1389 )  ;
assign n12435 =  ( n873 ) | ( n882 )  ;
assign n12436 =  ( n12435 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n12437 = ~ ( n12436 ) ;
assign n12438 =  ( n12434 ) ^ ( n12437 )  ;
assign n12439 =  ( n12438 ) ^ ( n941 )  ;
assign n12440 =  ( n12439 ) ^ ( n967 )  ;
assign n12441 =  ( n12440 ) ^ ( n999 )  ;
assign n12442 =  ( n12441 ) ^ ( n1064 )  ;
assign n12443 = ~ ( n2426 ) ;
assign n12444 =  ( n12443 ) | ( n2438 )  ;
assign n12445 = ~ ( n12444 ) ;
assign n12446 = ~ ( n2722 ) ;
assign n12447 = ~ ( n2742 ) ;
assign n12448 = ~ ( n3043 ) ;
assign n12449 =  ( n12447 ) | ( n12448 )  ;
assign n12450 =  ( n12449 ) | ( n3059 )  ;
assign n12451 = ~ ( n12450 ) ;
assign n12452 =  ( n12446 ) | ( n12451 )  ;
assign n12453 = ~ ( n2742 ) ;
assign n12454 =  ( n12453 ) | ( n3085 )  ;
assign n12455 = ~ ( n10688 ) ;
assign n12456 =  ( n12454 ) | ( n12455 )  ;
assign n12457 = ~ ( n12456 ) ;
assign n12458 =  ( n12452 ) | ( n12457 )  ;
assign n12459 = ~ ( n10709 ) ;
assign n12460 =  ( n12458 ) | ( n12459 )  ;
assign n12461 = ~ ( n2742 ) ;
assign n12462 =  ( n12461 ) | ( n3085 )  ;
assign n12463 = ~ ( n3392 ) ;
assign n12464 =  ( n12462 ) | ( n12463 )  ;
assign n12465 =  ( n12464 ) | ( n3672 )  ;
assign n12466 =  ( n12465 ) | ( n3985 )  ;
assign n12467 =  ( n12466 ) | ( n4253 )  ;
assign n12468 =  ( n12467 ) | ( n4458 )  ;
assign n12469 =  ( n12468 ) | ( n4710 )  ;
assign n12470 = ~ ( n4728 ) ;
assign n12471 =  ( n4722 ) | ( n12470 )  ;
assign n12472 =  ( n12471 ) | ( n4744 )  ;
assign n12473 = ~ ( n12472 ) ;
assign n12474 = ~ ( n4763 ) ;
assign n12475 = ~ ( n4889 ) ;
assign n12476 =  ( n12474 ) | ( n12475 )  ;
assign n12477 =  ( n12476 ) | ( n4900 )  ;
assign n12478 =  ( n12477 ) | ( n4913 )  ;
assign n12479 = ~ ( n12478 ) ;
assign n12480 =  ( n12473 ) | ( n12479 )  ;
assign n12481 =  ( n12480 ) | ( n10766 )  ;
assign n12482 =  ( n12481 ) | ( n10789 )  ;
assign n12483 = ~ ( n12482 ) ;
assign n12484 =  ( n12469 ) | ( n12483 )  ;
assign n12485 = ~ ( n12484 ) ;
assign n12486 =  ( n12460 ) | ( n12485 )  ;
assign n12487 = ~ ( n2742 ) ;
assign n12488 =  ( n12487 ) | ( n3085 )  ;
assign n12489 = ~ ( n3392 ) ;
assign n12490 =  ( n12488 ) | ( n12489 )  ;
assign n12491 =  ( n12490 ) | ( n3672 )  ;
assign n12492 =  ( n12491 ) | ( n3985 )  ;
assign n12493 =  ( n12492 ) | ( n4253 )  ;
assign n12494 =  ( n12493 ) | ( n4458 )  ;
assign n12495 =  ( n12494 ) | ( n4710 )  ;
assign n12496 = ~ ( n4763 ) ;
assign n12497 =  ( n12495 ) | ( n12496 )  ;
assign n12498 = ~ ( n4938 ) ;
assign n12499 =  ( n12497 ) | ( n12498 )  ;
assign n12500 =  ( n12499 ) | ( n5063 )  ;
assign n12501 =  ( n12500 ) | ( n5224 )  ;
assign n12502 =  ( n12501 ) | ( n5265 )  ;
assign n12503 =  ( n5366 ) ^ ( n5161 )  ;
assign n12504 =  ( n12503 ) ^ ( n5171 )  ;
assign n12505 =  ( n12504 ) ^ ( n4960 )  ;
assign n12506 =  ( n12505 ) ^ ( n4976 )  ;
assign n12507 =  ( n12506 ) ^ ( n4996 )  ;
assign n12508 =  ( n12507 ) ^ ( n5236 )  ;
assign n12509 = ~ ( n12508 ) ;
assign n12510 =  ( n12502 ) | ( n12509 )  ;
assign n12511 =  ( n5452 ) ^ ( n5325 )  ;
assign n12512 =  ( n12511 ) ^ ( n5083 )  ;
assign n12513 =  ( n12512 ) ^ ( n5099 )  ;
assign n12514 =  ( n12513 ) ^ ( n5116 )  ;
assign n12515 =  ( n12514 ) ^ ( n5141 )  ;
assign n12516 =  ( n12515 ) ^ ( n5129 )  ;
assign n12517 = ~ ( n12516 ) ;
assign n12518 =  ( n12510 ) | ( n12517 )  ;
assign n12519 =  ( n5489 ) ^ ( n5433 )  ;
assign n12520 =  ( n12519 ) ^ ( n5285 )  ;
assign n12521 =  ( n12520 ) ^ ( n5301 )  ;
assign n12522 =  ( n12521 ) ^ ( n5321 )  ;
assign n12523 = ~ ( n12522 ) ;
assign n12524 =  ( n12518 ) | ( n12523 )  ;
assign n12525 =  ( n5539 ) | ( n5600 )  ;
assign n12526 =  ( n12525 ) | ( n10836 )  ;
assign n12527 = ~ ( n12526 ) ;
assign n12528 =  ( n12524 ) | ( n12527 )  ;
assign n12529 = ~ ( n12528 ) ;
assign n12530 =  ( n12486 ) | ( n12529 )  ;
assign n12531 = ~ ( n12530 ) ;
assign n12532 =  ( n2453 ) | ( n12531 )  ;
assign n12533 = ~ ( n12532 ) ;
assign n12534 =  ( n12445 ) | ( n12533 )  ;
assign n12535 =  ( n12442 ) ^ ( n12534 )  ;
assign n12536 = ~ ( n12535 ) ;
assign n12537 = ~ ( n7022 ) ;
assign n12538 =  ( n12537 ) | ( n7045 )  ;
assign n12539 = ~ ( n12538 ) ;
assign n12540 =  ( n12539 ) ^ ( n6683 )  ;
assign n12541 = ~ ( n6690 ) ;
assign n12542 =  ( n6696 ) | ( n6711 )  ;
assign n12543 = ~ ( n12542 ) ;
assign n12544 =  ( n12541 ) | ( n12543 )  ;
assign n12545 =  ( n12540 ) ^ ( n12544 )  ;
assign n12546 = ~ ( n6330 ) ;
assign n12547 =  ( n6337 ) | ( n5909 )  ;
assign n12548 = ~ ( n12547 ) ;
assign n12549 =  ( n12546 ) | ( n12548 )  ;
assign n12550 = ~ ( n6356 ) ;
assign n12551 =  ( n12549 ) | ( n12550 )  ;
assign n12552 =  ( n12545 ) ^ ( n12551 )  ;
assign n12553 = ~ ( n6366 ) ;
assign n12554 = ~ ( n5902 ) ;
assign n12555 =  ( n12553 ) | ( n12554 )  ;
assign n12556 =  ( n12552 ) ^ ( n12555 )  ;
assign n12557 =  ( n6030 ) | ( n6039 )  ;
assign n12558 =  ( n12557 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n12559 = ~ ( n12558 ) ;
assign n12560 =  ( n12556 ) ^ ( n12559 )  ;
assign n12561 =  ( n5802 ) | ( n5811 )  ;
assign n12562 =  ( n12561 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12563 =  ( n12560 ) ^ ( n12562 )  ;
assign n12564 =  ( n5832 ) | ( n5841 )  ;
assign n12565 =  ( n12564 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12566 =  ( n12563 ) ^ ( n12565 )  ;
assign n12567 =  ( n5682 ) | ( n5691 )  ;
assign n12568 =  ( n12567 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12569 =  ( n12566 ) ^ ( n12568 )  ;
assign n12570 =  ( n5713 ) | ( n5722 )  ;
assign n12571 =  ( n12570 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12572 =  ( n12569 ) ^ ( n12571 )  ;
assign n12573 = ~ ( n7392 ) ;
assign n12574 =  ( n12573 ) | ( n7417 )  ;
assign n12575 = ~ ( n12574 ) ;
assign n12576 = ~ ( n7649 ) ;
assign n12577 =  ( n12576 ) | ( n7679 )  ;
assign n12578 = ~ ( n7719 ) ;
assign n12579 =  ( n12577 ) | ( n12578 )  ;
assign n12580 = ~ ( n12579 ) ;
assign n12581 = ~ ( n7765 ) ;
assign n12582 = ~ ( n8047 ) ;
assign n12583 =  ( n12581 ) | ( n12582 )  ;
assign n12584 =  ( n12583 ) | ( n8079 )  ;
assign n12585 = ~ ( n12584 ) ;
assign n12586 =  ( n12580 ) | ( n12585 )  ;
assign n12587 = ~ ( n7765 ) ;
assign n12588 =  ( n12587 ) | ( n8121 )  ;
assign n12589 = ~ ( n10939 ) ;
assign n12590 =  ( n12588 ) | ( n12589 )  ;
assign n12591 = ~ ( n12590 ) ;
assign n12592 =  ( n12586 ) | ( n12591 )  ;
assign n12593 =  ( n12592 ) | ( n10973 )  ;
assign n12594 = ~ ( n7765 ) ;
assign n12595 =  ( n12594 ) | ( n8121 )  ;
assign n12596 = ~ ( n8413 ) ;
assign n12597 =  ( n12595 ) | ( n12596 )  ;
assign n12598 = ~ ( n8717 ) ;
assign n12599 =  ( n12597 ) | ( n12598 )  ;
assign n12600 = ~ ( n9012 ) ;
assign n12601 =  ( n12599 ) | ( n12600 )  ;
assign n12602 = ~ ( n9252 ) ;
assign n12603 =  ( n12601 ) | ( n12602 )  ;
assign n12604 = ~ ( n9432 ) ;
assign n12605 =  ( n12603 ) | ( n12604 )  ;
assign n12606 = ~ ( n9649 ) ;
assign n12607 =  ( n12605 ) | ( n12606 )  ;
assign n12608 = ~ ( n9713 ) ;
assign n12609 = ~ ( n9751 ) ;
assign n12610 =  ( n12609 ) | ( n9808 )  ;
assign n12611 = ~ ( n9834 ) ;
assign n12612 =  ( n12610 ) | ( n12611 )  ;
assign n12613 = ~ ( n9864 ) ;
assign n12614 =  ( n12612 ) | ( n12613 )  ;
assign n12615 = ~ ( n12614 ) ;
assign n12616 =  ( n12608 ) | ( n12615 )  ;
assign n12617 = ~ ( n9751 ) ;
assign n12618 = ~ ( n9909 ) ;
assign n12619 =  ( n12617 ) | ( n12618 )  ;
assign n12620 = ~ ( n11024 ) ;
assign n12621 =  ( n12619 ) | ( n12620 )  ;
assign n12622 = ~ ( n12621 ) ;
assign n12623 =  ( n12616 ) | ( n12622 )  ;
assign n12624 =  ( n12623 ) | ( n11052 )  ;
assign n12625 = ~ ( n12624 ) ;
assign n12626 =  ( n12607 ) | ( n12625 )  ;
assign n12627 = ~ ( n12626 ) ;
assign n12628 =  ( n12593 ) | ( n12627 )  ;
assign n12629 = ~ ( n7765 ) ;
assign n12630 =  ( n12629 ) | ( n8121 )  ;
assign n12631 = ~ ( n8413 ) ;
assign n12632 =  ( n12630 ) | ( n12631 )  ;
assign n12633 = ~ ( n8717 ) ;
assign n12634 =  ( n12632 ) | ( n12633 )  ;
assign n12635 = ~ ( n9012 ) ;
assign n12636 =  ( n12634 ) | ( n12635 )  ;
assign n12637 = ~ ( n9252 ) ;
assign n12638 =  ( n12636 ) | ( n12637 )  ;
assign n12639 = ~ ( n9432 ) ;
assign n12640 =  ( n12638 ) | ( n12639 )  ;
assign n12641 = ~ ( n9649 ) ;
assign n12642 =  ( n12640 ) | ( n12641 )  ;
assign n12643 = ~ ( n9751 ) ;
assign n12644 =  ( n12642 ) | ( n12643 )  ;
assign n12645 = ~ ( n9909 ) ;
assign n12646 =  ( n12644 ) | ( n12645 )  ;
assign n12647 = ~ ( n10042 ) ;
assign n12648 =  ( n12646 ) | ( n12647 )  ;
assign n12649 = ~ ( n10208 ) ;
assign n12650 =  ( n12648 ) | ( n12649 )  ;
assign n12651 =  ( n12650 ) | ( n10274 )  ;
assign n12652 = ~ ( n10358 ) ;
assign n12653 =  ( n12651 ) | ( n12652 )  ;
assign n12654 = ~ ( n10430 ) ;
assign n12655 =  ( n12653 ) | ( n12654 )  ;
assign n12656 =  ( n12655 ) | ( n10467 )  ;
assign n12657 = ~ ( n11086 ) ;
assign n12658 =  ( n12656 ) | ( n12657 )  ;
assign n12659 = ~ ( n12658 ) ;
assign n12660 =  ( n12628 ) | ( n12659 )  ;
assign n12661 = ~ ( n12660 ) ;
assign n12662 =  ( n7445 ) | ( n12661 )  ;
assign n12663 = ~ ( n12662 ) ;
assign n12664 =  ( n12575 ) | ( n12663 )  ;
assign n12665 =  ( n12572 ) ^ ( n12664 )  ;
assign n12666 = ~ ( n12665 ) ;
assign n12667 =  ( n12536 ) | ( n12666 )  ;
assign n12668 = ~ ( n12667 ) ;
assign n12669 = ~ ( n2070 ) ;
assign n12670 =  ( n12669 ) | ( n2080 )  ;
assign n12671 = ~ ( n12670 ) ;
assign n12672 =  ( n12671 ) ^ ( n1740 )  ;
assign n12673 =  ( n12672 ) ^ ( n1755 )  ;
assign n12674 =  ( n12673 ) ^ ( n1379 )  ;
assign n12675 =  ( n12674 ) ^ ( n1389 )  ;
assign n12676 =  ( n873 ) | ( n882 )  ;
assign n12677 =  ( n12676 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n12678 = ~ ( n12677 ) ;
assign n12679 =  ( n12675 ) ^ ( n12678 )  ;
assign n12680 =  ( n12679 ) ^ ( n941 )  ;
assign n12681 =  ( n12680 ) ^ ( n967 )  ;
assign n12682 =  ( n12681 ) ^ ( n999 )  ;
assign n12683 =  ( n12682 ) ^ ( n1064 )  ;
assign n12684 =  ( n12683 ) ^ ( n12534 )  ;
assign n12685 = ~ ( n7022 ) ;
assign n12686 =  ( n12685 ) | ( n7045 )  ;
assign n12687 = ~ ( n12686 ) ;
assign n12688 =  ( n12684 ) ^ ( n12687 )  ;
assign n12689 =  ( n12688 ) ^ ( n6683 )  ;
assign n12690 = ~ ( n6690 ) ;
assign n12691 =  ( n6696 ) | ( n6711 )  ;
assign n12692 = ~ ( n12691 ) ;
assign n12693 =  ( n12690 ) | ( n12692 )  ;
assign n12694 =  ( n12689 ) ^ ( n12693 )  ;
assign n12695 = ~ ( n6330 ) ;
assign n12696 =  ( n6337 ) | ( n5909 )  ;
assign n12697 = ~ ( n12696 ) ;
assign n12698 =  ( n12695 ) | ( n12697 )  ;
assign n12699 = ~ ( n6356 ) ;
assign n12700 =  ( n12698 ) | ( n12699 )  ;
assign n12701 =  ( n12694 ) ^ ( n12700 )  ;
assign n12702 = ~ ( n6366 ) ;
assign n12703 = ~ ( n5902 ) ;
assign n12704 =  ( n12702 ) | ( n12703 )  ;
assign n12705 =  ( n12701 ) ^ ( n12704 )  ;
assign n12706 =  ( n6030 ) | ( n6039 )  ;
assign n12707 =  ( n12706 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n12708 = ~ ( n12707 ) ;
assign n12709 =  ( n12705 ) ^ ( n12708 )  ;
assign n12710 =  ( n5802 ) | ( n5811 )  ;
assign n12711 =  ( n12710 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12712 =  ( n12709 ) ^ ( n12711 )  ;
assign n12713 =  ( n5832 ) | ( n5841 )  ;
assign n12714 =  ( n12713 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12715 =  ( n12712 ) ^ ( n12714 )  ;
assign n12716 =  ( n5682 ) | ( n5691 )  ;
assign n12717 =  ( n12716 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12718 =  ( n12715 ) ^ ( n12717 )  ;
assign n12719 =  ( n5713 ) | ( n5722 )  ;
assign n12720 =  ( n12719 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12721 =  ( n12718 ) ^ ( n12720 )  ;
assign n12722 =  ( n12721 ) ^ ( n12664 )  ;
assign n12723 = ~ ( n12722 ) ;
assign n12724 =  ( bv_1_1_n5 ) ^ ( n2426 )  ;
assign n12725 =  ( n12724 ) ^ ( n2070 )  ;
assign n12726 =  ( n12725 ) ^ ( n1682 )  ;
assign n12727 =  ( n12726 ) ^ ( n1713 )  ;
assign n12728 =  ( n12727 ) ^ ( n1723 )  ;
assign n12729 =  ( n12728 ) ^ ( n1281 )  ;
assign n12730 =  ( n12729 ) ^ ( n1297 )  ;
assign n12731 =  ( n12730 ) ^ ( n1314 )  ;
assign n12732 =  ( n12731 ) ^ ( n1331 )  ;
assign n12733 =  ( n12732 ) ^ ( n1375 )  ;
assign n12734 =  ( n12733 ) ^ ( n12530 )  ;
assign n12735 = ~ ( n12734 ) ;
assign n12736 =  ( n12723 ) | ( n12735 )  ;
assign n12737 =  ( bv_1_1_n5 ) ^ ( n7392 )  ;
assign n12738 =  ( n12737 ) ^ ( n7022 )  ;
assign n12739 =  ( n12738 ) ^ ( n6589 )  ;
assign n12740 =  ( n12739 ) ^ ( n6634 )  ;
assign n12741 = ~ ( n6640 ) ;
assign n12742 = ~ ( n6173 ) ;
assign n12743 =  ( n12741 ) | ( n12742 )  ;
assign n12744 =  ( n12740 ) ^ ( n12743 )  ;
assign n12745 =  ( n6030 ) | ( n6039 )  ;
assign n12746 =  ( n12745 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n12747 =  ( n12744 ) ^ ( n12746 )  ;
assign n12748 =  ( n5802 ) | ( n5811 )  ;
assign n12749 =  ( n12748 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12750 =  ( n12747 ) ^ ( n12749 )  ;
assign n12751 =  ( n5832 ) | ( n5841 )  ;
assign n12752 =  ( n12751 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12753 =  ( n12750 ) ^ ( n12752 )  ;
assign n12754 =  ( n5682 ) | ( n5691 )  ;
assign n12755 =  ( n12754 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12756 =  ( n12753 ) ^ ( n12755 )  ;
assign n12757 =  ( n5713 ) | ( n5722 )  ;
assign n12758 =  ( n12757 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12759 =  ( n12756 ) ^ ( n12758 )  ;
assign n12760 =  ( n12759 ) ^ ( n12660 )  ;
assign n12761 = ~ ( n12760 ) ;
assign n12762 =  ( n12736 ) | ( n12761 )  ;
assign n12763 = ~ ( n12762 ) ;
assign n12764 =  ( n12668 ) | ( n12763 )  ;
assign n12765 = ~ ( n12722 ) ;
assign n12766 =  ( n2426 ) ^ ( n2070 )  ;
assign n12767 =  ( n12766 ) ^ ( n1682 )  ;
assign n12768 =  ( n12767 ) ^ ( n1713 )  ;
assign n12769 =  ( n12768 ) ^ ( n1723 )  ;
assign n12770 =  ( n12769 ) ^ ( n1281 )  ;
assign n12771 =  ( n12770 ) ^ ( n1297 )  ;
assign n12772 =  ( n12771 ) ^ ( n1314 )  ;
assign n12773 =  ( n12772 ) ^ ( n1331 )  ;
assign n12774 =  ( n12773 ) ^ ( n1375 )  ;
assign n12775 =  ( n12774 ) ^ ( n12530 )  ;
assign n12776 =  ( n12775 ) ^ ( n7392 )  ;
assign n12777 =  ( n12776 ) ^ ( n7022 )  ;
assign n12778 =  ( n12777 ) ^ ( n6589 )  ;
assign n12779 =  ( n12778 ) ^ ( n6634 )  ;
assign n12780 = ~ ( n6640 ) ;
assign n12781 = ~ ( n6173 ) ;
assign n12782 =  ( n12780 ) | ( n12781 )  ;
assign n12783 =  ( n12779 ) ^ ( n12782 )  ;
assign n12784 =  ( n6030 ) | ( n6039 )  ;
assign n12785 =  ( n12784 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n12786 =  ( n12783 ) ^ ( n12785 )  ;
assign n12787 =  ( n5802 ) | ( n5811 )  ;
assign n12788 =  ( n12787 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12789 =  ( n12786 ) ^ ( n12788 )  ;
assign n12790 =  ( n5832 ) | ( n5841 )  ;
assign n12791 =  ( n12790 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12792 =  ( n12789 ) ^ ( n12791 )  ;
assign n12793 =  ( n5682 ) | ( n5691 )  ;
assign n12794 =  ( n12793 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12795 =  ( n12792 ) ^ ( n12794 )  ;
assign n12796 =  ( n5713 ) | ( n5722 )  ;
assign n12797 =  ( n12796 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12798 =  ( n12795 ) ^ ( n12797 )  ;
assign n12799 =  ( n12798 ) ^ ( n12660 )  ;
assign n12800 = ~ ( n12799 ) ;
assign n12801 =  ( n12765 ) | ( n12800 )  ;
assign n12802 = ~ ( n2727 ) ;
assign n12803 =  ( n12802 ) ^ ( n2388 )  ;
assign n12804 =  ( n12803 ) ^ ( n2038 )  ;
assign n12805 =  ( n12804 ) ^ ( n2052 )  ;
assign n12806 =  ( n12805 ) ^ ( n1632 )  ;
assign n12807 =  ( n12806 ) ^ ( n1642 )  ;
assign n12808 =  ( n1475 ) | ( n1484 )  ;
assign n12809 =  ( n12808 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n12810 = ~ ( n12809 ) ;
assign n12811 =  ( n12807 ) ^ ( n12810 )  ;
assign n12812 =  ( n12811 ) ^ ( n1656 )  ;
assign n12813 =  ( n12812 ) ^ ( n1663 )  ;
assign n12814 =  ( n12813 ) ^ ( n1670 )  ;
assign n12815 =  ( n12814 ) ^ ( n1677 )  ;
assign n12816 =  ( n12815 ) ^ ( n2422 )  ;
assign n12817 = ~ ( n3043 ) ;
assign n12818 =  ( n12817 ) | ( n3059 )  ;
assign n12819 = ~ ( n12818 ) ;
assign n12820 = ~ ( n3366 ) ;
assign n12821 = ~ ( n3392 ) ;
assign n12822 = ~ ( n3623 ) ;
assign n12823 =  ( n12821 ) | ( n12822 )  ;
assign n12824 =  ( n12823 ) | ( n3646 )  ;
assign n12825 = ~ ( n12824 ) ;
assign n12826 =  ( n12820 ) | ( n12825 )  ;
assign n12827 = ~ ( n4184 ) ;
assign n12828 =  ( n12826 ) | ( n12827 )  ;
assign n12829 = ~ ( n3392 ) ;
assign n12830 =  ( n12829 ) | ( n3672 )  ;
assign n12831 =  ( n12830 ) | ( n3985 )  ;
assign n12832 =  ( n12831 ) | ( n4253 )  ;
assign n12833 = ~ ( n11234 ) ;
assign n12834 =  ( n12832 ) | ( n12833 )  ;
assign n12835 = ~ ( n12834 ) ;
assign n12836 =  ( n12828 ) | ( n12835 )  ;
assign n12837 = ~ ( n3392 ) ;
assign n12838 =  ( n12837 ) | ( n3672 )  ;
assign n12839 =  ( n12838 ) | ( n3985 )  ;
assign n12840 =  ( n12839 ) | ( n4253 )  ;
assign n12841 =  ( n12840 ) | ( n4458 )  ;
assign n12842 =  ( n12841 ) | ( n4710 )  ;
assign n12843 = ~ ( n4763 ) ;
assign n12844 =  ( n12842 ) | ( n12843 )  ;
assign n12845 = ~ ( n4938 ) ;
assign n12846 =  ( n12844 ) | ( n12845 )  ;
assign n12847 =  ( n5041 ) | ( n5203 )  ;
assign n12848 =  ( n12847 ) | ( n5345 )  ;
assign n12849 =  ( n12848 ) | ( n11288 )  ;
assign n12850 = ~ ( n12849 ) ;
assign n12851 =  ( n12846 ) | ( n12850 )  ;
assign n12852 = ~ ( n12851 ) ;
assign n12853 =  ( n12836 ) | ( n12852 )  ;
assign n12854 = ~ ( n3392 ) ;
assign n12855 =  ( n12854 ) | ( n3672 )  ;
assign n12856 =  ( n12855 ) | ( n3985 )  ;
assign n12857 =  ( n12856 ) | ( n4253 )  ;
assign n12858 =  ( n12857 ) | ( n4458 )  ;
assign n12859 =  ( n12858 ) | ( n4710 )  ;
assign n12860 = ~ ( n4763 ) ;
assign n12861 =  ( n12859 ) | ( n12860 )  ;
assign n12862 = ~ ( n4938 ) ;
assign n12863 =  ( n12861 ) | ( n12862 )  ;
assign n12864 =  ( n12863 ) | ( n5063 )  ;
assign n12865 =  ( n12864 ) | ( n5224 )  ;
assign n12866 =  ( n12865 ) | ( n5265 )  ;
assign n12867 =  ( n5366 ) ^ ( n5161 )  ;
assign n12868 =  ( n12867 ) ^ ( n5171 )  ;
assign n12869 =  ( n12868 ) ^ ( n4960 )  ;
assign n12870 =  ( n12869 ) ^ ( n4976 )  ;
assign n12871 =  ( n12870 ) ^ ( n4996 )  ;
assign n12872 =  ( n12871 ) ^ ( n5236 )  ;
assign n12873 = ~ ( n12872 ) ;
assign n12874 =  ( n12866 ) | ( n12873 )  ;
assign n12875 =  ( n5452 ) ^ ( n5325 )  ;
assign n12876 =  ( n12875 ) ^ ( n5083 )  ;
assign n12877 =  ( n12876 ) ^ ( n5099 )  ;
assign n12878 =  ( n12877 ) ^ ( n5116 )  ;
assign n12879 =  ( n12878 ) ^ ( n5141 )  ;
assign n12880 =  ( n12879 ) ^ ( n5129 )  ;
assign n12881 = ~ ( n12880 ) ;
assign n12882 =  ( n12874 ) | ( n12881 )  ;
assign n12883 =  ( n5489 ) ^ ( n5433 )  ;
assign n12884 =  ( n12883 ) ^ ( n5285 )  ;
assign n12885 =  ( n12884 ) ^ ( n5301 )  ;
assign n12886 =  ( n12885 ) ^ ( n5321 )  ;
assign n12887 = ~ ( n12886 ) ;
assign n12888 =  ( n12882 ) | ( n12887 )  ;
assign n12889 = ~ ( n5547 ) ;
assign n12890 =  ( n12888 ) | ( n12889 )  ;
assign n12891 =  ( n5594 ) ^ ( n5515 )  ;
assign n12892 =  ( n12891 ) ^ ( n5531 )  ;
assign n12893 = ~ ( n12892 ) ;
assign n12894 =  ( n12890 ) | ( n12893 )  ;
assign n12895 =  ( n5568 ) ^ ( n5583 )  ;
assign n12896 =  ( n12895 ) ^ ( n5580 )  ;
assign n12897 = ~ ( n12896 ) ;
assign n12898 =  ( n12894 ) | ( n12897 )  ;
assign n12899 = ~ ( n5648 ) ;
assign n12900 =  ( n12898 ) | ( n12899 )  ;
assign n12901 = ~ ( n5657 ) ;
assign n12902 =  ( n12900 ) | ( n12901 )  ;
assign n12903 = ki[1:1] ;
assign n12904 = ~ ( n12903 ) ;
assign n12905 =  ( n12902 ) | ( n12904 )  ;
assign n12906 = ~ ( n12905 ) ;
assign n12907 =  ( n12853 ) | ( n12906 )  ;
assign n12908 = ~ ( n12907 ) ;
assign n12909 =  ( n3085 ) | ( n12908 )  ;
assign n12910 = ~ ( n12909 ) ;
assign n12911 =  ( n12819 ) | ( n12910 )  ;
assign n12912 =  ( n12816 ) ^ ( n12911 )  ;
assign n12913 = ~ ( n12912 ) ;
assign n12914 = ~ ( n7649 ) ;
assign n12915 =  ( n12914 ) | ( n7679 )  ;
assign n12916 = ~ ( n12915 ) ;
assign n12917 = ~ ( n7281 ) ;
assign n12918 =  ( n7287 ) | ( n7311 )  ;
assign n12919 = ~ ( n12918 ) ;
assign n12920 =  ( n12917 ) | ( n12919 )  ;
assign n12921 =  ( n12916 ) ^ ( n12920 )  ;
assign n12922 =  ( n12921 ) ^ ( n6970 )  ;
assign n12923 = ~ ( n6977 ) ;
assign n12924 = ~ ( n6982 ) ;
assign n12925 =  ( n12923 ) | ( n12924 )  ;
assign n12926 =  ( n12922 ) ^ ( n12925 )  ;
assign n12927 = ~ ( n6517 ) ;
assign n12928 =  ( n6524 ) | ( n6150 )  ;
assign n12929 = ~ ( n12928 ) ;
assign n12930 =  ( n12927 ) | ( n12929 )  ;
assign n12931 = ~ ( n6543 ) ;
assign n12932 =  ( n12930 ) | ( n12931 )  ;
assign n12933 =  ( n12926 ) ^ ( n12932 )  ;
assign n12934 = ~ ( n6553 ) ;
assign n12935 = ~ ( n6173 ) ;
assign n12936 =  ( n12934 ) | ( n12935 )  ;
assign n12937 =  ( n12933 ) ^ ( n12936 )  ;
assign n12938 =  ( n6483 ) | ( n6492 )  ;
assign n12939 =  ( n12938 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n12940 = ~ ( n12939 ) ;
assign n12941 =  ( n12937 ) ^ ( n12940 )  ;
assign n12942 =  ( n6030 ) | ( n6039 )  ;
assign n12943 =  ( n12942 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n12944 =  ( n12941 ) ^ ( n12943 )  ;
assign n12945 =  ( n5802 ) | ( n5811 )  ;
assign n12946 =  ( n12945 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n12947 =  ( n12944 ) ^ ( n12946 )  ;
assign n12948 =  ( n5832 ) | ( n5841 )  ;
assign n12949 =  ( n12948 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n12950 =  ( n12947 ) ^ ( n12949 )  ;
assign n12951 =  ( n5682 ) | ( n5691 )  ;
assign n12952 =  ( n12951 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n12953 =  ( n12950 ) ^ ( n12952 )  ;
assign n12954 =  ( n5713 ) | ( n5722 )  ;
assign n12955 =  ( n12954 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n12956 =  ( n12953 ) ^ ( n12955 )  ;
assign n12957 = ~ ( n8047 ) ;
assign n12958 =  ( n12957 ) | ( n8079 )  ;
assign n12959 = ~ ( n12958 ) ;
assign n12960 = ~ ( n8279 ) ;
assign n12961 = ~ ( n8321 ) ;
assign n12962 =  ( n12960 ) | ( n12961 )  ;
assign n12963 = ~ ( n8364 ) ;
assign n12964 =  ( n12962 ) | ( n12963 )  ;
assign n12965 = ~ ( n12964 ) ;
assign n12966 = ~ ( n8413 ) ;
assign n12967 = ~ ( n8625 ) ;
assign n12968 =  ( n12966 ) | ( n12967 )  ;
assign n12969 = ~ ( n8669 ) ;
assign n12970 =  ( n12968 ) | ( n12969 )  ;
assign n12971 = ~ ( n12970 ) ;
assign n12972 =  ( n12965 ) | ( n12971 )  ;
assign n12973 = ~ ( n8413 ) ;
assign n12974 = ~ ( n8717 ) ;
assign n12975 =  ( n12973 ) | ( n12974 )  ;
assign n12976 = ~ ( n9172 ) ;
assign n12977 =  ( n12975 ) | ( n12976 )  ;
assign n12978 = ~ ( n12977 ) ;
assign n12979 =  ( n12972 ) | ( n12978 )  ;
assign n12980 =  ( n12979 ) | ( n11446 )  ;
assign n12981 = ~ ( n8413 ) ;
assign n12982 = ~ ( n8717 ) ;
assign n12983 =  ( n12981 ) | ( n12982 )  ;
assign n12984 = ~ ( n9012 ) ;
assign n12985 =  ( n12983 ) | ( n12984 )  ;
assign n12986 = ~ ( n9252 ) ;
assign n12987 =  ( n12985 ) | ( n12986 )  ;
assign n12988 = ~ ( n9432 ) ;
assign n12989 =  ( n12987 ) | ( n12988 )  ;
assign n12990 = ~ ( n9649 ) ;
assign n12991 =  ( n12989 ) | ( n12990 )  ;
assign n12992 = ~ ( n9751 ) ;
assign n12993 =  ( n12991 ) | ( n12992 )  ;
assign n12994 = ~ ( n9909 ) ;
assign n12995 =  ( n12993 ) | ( n12994 )  ;
assign n12996 = ~ ( n10005 ) ;
assign n12997 = ~ ( n10042 ) ;
assign n12998 = ~ ( n10140 ) ;
assign n12999 =  ( n12997 ) | ( n12998 )  ;
assign n13000 =  ( n12999 ) | ( n10158 )  ;
assign n13001 =  ( n13000 ) | ( n10180 )  ;
assign n13002 = ~ ( n13001 ) ;
assign n13003 =  ( n12996 ) | ( n13002 )  ;
assign n13004 = ~ ( n10314 ) ;
assign n13005 =  ( n13003 ) | ( n13004 )  ;
assign n13006 =  ( n13005 ) | ( n11508 )  ;
assign n13007 = ~ ( n13006 ) ;
assign n13008 =  ( n12995 ) | ( n13007 )  ;
assign n13009 = ~ ( n13008 ) ;
assign n13010 =  ( n12980 ) | ( n13009 )  ;
assign n13011 = ~ ( n8413 ) ;
assign n13012 = ~ ( n8717 ) ;
assign n13013 =  ( n13011 ) | ( n13012 )  ;
assign n13014 = ~ ( n9012 ) ;
assign n13015 =  ( n13013 ) | ( n13014 )  ;
assign n13016 = ~ ( n9252 ) ;
assign n13017 =  ( n13015 ) | ( n13016 )  ;
assign n13018 = ~ ( n9432 ) ;
assign n13019 =  ( n13017 ) | ( n13018 )  ;
assign n13020 = ~ ( n9649 ) ;
assign n13021 =  ( n13019 ) | ( n13020 )  ;
assign n13022 = ~ ( n9751 ) ;
assign n13023 =  ( n13021 ) | ( n13022 )  ;
assign n13024 = ~ ( n9909 ) ;
assign n13025 =  ( n13023 ) | ( n13024 )  ;
assign n13026 = ~ ( n10042 ) ;
assign n13027 =  ( n13025 ) | ( n13026 )  ;
assign n13028 = ~ ( n10208 ) ;
assign n13029 =  ( n13027 ) | ( n13028 )  ;
assign n13030 =  ( n13029 ) | ( n10274 )  ;
assign n13031 = ~ ( n10358 ) ;
assign n13032 =  ( n13030 ) | ( n13031 )  ;
assign n13033 = ~ ( n10430 ) ;
assign n13034 =  ( n13032 ) | ( n13033 )  ;
assign n13035 =  ( n13034 ) | ( n10467 )  ;
assign n13036 =  ( n13035 ) | ( n10489 )  ;
assign n13037 =  ( n13036 ) | ( n10550 )  ;
assign n13038 =  ( n7455 ) ^ ( n10522 )  ;
assign n13039 =  ( n13038 ) ^ ( n10519 )  ;
assign n13040 = ~ ( n13039 ) ;
assign n13041 =  ( n13037 ) | ( n13040 )  ;
assign n13042 = ~ ( n7455 ) ;
assign n13043 =  ( n13041 ) | ( n13042 )  ;
assign n13044 = ~ ( n10564 ) ;
assign n13045 =  ( n13043 ) | ( n13044 )  ;
assign n13046 = kd[1:1] ;
assign n13047 = ~ ( n13046 ) ;
assign n13048 =  ( n13045 ) | ( n13047 )  ;
assign n13049 = ~ ( n13048 ) ;
assign n13050 =  ( n13010 ) | ( n13049 )  ;
assign n13051 = ~ ( n13050 ) ;
assign n13052 =  ( n8121 ) | ( n13051 )  ;
assign n13053 = ~ ( n13052 ) ;
assign n13054 =  ( n12959 ) | ( n13053 )  ;
assign n13055 =  ( n12956 ) ^ ( n13054 )  ;
assign n13056 = ~ ( n13055 ) ;
assign n13057 =  ( n12913 ) | ( n13056 )  ;
assign n13058 = ~ ( n13057 ) ;
assign n13059 = ~ ( n2727 ) ;
assign n13060 =  ( n13059 ) ^ ( n2388 )  ;
assign n13061 =  ( n13060 ) ^ ( n2038 )  ;
assign n13062 =  ( n13061 ) ^ ( n2052 )  ;
assign n13063 =  ( n13062 ) ^ ( n1632 )  ;
assign n13064 =  ( n13063 ) ^ ( n1642 )  ;
assign n13065 =  ( n1475 ) | ( n1484 )  ;
assign n13066 =  ( n13065 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n13067 = ~ ( n13066 ) ;
assign n13068 =  ( n13064 ) ^ ( n13067 )  ;
assign n13069 =  ( n13068 ) ^ ( n1656 )  ;
assign n13070 =  ( n13069 ) ^ ( n1663 )  ;
assign n13071 =  ( n13070 ) ^ ( n1670 )  ;
assign n13072 =  ( n13071 ) ^ ( n1677 )  ;
assign n13073 =  ( n13072 ) ^ ( n2422 )  ;
assign n13074 =  ( n13073 ) ^ ( n12911 )  ;
assign n13075 = ~ ( n7649 ) ;
assign n13076 =  ( n13075 ) | ( n7679 )  ;
assign n13077 = ~ ( n13076 ) ;
assign n13078 =  ( n13074 ) ^ ( n13077 )  ;
assign n13079 = ~ ( n7281 ) ;
assign n13080 =  ( n7287 ) | ( n7311 )  ;
assign n13081 = ~ ( n13080 ) ;
assign n13082 =  ( n13079 ) | ( n13081 )  ;
assign n13083 =  ( n13078 ) ^ ( n13082 )  ;
assign n13084 =  ( n13083 ) ^ ( n6970 )  ;
assign n13085 = ~ ( n6977 ) ;
assign n13086 = ~ ( n6982 ) ;
assign n13087 =  ( n13085 ) | ( n13086 )  ;
assign n13088 =  ( n13084 ) ^ ( n13087 )  ;
assign n13089 = ~ ( n6517 ) ;
assign n13090 =  ( n6524 ) | ( n6150 )  ;
assign n13091 = ~ ( n13090 ) ;
assign n13092 =  ( n13089 ) | ( n13091 )  ;
assign n13093 = ~ ( n6543 ) ;
assign n13094 =  ( n13092 ) | ( n13093 )  ;
assign n13095 =  ( n13088 ) ^ ( n13094 )  ;
assign n13096 = ~ ( n6553 ) ;
assign n13097 = ~ ( n6173 ) ;
assign n13098 =  ( n13096 ) | ( n13097 )  ;
assign n13099 =  ( n13095 ) ^ ( n13098 )  ;
assign n13100 =  ( n6483 ) | ( n6492 )  ;
assign n13101 =  ( n13100 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13102 = ~ ( n13101 ) ;
assign n13103 =  ( n13099 ) ^ ( n13102 )  ;
assign n13104 =  ( n6030 ) | ( n6039 )  ;
assign n13105 =  ( n13104 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13106 =  ( n13103 ) ^ ( n13105 )  ;
assign n13107 =  ( n5802 ) | ( n5811 )  ;
assign n13108 =  ( n13107 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13109 =  ( n13106 ) ^ ( n13108 )  ;
assign n13110 =  ( n5832 ) | ( n5841 )  ;
assign n13111 =  ( n13110 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13112 =  ( n13109 ) ^ ( n13111 )  ;
assign n13113 =  ( n5682 ) | ( n5691 )  ;
assign n13114 =  ( n13113 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13115 =  ( n13112 ) ^ ( n13114 )  ;
assign n13116 =  ( n5713 ) | ( n5722 )  ;
assign n13117 =  ( n13116 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13118 =  ( n13115 ) ^ ( n13117 )  ;
assign n13119 =  ( n13118 ) ^ ( n13054 )  ;
assign n13120 = ~ ( n13119 ) ;
assign n13121 =  ( bv_1_1_n5 ) ^ ( n3043 )  ;
assign n13122 = ~ ( n2692 ) ;
assign n13123 =  ( n2675 ) | ( n13122 )  ;
assign n13124 =  ( n13121 ) ^ ( n13123 )  ;
assign n13125 =  ( n13124 ) ^ ( n2361 )  ;
assign n13126 =  ( n13125 ) ^ ( n2371 )  ;
assign n13127 =  ( n13126 ) ^ ( n1952 )  ;
assign n13128 =  ( n13127 ) ^ ( n1963 )  ;
assign n13129 =  ( n13128 ) ^ ( n1513 )  ;
assign n13130 =  ( n13129 ) ^ ( n1538 )  ;
assign n13131 =  ( n13130 ) ^ ( n1564 )  ;
assign n13132 =  ( n13131 ) ^ ( n1590 )  ;
assign n13133 =  ( n13132 ) ^ ( n1628 )  ;
assign n13134 =  ( n13133 ) ^ ( n2016 )  ;
assign n13135 =  ( n13134 ) ^ ( n12907 )  ;
assign n13136 = ~ ( n13135 ) ;
assign n13137 =  ( n13120 ) | ( n13136 )  ;
assign n13138 =  ( bv_1_1_n5 ) ^ ( n8047 )  ;
assign n13139 =  ( n13138 ) ^ ( n7649 )  ;
assign n13140 =  ( n13139 ) ^ ( n7265 )  ;
assign n13141 = ~ ( n7271 ) ;
assign n13142 = ~ ( n7277 ) ;
assign n13143 =  ( n13141 ) | ( n13142 )  ;
assign n13144 =  ( n13140 ) ^ ( n13143 )  ;
assign n13145 =  ( n13144 ) ^ ( n6888 )  ;
assign n13146 = ~ ( n6895 ) ;
assign n13147 = ~ ( n6366 ) ;
assign n13148 =  ( n13146 ) | ( n13147 )  ;
assign n13149 =  ( n13145 ) ^ ( n13148 )  ;
assign n13150 =  ( n6483 ) | ( n6492 )  ;
assign n13151 =  ( n13150 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13152 =  ( n13149 ) ^ ( n13151 )  ;
assign n13153 =  ( n6030 ) | ( n6039 )  ;
assign n13154 =  ( n13153 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13155 =  ( n13152 ) ^ ( n13154 )  ;
assign n13156 =  ( n5802 ) | ( n5811 )  ;
assign n13157 =  ( n13156 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13158 =  ( n13155 ) ^ ( n13157 )  ;
assign n13159 =  ( n5832 ) | ( n5841 )  ;
assign n13160 =  ( n13159 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13161 =  ( n13158 ) ^ ( n13160 )  ;
assign n13162 =  ( n5682 ) | ( n5691 )  ;
assign n13163 =  ( n13162 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13164 =  ( n13161 ) ^ ( n13163 )  ;
assign n13165 =  ( n5713 ) | ( n5722 )  ;
assign n13166 =  ( n13165 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13167 =  ( n13164 ) ^ ( n13166 )  ;
assign n13168 =  ( n13167 ) ^ ( n13050 )  ;
assign n13169 = ~ ( n13168 ) ;
assign n13170 =  ( n13137 ) | ( n13169 )  ;
assign n13171 = ~ ( n13170 ) ;
assign n13172 =  ( n13058 ) | ( n13171 )  ;
assign n13173 = ~ ( n13172 ) ;
assign n13174 =  ( n12801 ) | ( n13173 )  ;
assign n13175 = ~ ( n13174 ) ;
assign n13176 =  ( n12764 ) | ( n13175 )  ;
assign n13177 = ~ ( n12722 ) ;
assign n13178 =  ( n13177 ) | ( n12800 )  ;
assign n13179 = ~ ( n13119 ) ;
assign n13180 =  ( n13178 ) | ( n13179 )  ;
assign n13181 = ~ ( n2692 ) ;
assign n13182 =  ( n2675 ) | ( n13181 )  ;
assign n13183 =  ( n3043 ) ^ ( n13182 )  ;
assign n13184 =  ( n13183 ) ^ ( n2361 )  ;
assign n13185 =  ( n13184 ) ^ ( n2371 )  ;
assign n13186 =  ( n13185 ) ^ ( n1952 )  ;
assign n13187 =  ( n13186 ) ^ ( n1963 )  ;
assign n13188 =  ( n13187 ) ^ ( n1513 )  ;
assign n13189 =  ( n13188 ) ^ ( n1538 )  ;
assign n13190 =  ( n13189 ) ^ ( n1564 )  ;
assign n13191 =  ( n13190 ) ^ ( n1590 )  ;
assign n13192 =  ( n13191 ) ^ ( n1628 )  ;
assign n13193 =  ( n13192 ) ^ ( n2016 )  ;
assign n13194 =  ( n13193 ) ^ ( n12907 )  ;
assign n13195 =  ( n13194 ) ^ ( n8047 )  ;
assign n13196 =  ( n13195 ) ^ ( n7649 )  ;
assign n13197 =  ( n13196 ) ^ ( n7265 )  ;
assign n13198 = ~ ( n7271 ) ;
assign n13199 = ~ ( n7277 ) ;
assign n13200 =  ( n13198 ) | ( n13199 )  ;
assign n13201 =  ( n13197 ) ^ ( n13200 )  ;
assign n13202 =  ( n13201 ) ^ ( n6888 )  ;
assign n13203 = ~ ( n6895 ) ;
assign n13204 = ~ ( n6366 ) ;
assign n13205 =  ( n13203 ) | ( n13204 )  ;
assign n13206 =  ( n13202 ) ^ ( n13205 )  ;
assign n13207 =  ( n6483 ) | ( n6492 )  ;
assign n13208 =  ( n13207 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13209 =  ( n13206 ) ^ ( n13208 )  ;
assign n13210 =  ( n6030 ) | ( n6039 )  ;
assign n13211 =  ( n13210 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13212 =  ( n13209 ) ^ ( n13211 )  ;
assign n13213 =  ( n5802 ) | ( n5811 )  ;
assign n13214 =  ( n13213 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13215 =  ( n13212 ) ^ ( n13214 )  ;
assign n13216 =  ( n5832 ) | ( n5841 )  ;
assign n13217 =  ( n13216 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13218 =  ( n13215 ) ^ ( n13217 )  ;
assign n13219 =  ( n5682 ) | ( n5691 )  ;
assign n13220 =  ( n13219 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13221 =  ( n13218 ) ^ ( n13220 )  ;
assign n13222 =  ( n5713 ) | ( n5722 )  ;
assign n13223 =  ( n13222 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13224 =  ( n13221 ) ^ ( n13223 )  ;
assign n13225 =  ( n13224 ) ^ ( n13050 )  ;
assign n13226 = ~ ( n13225 ) ;
assign n13227 =  ( n13180 ) | ( n13226 )  ;
assign n13228 = ~ ( n3371 ) ;
assign n13229 = ~ ( n2973 ) ;
assign n13230 =  ( n13229 ) | ( n2994 )  ;
assign n13231 =  ( n13228 ) ^ ( n13230 )  ;
assign n13232 =  ( n2633 ) | ( n2643 )  ;
assign n13233 =  ( n13232 ) | ( n2657 )  ;
assign n13234 =  ( n13231 ) ^ ( n13233 )  ;
assign n13235 =  ( n13234 ) ^ ( n2672 )  ;
assign n13236 =  ( n13235 ) ^ ( n2227 )  ;
assign n13237 =  ( n13236 ) ^ ( n2237 )  ;
assign n13238 =  ( n13237 ) ^ ( n2314 )  ;
assign n13239 =  ( n1838 ) | ( n1847 )  ;
assign n13240 =  ( n13239 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n13241 = ~ ( n13240 ) ;
assign n13242 =  ( n13238 ) ^ ( n13241 )  ;
assign n13243 =  ( n13242 ) ^ ( n1879 )  ;
assign n13244 =  ( n13243 ) ^ ( n1896 )  ;
assign n13245 =  ( n13244 ) ^ ( n1913 )  ;
assign n13246 =  ( n13245 ) ^ ( n1948 )  ;
assign n13247 =  ( n13246 ) ^ ( n2357 )  ;
assign n13248 =  ( n13247 ) ^ ( n3039 )  ;
assign n13249 = ~ ( n3623 ) ;
assign n13250 =  ( n13249 ) | ( n3646 )  ;
assign n13251 = ~ ( n13250 ) ;
assign n13252 = ~ ( n3958 ) ;
assign n13253 =  ( n13252 ) | ( n4181 )  ;
assign n13254 = ~ ( n10705 ) ;
assign n13255 =  ( n13253 ) | ( n13254 )  ;
assign n13256 =  ( n3985 ) | ( n4253 )  ;
assign n13257 =  ( n13256 ) | ( n4458 )  ;
assign n13258 =  ( n13257 ) | ( n4710 )  ;
assign n13259 = ~ ( n11703 ) ;
assign n13260 =  ( n13258 ) | ( n13259 )  ;
assign n13261 = ~ ( n13260 ) ;
assign n13262 =  ( n13255 ) | ( n13261 )  ;
assign n13263 =  ( n3985 ) | ( n4253 )  ;
assign n13264 =  ( n13263 ) | ( n4458 )  ;
assign n13265 =  ( n13264 ) | ( n4710 )  ;
assign n13266 = ~ ( n4763 ) ;
assign n13267 =  ( n13265 ) | ( n13266 )  ;
assign n13268 = ~ ( n4938 ) ;
assign n13269 =  ( n13267 ) | ( n13268 )  ;
assign n13270 =  ( n13269 ) | ( n5063 )  ;
assign n13271 =  ( n13270 ) | ( n5224 )  ;
assign n13272 =  ( n5248 ) | ( n5341 )  ;
assign n13273 =  ( n13272 ) | ( n10785 )  ;
assign n13274 =  ( n13273 ) | ( n11760 )  ;
assign n13275 = ~ ( n13274 ) ;
assign n13276 =  ( n13271 ) | ( n13275 )  ;
assign n13277 = ~ ( n13276 ) ;
assign n13278 =  ( n13262 ) | ( n13277 )  ;
assign n13279 =  ( n3985 ) | ( n4253 )  ;
assign n13280 =  ( n13279 ) | ( n4458 )  ;
assign n13281 =  ( n13280 ) | ( n4710 )  ;
assign n13282 = ~ ( n4763 ) ;
assign n13283 =  ( n13281 ) | ( n13282 )  ;
assign n13284 = ~ ( n4938 ) ;
assign n13285 =  ( n13283 ) | ( n13284 )  ;
assign n13286 =  ( n13285 ) | ( n5063 )  ;
assign n13287 =  ( n13286 ) | ( n5224 )  ;
assign n13288 =  ( n13287 ) | ( n5265 )  ;
assign n13289 =  ( n5366 ) ^ ( n5161 )  ;
assign n13290 =  ( n13289 ) ^ ( n5171 )  ;
assign n13291 =  ( n13290 ) ^ ( n4960 )  ;
assign n13292 =  ( n13291 ) ^ ( n4976 )  ;
assign n13293 =  ( n13292 ) ^ ( n4996 )  ;
assign n13294 =  ( n13293 ) ^ ( n5236 )  ;
assign n13295 = ~ ( n13294 ) ;
assign n13296 =  ( n13288 ) | ( n13295 )  ;
assign n13297 =  ( n5452 ) ^ ( n5325 )  ;
assign n13298 =  ( n13297 ) ^ ( n5083 )  ;
assign n13299 =  ( n13298 ) ^ ( n5099 )  ;
assign n13300 =  ( n13299 ) ^ ( n5116 )  ;
assign n13301 =  ( n13300 ) ^ ( n5141 )  ;
assign n13302 =  ( n13301 ) ^ ( n5129 )  ;
assign n13303 = ~ ( n13302 ) ;
assign n13304 =  ( n13296 ) | ( n13303 )  ;
assign n13305 =  ( n5489 ) ^ ( n5433 )  ;
assign n13306 =  ( n13305 ) ^ ( n5285 )  ;
assign n13307 =  ( n13306 ) ^ ( n5301 )  ;
assign n13308 =  ( n13307 ) ^ ( n5321 )  ;
assign n13309 = ~ ( n13308 ) ;
assign n13310 =  ( n13304 ) | ( n13309 )  ;
assign n13311 = ~ ( n5547 ) ;
assign n13312 =  ( n13310 ) | ( n13311 )  ;
assign n13313 =  ( n5594 ) ^ ( n5515 )  ;
assign n13314 =  ( n13313 ) ^ ( n5531 )  ;
assign n13315 = ~ ( n13314 ) ;
assign n13316 =  ( n13312 ) | ( n13315 )  ;
assign n13317 =  ( n5568 ) ^ ( n5583 )  ;
assign n13318 =  ( n13317 ) ^ ( n5580 )  ;
assign n13319 = ~ ( n13318 ) ;
assign n13320 =  ( n13316 ) | ( n13319 )  ;
assign n13321 = ~ ( n5648 ) ;
assign n13322 =  ( n13320 ) | ( n13321 )  ;
assign n13323 = ~ ( n5657 ) ;
assign n13324 =  ( n13322 ) | ( n13323 )  ;
assign n13325 = ki[1:1] ;
assign n13326 = ~ ( n13325 ) ;
assign n13327 =  ( n13324 ) | ( n13326 )  ;
assign n13328 = ~ ( n13327 ) ;
assign n13329 =  ( n13278 ) | ( n13328 )  ;
assign n13330 = ~ ( n13329 ) ;
assign n13331 =  ( n3672 ) | ( n13330 )  ;
assign n13332 = ~ ( n13331 ) ;
assign n13333 =  ( n13251 ) | ( n13332 )  ;
assign n13334 =  ( n13248 ) ^ ( n13333 )  ;
assign n13335 = ~ ( n13334 ) ;
assign n13336 = ~ ( n8279 ) ;
assign n13337 = ~ ( n8321 ) ;
assign n13338 =  ( n13336 ) | ( n13337 )  ;
assign n13339 = ~ ( n13338 ) ;
assign n13340 =  ( n13339 ) ^ ( n7961 )  ;
assign n13341 =  ( n13340 ) ^ ( n7591 )  ;
assign n13342 = ~ ( n7597 ) ;
assign n13343 = ~ ( n7603 ) ;
assign n13344 =  ( n13342 ) | ( n13343 )  ;
assign n13345 =  ( n13341 ) ^ ( n13344 )  ;
assign n13346 = ~ ( n7133 ) ;
assign n13347 =  ( n7140 ) | ( n6337 )  ;
assign n13348 = ~ ( n13347 ) ;
assign n13349 =  ( n13346 ) | ( n13348 )  ;
assign n13350 = ~ ( n7159 ) ;
assign n13351 =  ( n13349 ) | ( n13350 )  ;
assign n13352 =  ( n13345 ) ^ ( n13351 )  ;
assign n13353 = ~ ( n7169 ) ;
assign n13354 = ~ ( n6366 ) ;
assign n13355 =  ( n13353 ) | ( n13354 )  ;
assign n13356 =  ( n13352 ) ^ ( n13355 )  ;
assign n13357 = ~ ( n5736 ) ;
assign n13358 =  ( n13357 ) | ( n5742 )  ;
assign n13359 =  ( n13356 ) ^ ( n13358 )  ;
assign n13360 =  ( n6825 ) | ( n6834 )  ;
assign n13361 =  ( n13360 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n13362 = ~ ( n13361 ) ;
assign n13363 =  ( n13359 ) ^ ( n13362 )  ;
assign n13364 =  ( n6483 ) | ( n6492 )  ;
assign n13365 =  ( n13364 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13366 =  ( n13363 ) ^ ( n13365 )  ;
assign n13367 =  ( n6030 ) | ( n6039 )  ;
assign n13368 =  ( n13367 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13369 =  ( n13366 ) ^ ( n13368 )  ;
assign n13370 =  ( n5802 ) | ( n5811 )  ;
assign n13371 =  ( n13370 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13372 =  ( n13369 ) ^ ( n13371 )  ;
assign n13373 =  ( n5832 ) | ( n5841 )  ;
assign n13374 =  ( n13373 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13375 =  ( n13372 ) ^ ( n13374 )  ;
assign n13376 =  ( n5682 ) | ( n5691 )  ;
assign n13377 =  ( n13376 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13378 =  ( n13375 ) ^ ( n13377 )  ;
assign n13379 =  ( n5713 ) | ( n5722 )  ;
assign n13380 =  ( n13379 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13381 =  ( n13378 ) ^ ( n13380 )  ;
assign n13382 = ~ ( n8625 ) ;
assign n13383 = ~ ( n8669 ) ;
assign n13384 =  ( n13382 ) | ( n13383 )  ;
assign n13385 = ~ ( n13384 ) ;
assign n13386 = ~ ( n8717 ) ;
assign n13387 = ~ ( n8880 ) ;
assign n13388 = ~ ( n8920 ) ;
assign n13389 =  ( n13387 ) | ( n13388 )  ;
assign n13390 = ~ ( n8963 ) ;
assign n13391 =  ( n13389 ) | ( n13390 )  ;
assign n13392 = ~ ( n13391 ) ;
assign n13393 =  ( n13392 ) | ( n9171 )  ;
assign n13394 = ~ ( n9012 ) ;
assign n13395 = ~ ( n9252 ) ;
assign n13396 =  ( n13394 ) | ( n13395 )  ;
assign n13397 = ~ ( n10966 ) ;
assign n13398 =  ( n13396 ) | ( n13397 )  ;
assign n13399 = ~ ( n13398 ) ;
assign n13400 =  ( n13393 ) | ( n13399 )  ;
assign n13401 =  ( n13400 ) | ( n11921 )  ;
assign n13402 = ~ ( n9012 ) ;
assign n13403 = ~ ( n9252 ) ;
assign n13404 =  ( n13402 ) | ( n13403 )  ;
assign n13405 = ~ ( n9432 ) ;
assign n13406 =  ( n13404 ) | ( n13405 )  ;
assign n13407 = ~ ( n9649 ) ;
assign n13408 =  ( n13406 ) | ( n13407 )  ;
assign n13409 = ~ ( n9751 ) ;
assign n13410 =  ( n13408 ) | ( n13409 )  ;
assign n13411 = ~ ( n9909 ) ;
assign n13412 =  ( n13410 ) | ( n13411 )  ;
assign n13413 = ~ ( n10042 ) ;
assign n13414 =  ( n13412 ) | ( n13413 )  ;
assign n13415 = ~ ( n10208 ) ;
assign n13416 =  ( n13414 ) | ( n13415 )  ;
assign n13417 = ~ ( n10249 ) ;
assign n13418 = ~ ( n10310 ) ;
assign n13419 =  ( n13417 ) | ( n13418 )  ;
assign n13420 = ~ ( n10358 ) ;
assign n13421 =  ( n10274 ) | ( n13420 )  ;
assign n13422 = ~ ( n11045 ) ;
assign n13423 =  ( n13421 ) | ( n13422 )  ;
assign n13424 = ~ ( n13423 ) ;
assign n13425 =  ( n13419 ) | ( n13424 )  ;
assign n13426 =  ( n13425 ) | ( n11971 )  ;
assign n13427 = ~ ( n13426 ) ;
assign n13428 =  ( n13416 ) | ( n13427 )  ;
assign n13429 = ~ ( n13428 ) ;
assign n13430 =  ( n13401 ) | ( n13429 )  ;
assign n13431 = ~ ( n9012 ) ;
assign n13432 = ~ ( n9252 ) ;
assign n13433 =  ( n13431 ) | ( n13432 )  ;
assign n13434 = ~ ( n9432 ) ;
assign n13435 =  ( n13433 ) | ( n13434 )  ;
assign n13436 = ~ ( n9649 ) ;
assign n13437 =  ( n13435 ) | ( n13436 )  ;
assign n13438 = ~ ( n9751 ) ;
assign n13439 =  ( n13437 ) | ( n13438 )  ;
assign n13440 = ~ ( n9909 ) ;
assign n13441 =  ( n13439 ) | ( n13440 )  ;
assign n13442 = ~ ( n10042 ) ;
assign n13443 =  ( n13441 ) | ( n13442 )  ;
assign n13444 = ~ ( n10208 ) ;
assign n13445 =  ( n13443 ) | ( n13444 )  ;
assign n13446 =  ( n13445 ) | ( n10274 )  ;
assign n13447 = ~ ( n10358 ) ;
assign n13448 =  ( n13446 ) | ( n13447 )  ;
assign n13449 = ~ ( n10430 ) ;
assign n13450 =  ( n13448 ) | ( n13449 )  ;
assign n13451 =  ( n13450 ) | ( n10467 )  ;
assign n13452 =  ( n13451 ) | ( n10489 )  ;
assign n13453 =  ( n13452 ) | ( n10550 )  ;
assign n13454 =  ( n7455 ) ^ ( n10522 )  ;
assign n13455 =  ( n13454 ) ^ ( n10519 )  ;
assign n13456 = ~ ( n13455 ) ;
assign n13457 =  ( n13453 ) | ( n13456 )  ;
assign n13458 = ~ ( n7455 ) ;
assign n13459 =  ( n13457 ) | ( n13458 )  ;
assign n13460 = ~ ( n10564 ) ;
assign n13461 =  ( n13459 ) | ( n13460 )  ;
assign n13462 = kd[1:1] ;
assign n13463 = ~ ( n13462 ) ;
assign n13464 =  ( n13461 ) | ( n13463 )  ;
assign n13465 = ~ ( n13464 ) ;
assign n13466 =  ( n13430 ) | ( n13465 )  ;
assign n13467 = ~ ( n13466 ) ;
assign n13468 =  ( n13386 ) | ( n13467 )  ;
assign n13469 = ~ ( n13468 ) ;
assign n13470 =  ( n13385 ) | ( n13469 )  ;
assign n13471 =  ( n13381 ) ^ ( n13470 )  ;
assign n13472 = ~ ( n13471 ) ;
assign n13473 =  ( n13335 ) | ( n13472 )  ;
assign n13474 = ~ ( n13473 ) ;
assign n13475 = ~ ( n3371 ) ;
assign n13476 = ~ ( n2973 ) ;
assign n13477 =  ( n13476 ) | ( n2994 )  ;
assign n13478 =  ( n13475 ) ^ ( n13477 )  ;
assign n13479 =  ( n2633 ) | ( n2643 )  ;
assign n13480 =  ( n13479 ) | ( n2657 )  ;
assign n13481 =  ( n13478 ) ^ ( n13480 )  ;
assign n13482 =  ( n13481 ) ^ ( n2672 )  ;
assign n13483 =  ( n13482 ) ^ ( n2227 )  ;
assign n13484 =  ( n13483 ) ^ ( n2237 )  ;
assign n13485 =  ( n13484 ) ^ ( n2314 )  ;
assign n13486 =  ( n1838 ) | ( n1847 )  ;
assign n13487 =  ( n13486 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n13488 = ~ ( n13487 ) ;
assign n13489 =  ( n13485 ) ^ ( n13488 )  ;
assign n13490 =  ( n13489 ) ^ ( n1879 )  ;
assign n13491 =  ( n13490 ) ^ ( n1896 )  ;
assign n13492 =  ( n13491 ) ^ ( n1913 )  ;
assign n13493 =  ( n13492 ) ^ ( n1948 )  ;
assign n13494 =  ( n13493 ) ^ ( n2357 )  ;
assign n13495 =  ( n13494 ) ^ ( n3039 )  ;
assign n13496 =  ( n13495 ) ^ ( n13333 )  ;
assign n13497 = ~ ( n8279 ) ;
assign n13498 = ~ ( n8321 ) ;
assign n13499 =  ( n13497 ) | ( n13498 )  ;
assign n13500 = ~ ( n13499 ) ;
assign n13501 =  ( n13496 ) ^ ( n13500 )  ;
assign n13502 =  ( n13501 ) ^ ( n7961 )  ;
assign n13503 =  ( n13502 ) ^ ( n7591 )  ;
assign n13504 = ~ ( n7597 ) ;
assign n13505 = ~ ( n7603 ) ;
assign n13506 =  ( n13504 ) | ( n13505 )  ;
assign n13507 =  ( n13503 ) ^ ( n13506 )  ;
assign n13508 = ~ ( n7133 ) ;
assign n13509 =  ( n7140 ) | ( n6337 )  ;
assign n13510 = ~ ( n13509 ) ;
assign n13511 =  ( n13508 ) | ( n13510 )  ;
assign n13512 = ~ ( n7159 ) ;
assign n13513 =  ( n13511 ) | ( n13512 )  ;
assign n13514 =  ( n13507 ) ^ ( n13513 )  ;
assign n13515 = ~ ( n7169 ) ;
assign n13516 = ~ ( n6366 ) ;
assign n13517 =  ( n13515 ) | ( n13516 )  ;
assign n13518 =  ( n13514 ) ^ ( n13517 )  ;
assign n13519 = ~ ( n5736 ) ;
assign n13520 =  ( n13519 ) | ( n5742 )  ;
assign n13521 =  ( n13518 ) ^ ( n13520 )  ;
assign n13522 =  ( n6825 ) | ( n6834 )  ;
assign n13523 =  ( n13522 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n13524 = ~ ( n13523 ) ;
assign n13525 =  ( n13521 ) ^ ( n13524 )  ;
assign n13526 =  ( n6483 ) | ( n6492 )  ;
assign n13527 =  ( n13526 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13528 =  ( n13525 ) ^ ( n13527 )  ;
assign n13529 =  ( n6030 ) | ( n6039 )  ;
assign n13530 =  ( n13529 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13531 =  ( n13528 ) ^ ( n13530 )  ;
assign n13532 =  ( n5802 ) | ( n5811 )  ;
assign n13533 =  ( n13532 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13534 =  ( n13531 ) ^ ( n13533 )  ;
assign n13535 =  ( n5832 ) | ( n5841 )  ;
assign n13536 =  ( n13535 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13537 =  ( n13534 ) ^ ( n13536 )  ;
assign n13538 =  ( n5682 ) | ( n5691 )  ;
assign n13539 =  ( n13538 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13540 =  ( n13537 ) ^ ( n13539 )  ;
assign n13541 =  ( n5713 ) | ( n5722 )  ;
assign n13542 =  ( n13541 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13543 =  ( n13540 ) ^ ( n13542 )  ;
assign n13544 =  ( n13543 ) ^ ( n13470 )  ;
assign n13545 = ~ ( n13544 ) ;
assign n13546 =  ( bv_1_1_n5 ) ^ ( n3623 )  ;
assign n13547 = ~ ( n3323 ) ;
assign n13548 =  ( n3306 ) | ( n13547 )  ;
assign n13549 =  ( n13546 ) ^ ( n13548 )  ;
assign n13550 = ~ ( n2928 ) ;
assign n13551 = ~ ( n2939 ) ;
assign n13552 =  ( n13550 ) | ( n13551 )  ;
assign n13553 = ~ ( n2954 ) ;
assign n13554 =  ( n13552 ) | ( n13553 )  ;
assign n13555 =  ( n13549 ) ^ ( n13554 )  ;
assign n13556 =  ( n13555 ) ^ ( n2971 )  ;
assign n13557 =  ( n13556 ) ^ ( n2552 )  ;
assign n13558 =  ( n13557 ) ^ ( n2561 )  ;
assign n13559 =  ( n13558 ) ^ ( n2624 )  ;
assign n13560 =  ( n13559 ) ^ ( n2144 )  ;
assign n13561 =  ( n13560 ) ^ ( n2160 )  ;
assign n13562 =  ( n13561 ) ^ ( n2177 )  ;
assign n13563 =  ( n13562 ) ^ ( n2194 )  ;
assign n13564 =  ( n13563 ) ^ ( n2223 )  ;
assign n13565 =  ( n13564 ) ^ ( n2263 )  ;
assign n13566 =  ( n13565 ) ^ ( n2309 )  ;
assign n13567 =  ( n13566 ) ^ ( n13329 )  ;
assign n13568 = ~ ( n13567 ) ;
assign n13569 =  ( n13545 ) | ( n13568 )  ;
assign n13570 =  ( bv_1_1_n5 ) ^ ( n8625 )  ;
assign n13571 =  ( n13570 ) ^ ( n8279 )  ;
assign n13572 =  ( n13571 ) ^ ( n7899 )  ;
assign n13573 = ~ ( n7905 ) ;
assign n13574 = ~ ( n7911 ) ;
assign n13575 =  ( n13573 ) | ( n13574 )  ;
assign n13576 =  ( n13572 ) ^ ( n13575 )  ;
assign n13577 = ~ ( n7467 ) ;
assign n13578 =  ( n7473 ) | ( n6524 )  ;
assign n13579 = ~ ( n13578 ) ;
assign n13580 =  ( n13577 ) | ( n13579 )  ;
assign n13581 = ~ ( n7491 ) ;
assign n13582 =  ( n13580 ) | ( n13581 )  ;
assign n13583 =  ( n13576 ) ^ ( n13582 )  ;
assign n13584 = ~ ( n7498 ) ;
assign n13585 = ~ ( n6553 ) ;
assign n13586 =  ( n13584 ) | ( n13585 )  ;
assign n13587 =  ( n13583 ) ^ ( n13586 )  ;
assign n13588 = ~ ( n5902 ) ;
assign n13589 = ~ ( n5913 ) ;
assign n13590 =  ( n13588 ) | ( n13589 )  ;
assign n13591 =  ( n13587 ) ^ ( n13590 )  ;
assign n13592 =  ( n6825 ) | ( n6834 )  ;
assign n13593 =  ( n13592 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n13594 =  ( n13591 ) ^ ( n13593 )  ;
assign n13595 =  ( n6483 ) | ( n6492 )  ;
assign n13596 =  ( n13595 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13597 =  ( n13594 ) ^ ( n13596 )  ;
assign n13598 =  ( n6030 ) | ( n6039 )  ;
assign n13599 =  ( n13598 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13600 =  ( n13597 ) ^ ( n13599 )  ;
assign n13601 =  ( n5802 ) | ( n5811 )  ;
assign n13602 =  ( n13601 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13603 =  ( n13600 ) ^ ( n13602 )  ;
assign n13604 =  ( n5832 ) | ( n5841 )  ;
assign n13605 =  ( n13604 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13606 =  ( n13603 ) ^ ( n13605 )  ;
assign n13607 =  ( n5682 ) | ( n5691 )  ;
assign n13608 =  ( n13607 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13609 =  ( n13606 ) ^ ( n13608 )  ;
assign n13610 =  ( n5713 ) | ( n5722 )  ;
assign n13611 =  ( n13610 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13612 =  ( n13609 ) ^ ( n13611 )  ;
assign n13613 =  ( n13612 ) ^ ( n13466 )  ;
assign n13614 = ~ ( n13613 ) ;
assign n13615 =  ( n13569 ) | ( n13614 )  ;
assign n13616 = ~ ( n13615 ) ;
assign n13617 =  ( n13474 ) | ( n13616 )  ;
assign n13618 = ~ ( n13544 ) ;
assign n13619 = ~ ( n3323 ) ;
assign n13620 =  ( n3306 ) | ( n13619 )  ;
assign n13621 =  ( n3623 ) ^ ( n13620 )  ;
assign n13622 = ~ ( n2928 ) ;
assign n13623 = ~ ( n2939 ) ;
assign n13624 =  ( n13622 ) | ( n13623 )  ;
assign n13625 = ~ ( n2954 ) ;
assign n13626 =  ( n13624 ) | ( n13625 )  ;
assign n13627 =  ( n13621 ) ^ ( n13626 )  ;
assign n13628 =  ( n13627 ) ^ ( n2971 )  ;
assign n13629 =  ( n13628 ) ^ ( n2552 )  ;
assign n13630 =  ( n13629 ) ^ ( n2561 )  ;
assign n13631 =  ( n13630 ) ^ ( n2624 )  ;
assign n13632 =  ( n13631 ) ^ ( n2144 )  ;
assign n13633 =  ( n13632 ) ^ ( n2160 )  ;
assign n13634 =  ( n13633 ) ^ ( n2177 )  ;
assign n13635 =  ( n13634 ) ^ ( n2194 )  ;
assign n13636 =  ( n13635 ) ^ ( n2223 )  ;
assign n13637 =  ( n13636 ) ^ ( n2263 )  ;
assign n13638 =  ( n13637 ) ^ ( n2309 )  ;
assign n13639 =  ( n13638 ) ^ ( n13329 )  ;
assign n13640 =  ( n13639 ) ^ ( n8625 )  ;
assign n13641 =  ( n13640 ) ^ ( n8279 )  ;
assign n13642 =  ( n13641 ) ^ ( n7899 )  ;
assign n13643 = ~ ( n7905 ) ;
assign n13644 = ~ ( n7911 ) ;
assign n13645 =  ( n13643 ) | ( n13644 )  ;
assign n13646 =  ( n13642 ) ^ ( n13645 )  ;
assign n13647 = ~ ( n7467 ) ;
assign n13648 =  ( n7473 ) | ( n6524 )  ;
assign n13649 = ~ ( n13648 ) ;
assign n13650 =  ( n13647 ) | ( n13649 )  ;
assign n13651 = ~ ( n7491 ) ;
assign n13652 =  ( n13650 ) | ( n13651 )  ;
assign n13653 =  ( n13646 ) ^ ( n13652 )  ;
assign n13654 = ~ ( n7498 ) ;
assign n13655 = ~ ( n6553 ) ;
assign n13656 =  ( n13654 ) | ( n13655 )  ;
assign n13657 =  ( n13653 ) ^ ( n13656 )  ;
assign n13658 = ~ ( n5902 ) ;
assign n13659 = ~ ( n5913 ) ;
assign n13660 =  ( n13658 ) | ( n13659 )  ;
assign n13661 =  ( n13657 ) ^ ( n13660 )  ;
assign n13662 =  ( n6825 ) | ( n6834 )  ;
assign n13663 =  ( n13662 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n13664 =  ( n13661 ) ^ ( n13663 )  ;
assign n13665 =  ( n6483 ) | ( n6492 )  ;
assign n13666 =  ( n13665 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13667 =  ( n13664 ) ^ ( n13666 )  ;
assign n13668 =  ( n6030 ) | ( n6039 )  ;
assign n13669 =  ( n13668 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13670 =  ( n13667 ) ^ ( n13669 )  ;
assign n13671 =  ( n5802 ) | ( n5811 )  ;
assign n13672 =  ( n13671 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13673 =  ( n13670 ) ^ ( n13672 )  ;
assign n13674 =  ( n5832 ) | ( n5841 )  ;
assign n13675 =  ( n13674 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13676 =  ( n13673 ) ^ ( n13675 )  ;
assign n13677 =  ( n5682 ) | ( n5691 )  ;
assign n13678 =  ( n13677 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13679 =  ( n13676 ) ^ ( n13678 )  ;
assign n13680 =  ( n5713 ) | ( n5722 )  ;
assign n13681 =  ( n13680 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13682 =  ( n13679 ) ^ ( n13681 )  ;
assign n13683 =  ( n13682 ) ^ ( n13466 )  ;
assign n13684 = ~ ( n13683 ) ;
assign n13685 =  ( n13618 ) | ( n13684 )  ;
assign n13686 = ~ ( n3963 ) ;
assign n13687 =  ( bv_1_1_n5 ) ^ ( n13686 )  ;
assign n13688 = ~ ( n3583 ) ;
assign n13689 =  ( n3567 ) | ( n13688 )  ;
assign n13690 =  ( n13687 ) ^ ( n13689 )  ;
assign n13691 =  ( n3264 ) | ( n3274 )  ;
assign n13692 =  ( n13691 ) | ( n3288 )  ;
assign n13693 =  ( n13690 ) ^ ( n13692 )  ;
assign n13694 =  ( n13693 ) ^ ( n3303 )  ;
assign n13695 =  ( n13694 ) ^ ( n2846 )  ;
assign n13696 =  ( n13695 ) ^ ( n2856 )  ;
assign n13697 =  ( n13696 ) ^ ( n2919 )  ;
assign n13698 = ~ ( n2468 ) ;
assign n13699 =  ( n13697 ) ^ ( n13698 )  ;
assign n13700 =  ( n13699 ) ^ ( n2483 )  ;
assign n13701 =  ( n13700 ) ^ ( n2500 )  ;
assign n13702 =  ( n13701 ) ^ ( n2517 )  ;
assign n13703 =  ( n13702 ) ^ ( n2548 )  ;
assign n13704 =  ( n13703 ) ^ ( n2578 )  ;
assign n13705 =  ( n13704 ) ^ ( n2594 )  ;
assign n13706 =  ( n13705 ) ^ ( n2620 )  ;
assign n13707 =  ( n4123 ) | ( n4142 )  ;
assign n13708 = ~ ( n13707 ) ;
assign n13709 =  ( n13708 ) | ( n4160 )  ;
assign n13710 =  ( n13709 ) | ( n4179 )  ;
assign n13711 = ~ ( n13710 ) ;
assign n13712 = ~ ( n5668 ) ;
assign n13713 =  ( n4253 ) | ( n13712 )  ;
assign n13714 = ~ ( n13713 ) ;
assign n13715 =  ( n13711 ) | ( n13714 )  ;
assign n13716 =  ( n13706 ) ^ ( n13715 )  ;
assign n13717 = ~ ( n13716 ) ;
assign n13718 = ~ ( n8880 ) ;
assign n13719 = ~ ( n8920 ) ;
assign n13720 =  ( n13718 ) | ( n13719 )  ;
assign n13721 = ~ ( n13720 ) ;
assign n13722 =  ( bv_1_1_n5 ) ^ ( n13721 )  ;
assign n13723 =  ( n13722 ) ^ ( n8541 )  ;
assign n13724 =  ( n13723 ) ^ ( n8227 )  ;
assign n13725 =  ( n13724 ) ^ ( n8233 )  ;
assign n13726 = ~ ( n7779 ) ;
assign n13727 =  ( n7784 ) | ( n6524 )  ;
assign n13728 = ~ ( n13727 ) ;
assign n13729 =  ( n13726 ) | ( n13728 )  ;
assign n13730 = ~ ( n7801 ) ;
assign n13731 =  ( n13729 ) | ( n13730 )  ;
assign n13732 =  ( n13725 ) ^ ( n13731 )  ;
assign n13733 = ~ ( n7809 ) ;
assign n13734 = ~ ( n6553 ) ;
assign n13735 =  ( n13733 ) | ( n13734 )  ;
assign n13736 =  ( n13732 ) ^ ( n13735 )  ;
assign n13737 = ~ ( n5902 ) ;
assign n13738 = ~ ( n5913 ) ;
assign n13739 =  ( n13737 ) | ( n13738 )  ;
assign n13740 =  ( n13736 ) ^ ( n13739 )  ;
assign n13741 = ~ ( n7455 ) ;
assign n13742 =  ( n13740 ) ^ ( n13741 )  ;
assign n13743 =  ( n6825 ) | ( n6834 )  ;
assign n13744 =  ( n13743 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n13745 =  ( n13742 ) ^ ( n13744 )  ;
assign n13746 =  ( n6483 ) | ( n6492 )  ;
assign n13747 =  ( n13746 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13748 =  ( n13745 ) ^ ( n13747 )  ;
assign n13749 =  ( n6030 ) | ( n6039 )  ;
assign n13750 =  ( n13749 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13751 =  ( n13748 ) ^ ( n13750 )  ;
assign n13752 =  ( n5802 ) | ( n5811 )  ;
assign n13753 =  ( n13752 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13754 =  ( n13751 ) ^ ( n13753 )  ;
assign n13755 =  ( n5832 ) | ( n5841 )  ;
assign n13756 =  ( n13755 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13757 =  ( n13754 ) ^ ( n13756 )  ;
assign n13758 =  ( n5682 ) | ( n5691 )  ;
assign n13759 =  ( n13758 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13760 =  ( n13757 ) ^ ( n13759 )  ;
assign n13761 =  ( n5713 ) | ( n5722 )  ;
assign n13762 =  ( n13761 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13763 =  ( n13760 ) ^ ( n13762 )  ;
assign n13764 = ~ ( n9088 ) ;
assign n13765 = ~ ( n9126 ) ;
assign n13766 =  ( n13764 ) | ( n13765 )  ;
assign n13767 = ~ ( n9168 ) ;
assign n13768 =  ( n13766 ) | ( n13767 )  ;
assign n13769 = ~ ( n13768 ) ;
assign n13770 = ~ ( n9252 ) ;
assign n13771 = ~ ( n10575 ) ;
assign n13772 =  ( n13770 ) | ( n13771 )  ;
assign n13773 = ~ ( n13772 ) ;
assign n13774 =  ( n13769 ) | ( n13773 )  ;
assign n13775 =  ( n13763 ) ^ ( n13774 )  ;
assign n13776 = ~ ( n13775 ) ;
assign n13777 =  ( n13717 ) | ( n13776 )  ;
assign n13778 = ~ ( n13777 ) ;
assign n13779 = ~ ( n3963 ) ;
assign n13780 = ~ ( n3583 ) ;
assign n13781 =  ( n3567 ) | ( n13780 )  ;
assign n13782 =  ( n13779 ) ^ ( n13781 )  ;
assign n13783 =  ( n3264 ) | ( n3274 )  ;
assign n13784 =  ( n13783 ) | ( n3288 )  ;
assign n13785 =  ( n13782 ) ^ ( n13784 )  ;
assign n13786 =  ( n13785 ) ^ ( n3303 )  ;
assign n13787 =  ( n13786 ) ^ ( n2846 )  ;
assign n13788 =  ( n13787 ) ^ ( n2856 )  ;
assign n13789 =  ( n13788 ) ^ ( n2919 )  ;
assign n13790 = ~ ( n2468 ) ;
assign n13791 =  ( n13789 ) ^ ( n13790 )  ;
assign n13792 =  ( n13791 ) ^ ( n2483 )  ;
assign n13793 =  ( n13792 ) ^ ( n2500 )  ;
assign n13794 =  ( n13793 ) ^ ( n2517 )  ;
assign n13795 =  ( n13794 ) ^ ( n2548 )  ;
assign n13796 =  ( n13795 ) ^ ( n2578 )  ;
assign n13797 =  ( n13796 ) ^ ( n2594 )  ;
assign n13798 =  ( n13797 ) ^ ( n2620 )  ;
assign n13799 =  ( n13798 ) ^ ( n13715 )  ;
assign n13800 = ~ ( n8880 ) ;
assign n13801 = ~ ( n8920 ) ;
assign n13802 =  ( n13800 ) | ( n13801 )  ;
assign n13803 = ~ ( n13802 ) ;
assign n13804 =  ( n13799 ) ^ ( n13803 )  ;
assign n13805 =  ( n13804 ) ^ ( n8541 )  ;
assign n13806 =  ( n13805 ) ^ ( n8227 )  ;
assign n13807 =  ( n13806 ) ^ ( n8233 )  ;
assign n13808 = ~ ( n7779 ) ;
assign n13809 =  ( n7784 ) | ( n6524 )  ;
assign n13810 = ~ ( n13809 ) ;
assign n13811 =  ( n13808 ) | ( n13810 )  ;
assign n13812 = ~ ( n7801 ) ;
assign n13813 =  ( n13811 ) | ( n13812 )  ;
assign n13814 =  ( n13807 ) ^ ( n13813 )  ;
assign n13815 = ~ ( n7809 ) ;
assign n13816 = ~ ( n6553 ) ;
assign n13817 =  ( n13815 ) | ( n13816 )  ;
assign n13818 =  ( n13814 ) ^ ( n13817 )  ;
assign n13819 = ~ ( n5902 ) ;
assign n13820 = ~ ( n5913 ) ;
assign n13821 =  ( n13819 ) | ( n13820 )  ;
assign n13822 =  ( n13818 ) ^ ( n13821 )  ;
assign n13823 = ~ ( n7455 ) ;
assign n13824 =  ( n13822 ) ^ ( n13823 )  ;
assign n13825 =  ( n6825 ) | ( n6834 )  ;
assign n13826 =  ( n13825 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n13827 =  ( n13824 ) ^ ( n13826 )  ;
assign n13828 =  ( n6483 ) | ( n6492 )  ;
assign n13829 =  ( n13828 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13830 =  ( n13827 ) ^ ( n13829 )  ;
assign n13831 =  ( n6030 ) | ( n6039 )  ;
assign n13832 =  ( n13831 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13833 =  ( n13830 ) ^ ( n13832 )  ;
assign n13834 =  ( n5802 ) | ( n5811 )  ;
assign n13835 =  ( n13834 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13836 =  ( n13833 ) ^ ( n13835 )  ;
assign n13837 =  ( n5832 ) | ( n5841 )  ;
assign n13838 =  ( n13837 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13839 =  ( n13836 ) ^ ( n13838 )  ;
assign n13840 =  ( n5682 ) | ( n5691 )  ;
assign n13841 =  ( n13840 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13842 =  ( n13839 ) ^ ( n13841 )  ;
assign n13843 =  ( n5713 ) | ( n5722 )  ;
assign n13844 =  ( n13843 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13845 =  ( n13842 ) ^ ( n13844 )  ;
assign n13846 =  ( n13845 ) ^ ( n13774 )  ;
assign n13847 = ~ ( n13846 ) ;
assign n13848 = ~ ( n3918 ) ;
assign n13849 =  ( n3902 ) | ( n13848 )  ;
assign n13850 =  ( n4234 ) ^ ( n13849 )  ;
assign n13851 =  ( n3519 ) | ( n3531 )  ;
assign n13852 =  ( n13851 ) | ( n3547 )  ;
assign n13853 =  ( n13850 ) ^ ( n13852 )  ;
assign n13854 =  ( n13853 ) ^ ( n3564 )  ;
assign n13855 =  ( n13854 ) ^ ( n3189 )  ;
assign n13856 =  ( n13855 ) ^ ( n3199 )  ;
assign n13857 =  ( n13856 ) ^ ( n3255 )  ;
assign n13858 =  ( n13857 ) ^ ( n2763 )  ;
assign n13859 =  ( n13858 ) ^ ( n2779 )  ;
assign n13860 =  ( n13859 ) ^ ( n2796 )  ;
assign n13861 =  ( n13860 ) ^ ( n2813 )  ;
assign n13862 =  ( n13861 ) ^ ( n2842 )  ;
assign n13863 =  ( n13862 ) ^ ( n2873 )  ;
assign n13864 =  ( n13863 ) ^ ( n2889 )  ;
assign n13865 =  ( n13864 ) ^ ( n2915 )  ;
assign n13866 =  ( n13865 ) ^ ( n5668 )  ;
assign n13867 = ~ ( n13866 ) ;
assign n13868 =  ( n13847 ) | ( n13867 )  ;
assign n13869 = ~ ( n9088 ) ;
assign n13870 = ~ ( n9126 ) ;
assign n13871 =  ( n13869 ) | ( n13870 )  ;
assign n13872 = ~ ( n13871 ) ;
assign n13873 =  ( n13872 ) ^ ( n8880 )  ;
assign n13874 =  ( n13873 ) ^ ( n8490 )  ;
assign n13875 = ~ ( n7905 ) ;
assign n13876 =  ( n8179 ) | ( n8427 )  ;
assign n13877 = ~ ( n13876 ) ;
assign n13878 =  ( n13875 ) | ( n13877 )  ;
assign n13879 =  ( n13874 ) ^ ( n13878 )  ;
assign n13880 = ~ ( n7779 ) ;
assign n13881 =  ( n7784 ) | ( n6524 )  ;
assign n13882 = ~ ( n13881 ) ;
assign n13883 =  ( n13880 ) | ( n13882 )  ;
assign n13884 = ~ ( n7801 ) ;
assign n13885 =  ( n13883 ) | ( n13884 )  ;
assign n13886 =  ( n13879 ) ^ ( n13885 )  ;
assign n13887 = ~ ( n7809 ) ;
assign n13888 = ~ ( n6553 ) ;
assign n13889 =  ( n13887 ) | ( n13888 )  ;
assign n13890 =  ( n13886 ) ^ ( n13889 )  ;
assign n13891 =  ( n13890 ) ^ ( n8164 )  ;
assign n13892 =  ( n13891 ) ^ ( n7455 )  ;
assign n13893 =  ( n6825 ) | ( n6834 )  ;
assign n13894 =  ( n13893 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n13895 =  ( n13892 ) ^ ( n13894 )  ;
assign n13896 =  ( n6483 ) | ( n6492 )  ;
assign n13897 =  ( n13896 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n13898 =  ( n13895 ) ^ ( n13897 )  ;
assign n13899 =  ( n6030 ) | ( n6039 )  ;
assign n13900 =  ( n13899 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n13901 =  ( n13898 ) ^ ( n13900 )  ;
assign n13902 =  ( n5802 ) | ( n5811 )  ;
assign n13903 =  ( n13902 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n13904 =  ( n13901 ) ^ ( n13903 )  ;
assign n13905 =  ( n5832 ) | ( n5841 )  ;
assign n13906 =  ( n13905 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n13907 =  ( n13904 ) ^ ( n13906 )  ;
assign n13908 =  ( n5682 ) | ( n5691 )  ;
assign n13909 =  ( n13908 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n13910 =  ( n13907 ) ^ ( n13909 )  ;
assign n13911 =  ( n5713 ) | ( n5722 )  ;
assign n13912 =  ( n13911 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n13913 =  ( n13910 ) ^ ( n13912 )  ;
assign n13914 =  ( n13913 ) ^ ( n10575 )  ;
assign n13915 = ~ ( n13914 ) ;
assign n13916 =  ( n13868 ) | ( n13915 )  ;
assign n13917 = ~ ( n13916 ) ;
assign n13918 =  ( n13778 ) | ( n13917 )  ;
assign n13919 = ~ ( n13918 ) ;
assign n13920 =  ( n13685 ) | ( n13919 )  ;
assign n13921 = ~ ( n13920 ) ;
assign n13922 =  ( n13617 ) | ( n13921 )  ;
assign n13923 = ~ ( n13922 ) ;
assign n13924 =  ( n13227 ) | ( n13923 )  ;
assign n13925 = ~ ( n13924 ) ;
assign n13926 =  ( n13176 ) | ( n13925 )  ;
assign n13927 = ~ ( n13926 ) ;
assign n13928 =  ( n12427 ) | ( n13927 )  ;
assign n13929 = ~ ( n13928 ) ;
assign n13930 =  ( n12387 ) | ( n13929 )  ;
assign n13931 = ~ ( n11115 ) ;
assign n13932 =  ( n13931 ) | ( n11145 )  ;
assign n13933 = ~ ( n11570 ) ;
assign n13934 =  ( n13932 ) | ( n13933 )  ;
assign n13935 =  ( n13934 ) | ( n11619 )  ;
assign n13936 = ~ ( n12036 ) ;
assign n13937 =  ( n13935 ) | ( n13936 )  ;
assign n13938 =  ( n13937 ) | ( n12090 )  ;
assign n13939 = ~ ( n12343 ) ;
assign n13940 =  ( n13938 ) | ( n13939 )  ;
assign n13941 =  ( n13940 ) | ( n12426 )  ;
assign n13942 = ~ ( n12722 ) ;
assign n13943 =  ( n13941 ) | ( n13942 )  ;
assign n13944 =  ( n13943 ) | ( n12800 )  ;
assign n13945 = ~ ( n13119 ) ;
assign n13946 =  ( n13944 ) | ( n13945 )  ;
assign n13947 =  ( n13946 ) | ( n13226 )  ;
assign n13948 = ~ ( n13544 ) ;
assign n13949 =  ( n13947 ) | ( n13948 )  ;
assign n13950 = ~ ( n13683 ) ;
assign n13951 =  ( n13949 ) | ( n13950 )  ;
assign n13952 = ~ ( n13846 ) ;
assign n13953 =  ( n13951 ) | ( n13952 )  ;
assign n13954 = ~ ( n3918 ) ;
assign n13955 =  ( n3902 ) | ( n13954 )  ;
assign n13956 =  ( n4234 ) ^ ( n13955 )  ;
assign n13957 =  ( n3519 ) | ( n3531 )  ;
assign n13958 =  ( n13957 ) | ( n3547 )  ;
assign n13959 =  ( n13956 ) ^ ( n13958 )  ;
assign n13960 =  ( n13959 ) ^ ( n3564 )  ;
assign n13961 =  ( n13960 ) ^ ( n3189 )  ;
assign n13962 =  ( n13961 ) ^ ( n3199 )  ;
assign n13963 =  ( n13962 ) ^ ( n3255 )  ;
assign n13964 =  ( n13963 ) ^ ( n2763 )  ;
assign n13965 =  ( n13964 ) ^ ( n2779 )  ;
assign n13966 =  ( n13965 ) ^ ( n2796 )  ;
assign n13967 =  ( n13966 ) ^ ( n2813 )  ;
assign n13968 =  ( n13967 ) ^ ( n2842 )  ;
assign n13969 =  ( n13968 ) ^ ( n2873 )  ;
assign n13970 =  ( n13969 ) ^ ( n2889 )  ;
assign n13971 =  ( n13970 ) ^ ( n2915 )  ;
assign n13972 =  ( n13971 ) ^ ( n5668 )  ;
assign n13973 = ~ ( n9088 ) ;
assign n13974 = ~ ( n9126 ) ;
assign n13975 =  ( n13973 ) | ( n13974 )  ;
assign n13976 = ~ ( n13975 ) ;
assign n13977 =  ( n13972 ) ^ ( n13976 )  ;
assign n13978 =  ( n13977 ) ^ ( n8880 )  ;
assign n13979 =  ( n13978 ) ^ ( n8490 )  ;
assign n13980 = ~ ( n7905 ) ;
assign n13981 =  ( n8179 ) | ( n8427 )  ;
assign n13982 = ~ ( n13981 ) ;
assign n13983 =  ( n13980 ) | ( n13982 )  ;
assign n13984 =  ( n13979 ) ^ ( n13983 )  ;
assign n13985 = ~ ( n7779 ) ;
assign n13986 =  ( n7784 ) | ( n6524 )  ;
assign n13987 = ~ ( n13986 ) ;
assign n13988 =  ( n13985 ) | ( n13987 )  ;
assign n13989 = ~ ( n7801 ) ;
assign n13990 =  ( n13988 ) | ( n13989 )  ;
assign n13991 =  ( n13984 ) ^ ( n13990 )  ;
assign n13992 = ~ ( n7809 ) ;
assign n13993 = ~ ( n6553 ) ;
assign n13994 =  ( n13992 ) | ( n13993 )  ;
assign n13995 =  ( n13991 ) ^ ( n13994 )  ;
assign n13996 =  ( n13995 ) ^ ( n8164 )  ;
assign n13997 =  ( n13996 ) ^ ( n7455 )  ;
assign n13998 =  ( n6825 ) | ( n6834 )  ;
assign n13999 =  ( n13998 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14000 =  ( n13997 ) ^ ( n13999 )  ;
assign n14001 =  ( n6483 ) | ( n6492 )  ;
assign n14002 =  ( n14001 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14003 =  ( n14000 ) ^ ( n14002 )  ;
assign n14004 =  ( n6030 ) | ( n6039 )  ;
assign n14005 =  ( n14004 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14006 =  ( n14003 ) ^ ( n14005 )  ;
assign n14007 =  ( n5802 ) | ( n5811 )  ;
assign n14008 =  ( n14007 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14009 =  ( n14006 ) ^ ( n14008 )  ;
assign n14010 =  ( n5832 ) | ( n5841 )  ;
assign n14011 =  ( n14010 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14012 =  ( n14009 ) ^ ( n14011 )  ;
assign n14013 =  ( n5682 ) | ( n5691 )  ;
assign n14014 =  ( n14013 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n14015 =  ( n14012 ) ^ ( n14014 )  ;
assign n14016 =  ( n5713 ) | ( n5722 )  ;
assign n14017 =  ( n14016 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n14018 =  ( n14015 ) ^ ( n14017 )  ;
assign n14019 =  ( n14018 ) ^ ( n10575 )  ;
assign n14020 = ~ ( n14019 ) ;
assign n14021 =  ( n13953 ) | ( n14020 )  ;
assign n14022 =  ( n4123 ) | ( n4142 )  ;
assign n14023 =  ( n4440 ) ^ ( n14022 )  ;
assign n14024 =  ( n3856 ) | ( n3866 )  ;
assign n14025 =  ( n14024 ) | ( n3884 )  ;
assign n14026 =  ( n14023 ) ^ ( n14025 )  ;
assign n14027 =  ( n14026 ) ^ ( n3899 )  ;
assign n14028 =  ( n14027 ) ^ ( n3496 )  ;
assign n14029 =  ( n14028 ) ^ ( n3506 )  ;
assign n14030 =  ( n14029 ) ^ ( n3106 )  ;
assign n14031 =  ( n14030 ) ^ ( n3122 )  ;
assign n14032 =  ( n14031 ) ^ ( n3139 )  ;
assign n14033 =  ( n14032 ) ^ ( n3156 )  ;
assign n14034 =  ( n14033 ) ^ ( n3185 )  ;
assign n14035 =  ( n14034 ) ^ ( n3216 )  ;
assign n14036 =  ( n14035 ) ^ ( n3232 )  ;
assign n14037 =  ( n14036 ) ^ ( n3251 )  ;
assign n14038 =  ( n14037 ) ^ ( n3248 )  ;
assign n14039 = ~ ( n4659 ) ;
assign n14040 =  ( n4647 ) | ( n14039 )  ;
assign n14041 = ~ ( n14040 ) ;
assign n14042 =  ( n14041 ) | ( n4674 )  ;
assign n14043 =  ( n14042 ) | ( n4688 )  ;
assign n14044 = ~ ( n14043 ) ;
assign n14045 = ~ ( n10841 ) ;
assign n14046 =  ( n4710 ) | ( n14045 )  ;
assign n14047 = ~ ( n14046 ) ;
assign n14048 =  ( n14044 ) | ( n14047 )  ;
assign n14049 =  ( n14038 ) ^ ( n14048 )  ;
assign n14050 = ~ ( n14049 ) ;
assign n14051 = ~ ( n9314 ) ;
assign n14052 = ~ ( n9348 ) ;
assign n14053 =  ( n14051 ) | ( n14052 )  ;
assign n14054 = ~ ( n14053 ) ;
assign n14055 =  ( n14054 ) ^ ( n9088 )  ;
assign n14056 =  ( n14055 ) ^ ( n8829 )  ;
assign n14057 = ~ ( n7905 ) ;
assign n14058 = ~ ( n8835 ) ;
assign n14059 =  ( n14057 ) | ( n14058 )  ;
assign n14060 =  ( n14056 ) ^ ( n14059 )  ;
assign n14061 = ~ ( n7779 ) ;
assign n14062 =  ( n7784 ) | ( n6524 )  ;
assign n14063 = ~ ( n14062 ) ;
assign n14064 =  ( n14061 ) | ( n14063 )  ;
assign n14065 = ~ ( n7801 ) ;
assign n14066 =  ( n14064 ) | ( n14065 )  ;
assign n14067 =  ( n14060 ) ^ ( n14066 )  ;
assign n14068 = ~ ( n7809 ) ;
assign n14069 = ~ ( n6553 ) ;
assign n14070 =  ( n14068 ) | ( n14069 )  ;
assign n14071 =  ( n14067 ) ^ ( n14070 )  ;
assign n14072 =  ( n14071 ) ^ ( n7455 )  ;
assign n14073 =  ( n6825 ) | ( n6834 )  ;
assign n14074 =  ( n14073 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14075 =  ( n14072 ) ^ ( n14074 )  ;
assign n14076 =  ( n6483 ) | ( n6492 )  ;
assign n14077 =  ( n14076 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14078 =  ( n14075 ) ^ ( n14077 )  ;
assign n14079 =  ( n6030 ) | ( n6039 )  ;
assign n14080 =  ( n14079 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14081 =  ( n14078 ) ^ ( n14080 )  ;
assign n14082 =  ( n5802 ) | ( n5811 )  ;
assign n14083 =  ( n14082 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14084 =  ( n14081 ) ^ ( n14083 )  ;
assign n14085 =  ( n5832 ) | ( n5841 )  ;
assign n14086 =  ( n14085 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14087 =  ( n14084 ) ^ ( n14086 )  ;
assign n14088 =  ( n5682 ) | ( n5691 )  ;
assign n14089 =  ( n14088 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n14090 =  ( n14087 ) ^ ( n14089 )  ;
assign n14091 =  ( n14090 ) ^ ( n8160 )  ;
assign n14092 =  ( n14091 ) ^ ( n8157 )  ;
assign n14093 = ~ ( n9538 ) ;
assign n14094 = ~ ( n9569 ) ;
assign n14095 =  ( n14093 ) | ( n14094 )  ;
assign n14096 = ~ ( n9605 ) ;
assign n14097 =  ( n14095 ) | ( n14096 )  ;
assign n14098 = ~ ( n14097 ) ;
assign n14099 = ~ ( n9649 ) ;
assign n14100 = ~ ( n11090 ) ;
assign n14101 =  ( n14099 ) | ( n14100 )  ;
assign n14102 = ~ ( n14101 ) ;
assign n14103 =  ( n14098 ) | ( n14102 )  ;
assign n14104 =  ( n14092 ) ^ ( n14103 )  ;
assign n14105 = ~ ( n14104 ) ;
assign n14106 =  ( n14050 ) | ( n14105 )  ;
assign n14107 = ~ ( n14106 ) ;
assign n14108 =  ( n4123 ) | ( n4142 )  ;
assign n14109 =  ( n4440 ) ^ ( n14108 )  ;
assign n14110 =  ( n3856 ) | ( n3866 )  ;
assign n14111 =  ( n14110 ) | ( n3884 )  ;
assign n14112 =  ( n14109 ) ^ ( n14111 )  ;
assign n14113 =  ( n14112 ) ^ ( n3899 )  ;
assign n14114 =  ( n14113 ) ^ ( n3496 )  ;
assign n14115 =  ( n14114 ) ^ ( n3506 )  ;
assign n14116 =  ( n14115 ) ^ ( n3106 )  ;
assign n14117 =  ( n14116 ) ^ ( n3122 )  ;
assign n14118 =  ( n14117 ) ^ ( n3139 )  ;
assign n14119 =  ( n14118 ) ^ ( n3156 )  ;
assign n14120 =  ( n14119 ) ^ ( n3185 )  ;
assign n14121 =  ( n14120 ) ^ ( n3216 )  ;
assign n14122 =  ( n14121 ) ^ ( n3232 )  ;
assign n14123 =  ( n14122 ) ^ ( n3251 )  ;
assign n14124 =  ( n14123 ) ^ ( n3248 )  ;
assign n14125 =  ( n14124 ) ^ ( n14048 )  ;
assign n14126 = ~ ( n9314 ) ;
assign n14127 = ~ ( n9348 ) ;
assign n14128 =  ( n14126 ) | ( n14127 )  ;
assign n14129 = ~ ( n14128 ) ;
assign n14130 =  ( n14125 ) ^ ( n14129 )  ;
assign n14131 =  ( n14130 ) ^ ( n9088 )  ;
assign n14132 =  ( n14131 ) ^ ( n8829 )  ;
assign n14133 = ~ ( n7905 ) ;
assign n14134 = ~ ( n8835 ) ;
assign n14135 =  ( n14133 ) | ( n14134 )  ;
assign n14136 =  ( n14132 ) ^ ( n14135 )  ;
assign n14137 = ~ ( n7779 ) ;
assign n14138 =  ( n7784 ) | ( n6524 )  ;
assign n14139 = ~ ( n14138 ) ;
assign n14140 =  ( n14137 ) | ( n14139 )  ;
assign n14141 = ~ ( n7801 ) ;
assign n14142 =  ( n14140 ) | ( n14141 )  ;
assign n14143 =  ( n14136 ) ^ ( n14142 )  ;
assign n14144 = ~ ( n7809 ) ;
assign n14145 = ~ ( n6553 ) ;
assign n14146 =  ( n14144 ) | ( n14145 )  ;
assign n14147 =  ( n14143 ) ^ ( n14146 )  ;
assign n14148 =  ( n14147 ) ^ ( n7455 )  ;
assign n14149 =  ( n6825 ) | ( n6834 )  ;
assign n14150 =  ( n14149 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14151 =  ( n14148 ) ^ ( n14150 )  ;
assign n14152 =  ( n6483 ) | ( n6492 )  ;
assign n14153 =  ( n14152 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14154 =  ( n14151 ) ^ ( n14153 )  ;
assign n14155 =  ( n6030 ) | ( n6039 )  ;
assign n14156 =  ( n14155 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14157 =  ( n14154 ) ^ ( n14156 )  ;
assign n14158 =  ( n5802 ) | ( n5811 )  ;
assign n14159 =  ( n14158 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14160 =  ( n14157 ) ^ ( n14159 )  ;
assign n14161 =  ( n5832 ) | ( n5841 )  ;
assign n14162 =  ( n14161 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14163 =  ( n14160 ) ^ ( n14162 )  ;
assign n14164 =  ( n5682 ) | ( n5691 )  ;
assign n14165 =  ( n14164 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n14166 =  ( n14163 ) ^ ( n14165 )  ;
assign n14167 =  ( n14166 ) ^ ( n8160 )  ;
assign n14168 =  ( n14167 ) ^ ( n8157 )  ;
assign n14169 =  ( n14168 ) ^ ( n14103 )  ;
assign n14170 = ~ ( n14169 ) ;
assign n14171 = ~ ( n4695 ) ;
assign n14172 =  ( n4390 ) | ( n4403 )  ;
assign n14173 =  ( n14171 ) ^ ( n14172 )  ;
assign n14174 =  ( n14173 ) ^ ( n4111 )  ;
assign n14175 =  ( n14174 ) ^ ( n3776 )  ;
assign n14176 =  ( n14175 ) ^ ( n3786 )  ;
assign n14177 =  ( n14176 ) ^ ( n3847 )  ;
assign n14178 =  ( n14177 ) ^ ( n3413 )  ;
assign n14179 =  ( n14178 ) ^ ( n3429 )  ;
assign n14180 =  ( n14179 ) ^ ( n3446 )  ;
assign n14181 =  ( n14180 ) ^ ( n3463 )  ;
assign n14182 =  ( n14181 ) ^ ( n3492 )  ;
assign n14183 =  ( n14182 ) ^ ( n3881 )  ;
assign n14184 =  ( n14183 ) ^ ( n4139 )  ;
assign n14185 =  ( n14184 ) ^ ( n10841 )  ;
assign n14186 = ~ ( n14185 ) ;
assign n14187 =  ( n14170 ) | ( n14186 )  ;
assign n14188 = ~ ( n9538 ) ;
assign n14189 = ~ ( n9569 ) ;
assign n14190 =  ( n14188 ) | ( n14189 )  ;
assign n14191 = ~ ( n14190 ) ;
assign n14192 =  ( n14191 ) ^ ( n9314 )  ;
assign n14193 =  ( n14192 ) ^ ( n9018 )  ;
assign n14194 = ~ ( n7779 ) ;
assign n14195 =  ( n7784 ) | ( n6524 )  ;
assign n14196 = ~ ( n14195 ) ;
assign n14197 =  ( n14194 ) | ( n14196 )  ;
assign n14198 = ~ ( n7801 ) ;
assign n14199 =  ( n14197 ) | ( n14198 )  ;
assign n14200 =  ( n14193 ) ^ ( n14199 )  ;
assign n14201 = ~ ( n7809 ) ;
assign n14202 = ~ ( n6553 ) ;
assign n14203 =  ( n14201 ) | ( n14202 )  ;
assign n14204 =  ( n14200 ) ^ ( n14203 )  ;
assign n14205 = ~ ( n8761 ) ;
assign n14206 =  ( n14205 ) | ( n8771 )  ;
assign n14207 =  ( n14204 ) ^ ( n14206 )  ;
assign n14208 =  ( n14207 ) ^ ( n7455 )  ;
assign n14209 =  ( n6825 ) | ( n6834 )  ;
assign n14210 =  ( n14209 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14211 =  ( n14208 ) ^ ( n14210 )  ;
assign n14212 =  ( n6483 ) | ( n6492 )  ;
assign n14213 =  ( n14212 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14214 =  ( n14211 ) ^ ( n14213 )  ;
assign n14215 =  ( n6030 ) | ( n6039 )  ;
assign n14216 =  ( n14215 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14217 =  ( n14214 ) ^ ( n14216 )  ;
assign n14218 =  ( n5802 ) | ( n5811 )  ;
assign n14219 =  ( n14218 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14220 =  ( n14217 ) ^ ( n14219 )  ;
assign n14221 =  ( n5832 ) | ( n5841 )  ;
assign n14222 =  ( n14221 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14223 =  ( n14220 ) ^ ( n14222 )  ;
assign n14224 =  ( n5682 ) | ( n5691 )  ;
assign n14225 =  ( n14224 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n14226 =  ( n14223 ) ^ ( n14225 )  ;
assign n14227 =  ( n14226 ) ^ ( n11090 )  ;
assign n14228 = ~ ( n14227 ) ;
assign n14229 =  ( n14187 ) | ( n14228 )  ;
assign n14230 = ~ ( n14229 ) ;
assign n14231 =  ( n14107 ) | ( n14230 )  ;
assign n14232 = ~ ( n14169 ) ;
assign n14233 = ~ ( n4695 ) ;
assign n14234 =  ( n4390 ) | ( n4403 )  ;
assign n14235 =  ( n14233 ) ^ ( n14234 )  ;
assign n14236 =  ( n14235 ) ^ ( n4111 )  ;
assign n14237 =  ( n14236 ) ^ ( n3776 )  ;
assign n14238 =  ( n14237 ) ^ ( n3786 )  ;
assign n14239 =  ( n14238 ) ^ ( n3847 )  ;
assign n14240 =  ( n14239 ) ^ ( n3413 )  ;
assign n14241 =  ( n14240 ) ^ ( n3429 )  ;
assign n14242 =  ( n14241 ) ^ ( n3446 )  ;
assign n14243 =  ( n14242 ) ^ ( n3463 )  ;
assign n14244 =  ( n14243 ) ^ ( n3492 )  ;
assign n14245 =  ( n14244 ) ^ ( n3881 )  ;
assign n14246 =  ( n14245 ) ^ ( n4139 )  ;
assign n14247 =  ( n14246 ) ^ ( n10841 )  ;
assign n14248 = ~ ( n9538 ) ;
assign n14249 = ~ ( n9569 ) ;
assign n14250 =  ( n14248 ) | ( n14249 )  ;
assign n14251 = ~ ( n14250 ) ;
assign n14252 =  ( n14247 ) ^ ( n14251 )  ;
assign n14253 =  ( n14252 ) ^ ( n9314 )  ;
assign n14254 =  ( n14253 ) ^ ( n9018 )  ;
assign n14255 = ~ ( n7779 ) ;
assign n14256 =  ( n7784 ) | ( n6524 )  ;
assign n14257 = ~ ( n14256 ) ;
assign n14258 =  ( n14255 ) | ( n14257 )  ;
assign n14259 = ~ ( n7801 ) ;
assign n14260 =  ( n14258 ) | ( n14259 )  ;
assign n14261 =  ( n14254 ) ^ ( n14260 )  ;
assign n14262 = ~ ( n7809 ) ;
assign n14263 = ~ ( n6553 ) ;
assign n14264 =  ( n14262 ) | ( n14263 )  ;
assign n14265 =  ( n14261 ) ^ ( n14264 )  ;
assign n14266 = ~ ( n8761 ) ;
assign n14267 =  ( n14266 ) | ( n8771 )  ;
assign n14268 =  ( n14265 ) ^ ( n14267 )  ;
assign n14269 =  ( n14268 ) ^ ( n7455 )  ;
assign n14270 =  ( n6825 ) | ( n6834 )  ;
assign n14271 =  ( n14270 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14272 =  ( n14269 ) ^ ( n14271 )  ;
assign n14273 =  ( n6483 ) | ( n6492 )  ;
assign n14274 =  ( n14273 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14275 =  ( n14272 ) ^ ( n14274 )  ;
assign n14276 =  ( n6030 ) | ( n6039 )  ;
assign n14277 =  ( n14276 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14278 =  ( n14275 ) ^ ( n14277 )  ;
assign n14279 =  ( n5802 ) | ( n5811 )  ;
assign n14280 =  ( n14279 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14281 =  ( n14278 ) ^ ( n14280 )  ;
assign n14282 =  ( n5832 ) | ( n5841 )  ;
assign n14283 =  ( n14282 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14284 =  ( n14281 ) ^ ( n14283 )  ;
assign n14285 =  ( n5682 ) | ( n5691 )  ;
assign n14286 =  ( n14285 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n14287 =  ( n14284 ) ^ ( n14286 )  ;
assign n14288 =  ( n14287 ) ^ ( n11090 )  ;
assign n14289 = ~ ( n14288 ) ;
assign n14290 =  ( n14232 ) | ( n14289 )  ;
assign n14291 = ~ ( n4728 ) ;
assign n14292 =  ( n4722 ) | ( n14291 )  ;
assign n14293 = ~ ( n14292 ) ;
assign n14294 = ~ ( n4659 ) ;
assign n14295 =  ( n4647 ) | ( n14294 )  ;
assign n14296 =  ( n14293 ) ^ ( n14295 )  ;
assign n14297 =  ( n14296 ) ^ ( n4380 )  ;
assign n14298 =  ( n14297 ) ^ ( n4088 )  ;
assign n14299 =  ( n14298 ) ^ ( n4098 )  ;
assign n14300 =  ( n14299 ) ^ ( n3693 )  ;
assign n14301 =  ( n14300 ) ^ ( n3709 )  ;
assign n14302 =  ( n14301 ) ^ ( n3726 )  ;
assign n14303 =  ( n14302 ) ^ ( n3743 )  ;
assign n14304 =  ( n14303 ) ^ ( n3772 )  ;
assign n14305 =  ( n14304 ) ^ ( n3812 )  ;
assign n14306 =  ( n14305 ) ^ ( n3836 )  ;
assign n14307 =  ( n14306 ) ^ ( n3824 )  ;
assign n14308 = ~ ( n4889 ) ;
assign n14309 =  ( n14308 ) | ( n4900 )  ;
assign n14310 =  ( n14309 ) | ( n4913 )  ;
assign n14311 = ~ ( n14310 ) ;
assign n14312 = ~ ( n4938 ) ;
assign n14313 =  ( n5041 ) | ( n5203 )  ;
assign n14314 =  ( n14313 ) | ( n5345 )  ;
assign n14315 =  ( n14314 ) | ( n11288 )  ;
assign n14316 =  ( n14315 ) | ( n11331 )  ;
assign n14317 = ~ ( n14316 ) ;
assign n14318 =  ( n14312 ) | ( n14317 )  ;
assign n14319 = ~ ( n14318 ) ;
assign n14320 =  ( n14311 ) | ( n14319 )  ;
assign n14321 =  ( n14307 ) ^ ( n14320 )  ;
assign n14322 = ~ ( n14321 ) ;
assign n14323 = ~ ( n9719 ) ;
assign n14324 =  ( n14323 ) ^ ( n9538 )  ;
assign n14325 =  ( n14324 ) ^ ( n9018 )  ;
assign n14326 = ~ ( n7779 ) ;
assign n14327 =  ( n7784 ) | ( n6524 )  ;
assign n14328 = ~ ( n14327 ) ;
assign n14329 =  ( n14326 ) | ( n14328 )  ;
assign n14330 = ~ ( n7801 ) ;
assign n14331 =  ( n14329 ) | ( n14330 )  ;
assign n14332 =  ( n14325 ) ^ ( n14331 )  ;
assign n14333 = ~ ( n7809 ) ;
assign n14334 = ~ ( n6553 ) ;
assign n14335 =  ( n14333 ) | ( n14334 )  ;
assign n14336 =  ( n14332 ) ^ ( n14335 )  ;
assign n14337 =  ( n14336 ) ^ ( n7455 )  ;
assign n14338 =  ( n6825 ) | ( n6834 )  ;
assign n14339 =  ( n14338 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14340 =  ( n14337 ) ^ ( n14339 )  ;
assign n14341 =  ( n6483 ) | ( n6492 )  ;
assign n14342 =  ( n14341 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14343 =  ( n14340 ) ^ ( n14342 )  ;
assign n14344 =  ( n6030 ) | ( n6039 )  ;
assign n14345 =  ( n14344 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14346 =  ( n14343 ) ^ ( n14345 )  ;
assign n14347 =  ( n5802 ) | ( n5811 )  ;
assign n14348 =  ( n14347 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14349 =  ( n14346 ) ^ ( n14348 )  ;
assign n14350 =  ( n5832 ) | ( n5841 )  ;
assign n14351 =  ( n14350 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14352 =  ( n14349 ) ^ ( n14351 )  ;
assign n14353 =  ( n14352 ) ^ ( n8759 )  ;
assign n14354 =  ( n14353 ) ^ ( n8756 )  ;
assign n14355 = ~ ( n9834 ) ;
assign n14356 =  ( n9808 ) | ( n14355 )  ;
assign n14357 = ~ ( n9864 ) ;
assign n14358 =  ( n14356 ) | ( n14357 )  ;
assign n14359 = ~ ( n14358 ) ;
assign n14360 = ~ ( n9909 ) ;
assign n14361 = ~ ( n11533 ) ;
assign n14362 =  ( n14360 ) | ( n14361 )  ;
assign n14363 = ~ ( n14362 ) ;
assign n14364 =  ( n14359 ) | ( n14363 )  ;
assign n14365 =  ( n14354 ) ^ ( n14364 )  ;
assign n14366 = ~ ( n14365 ) ;
assign n14367 =  ( n14322 ) | ( n14366 )  ;
assign n14368 = ~ ( n14367 ) ;
assign n14369 = ~ ( n4728 ) ;
assign n14370 =  ( n4722 ) | ( n14369 )  ;
assign n14371 = ~ ( n14370 ) ;
assign n14372 = ~ ( n4659 ) ;
assign n14373 =  ( n4647 ) | ( n14372 )  ;
assign n14374 =  ( n14371 ) ^ ( n14373 )  ;
assign n14375 =  ( n14374 ) ^ ( n4380 )  ;
assign n14376 =  ( n14375 ) ^ ( n4088 )  ;
assign n14377 =  ( n14376 ) ^ ( n4098 )  ;
assign n14378 =  ( n14377 ) ^ ( n3693 )  ;
assign n14379 =  ( n14378 ) ^ ( n3709 )  ;
assign n14380 =  ( n14379 ) ^ ( n3726 )  ;
assign n14381 =  ( n14380 ) ^ ( n3743 )  ;
assign n14382 =  ( n14381 ) ^ ( n3772 )  ;
assign n14383 =  ( n14382 ) ^ ( n3812 )  ;
assign n14384 =  ( n14383 ) ^ ( n3836 )  ;
assign n14385 =  ( n14384 ) ^ ( n3824 )  ;
assign n14386 =  ( n14385 ) ^ ( n14320 )  ;
assign n14387 = ~ ( n9719 ) ;
assign n14388 =  ( n14386 ) ^ ( n14387 )  ;
assign n14389 =  ( n14388 ) ^ ( n9538 )  ;
assign n14390 =  ( n14389 ) ^ ( n9018 )  ;
assign n14391 = ~ ( n7779 ) ;
assign n14392 =  ( n7784 ) | ( n6524 )  ;
assign n14393 = ~ ( n14392 ) ;
assign n14394 =  ( n14391 ) | ( n14393 )  ;
assign n14395 = ~ ( n7801 ) ;
assign n14396 =  ( n14394 ) | ( n14395 )  ;
assign n14397 =  ( n14390 ) ^ ( n14396 )  ;
assign n14398 = ~ ( n7809 ) ;
assign n14399 = ~ ( n6553 ) ;
assign n14400 =  ( n14398 ) | ( n14399 )  ;
assign n14401 =  ( n14397 ) ^ ( n14400 )  ;
assign n14402 =  ( n14401 ) ^ ( n7455 )  ;
assign n14403 =  ( n6825 ) | ( n6834 )  ;
assign n14404 =  ( n14403 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14405 =  ( n14402 ) ^ ( n14404 )  ;
assign n14406 =  ( n6483 ) | ( n6492 )  ;
assign n14407 =  ( n14406 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14408 =  ( n14405 ) ^ ( n14407 )  ;
assign n14409 =  ( n6030 ) | ( n6039 )  ;
assign n14410 =  ( n14409 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14411 =  ( n14408 ) ^ ( n14410 )  ;
assign n14412 =  ( n5802 ) | ( n5811 )  ;
assign n14413 =  ( n14412 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14414 =  ( n14411 ) ^ ( n14413 )  ;
assign n14415 =  ( n5832 ) | ( n5841 )  ;
assign n14416 =  ( n14415 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14417 =  ( n14414 ) ^ ( n14416 )  ;
assign n14418 =  ( n14417 ) ^ ( n8759 )  ;
assign n14419 =  ( n14418 ) ^ ( n8756 )  ;
assign n14420 =  ( n14419 ) ^ ( n14364 )  ;
assign n14421 = ~ ( n14420 ) ;
assign n14422 = ~ ( n4889 ) ;
assign n14423 =  ( n14422 ) | ( n4900 )  ;
assign n14424 = ~ ( n14423 ) ;
assign n14425 =  ( n4605 ) | ( n4615 )  ;
assign n14426 =  ( n14425 ) | ( n4629 )  ;
assign n14427 =  ( n14424 ) ^ ( n14426 )  ;
assign n14428 =  ( n14427 ) ^ ( n4644 )  ;
assign n14429 =  ( n14428 ) ^ ( n4357 )  ;
assign n14430 =  ( n14429 ) ^ ( n4367 )  ;
assign n14431 =  ( n14430 ) ^ ( n4005 )  ;
assign n14432 =  ( n14431 ) ^ ( n4021 )  ;
assign n14433 =  ( n14432 ) ^ ( n4038 )  ;
assign n14434 =  ( n14433 ) ^ ( n4055 )  ;
assign n14435 =  ( n14434 ) ^ ( n4084 )  ;
assign n14436 =  ( n14435 ) ^ ( n4728 )  ;
assign n14437 =  ( n5041 ) | ( n5203 )  ;
assign n14438 =  ( n14437 ) | ( n5345 )  ;
assign n14439 =  ( n14438 ) | ( n11288 )  ;
assign n14440 =  ( n14439 ) | ( n11331 )  ;
assign n14441 =  ( n14436 ) ^ ( n14440 )  ;
assign n14442 = ~ ( n14441 ) ;
assign n14443 =  ( n14421 ) | ( n14442 )  ;
assign n14444 = ~ ( n9834 ) ;
assign n14445 =  ( n9808 ) | ( n14444 )  ;
assign n14446 = ~ ( n14445 ) ;
assign n14447 =  ( n14446 ) ^ ( n9523 )  ;
assign n14448 =  ( n14447 ) ^ ( n9529 )  ;
assign n14449 = ~ ( n7779 ) ;
assign n14450 =  ( n7784 ) | ( n6524 )  ;
assign n14451 = ~ ( n14450 ) ;
assign n14452 =  ( n14449 ) | ( n14451 )  ;
assign n14453 = ~ ( n7801 ) ;
assign n14454 =  ( n14452 ) | ( n14453 )  ;
assign n14455 =  ( n14448 ) ^ ( n14454 )  ;
assign n14456 = ~ ( n7809 ) ;
assign n14457 = ~ ( n6553 ) ;
assign n14458 =  ( n14456 ) | ( n14457 )  ;
assign n14459 =  ( n14455 ) ^ ( n14458 )  ;
assign n14460 =  ( n14459 ) ^ ( n7455 )  ;
assign n14461 =  ( n6825 ) | ( n6834 )  ;
assign n14462 =  ( n14461 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14463 =  ( n14460 ) ^ ( n14462 )  ;
assign n14464 =  ( n6483 ) | ( n6492 )  ;
assign n14465 =  ( n14464 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14466 =  ( n14463 ) ^ ( n14465 )  ;
assign n14467 =  ( n6030 ) | ( n6039 )  ;
assign n14468 =  ( n14467 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14469 =  ( n14466 ) ^ ( n14468 )  ;
assign n14470 =  ( n5802 ) | ( n5811 )  ;
assign n14471 =  ( n14470 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14472 =  ( n14469 ) ^ ( n14471 )  ;
assign n14473 =  ( n5832 ) | ( n5841 )  ;
assign n14474 =  ( n14473 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14475 =  ( n14472 ) ^ ( n14474 )  ;
assign n14476 =  ( n14475 ) ^ ( n11533 )  ;
assign n14477 = ~ ( n14476 ) ;
assign n14478 =  ( n14443 ) | ( n14477 )  ;
assign n14479 = ~ ( n14478 ) ;
assign n14480 =  ( n14368 ) | ( n14479 )  ;
assign n14481 = ~ ( n14480 ) ;
assign n14482 =  ( n14290 ) | ( n14481 )  ;
assign n14483 = ~ ( n14482 ) ;
assign n14484 =  ( n14231 ) | ( n14483 )  ;
assign n14485 = ~ ( n14169 ) ;
assign n14486 = ~ ( n14288 ) ;
assign n14487 =  ( n14485 ) | ( n14486 )  ;
assign n14488 = ~ ( n14420 ) ;
assign n14489 =  ( n14487 ) | ( n14488 )  ;
assign n14490 = ~ ( n4889 ) ;
assign n14491 =  ( n14490 ) | ( n4900 )  ;
assign n14492 = ~ ( n14491 ) ;
assign n14493 =  ( n4605 ) | ( n4615 )  ;
assign n14494 =  ( n14493 ) | ( n4629 )  ;
assign n14495 =  ( n14492 ) ^ ( n14494 )  ;
assign n14496 =  ( n14495 ) ^ ( n4644 )  ;
assign n14497 =  ( n14496 ) ^ ( n4357 )  ;
assign n14498 =  ( n14497 ) ^ ( n4367 )  ;
assign n14499 =  ( n14498 ) ^ ( n4005 )  ;
assign n14500 =  ( n14499 ) ^ ( n4021 )  ;
assign n14501 =  ( n14500 ) ^ ( n4038 )  ;
assign n14502 =  ( n14501 ) ^ ( n4055 )  ;
assign n14503 =  ( n14502 ) ^ ( n4084 )  ;
assign n14504 =  ( n14503 ) ^ ( n4728 )  ;
assign n14505 =  ( n5041 ) | ( n5203 )  ;
assign n14506 =  ( n14505 ) | ( n5345 )  ;
assign n14507 =  ( n14506 ) | ( n11288 )  ;
assign n14508 =  ( n14507 ) | ( n11331 )  ;
assign n14509 =  ( n14504 ) ^ ( n14508 )  ;
assign n14510 = ~ ( n9834 ) ;
assign n14511 =  ( n9808 ) | ( n14510 )  ;
assign n14512 = ~ ( n14511 ) ;
assign n14513 =  ( n14509 ) ^ ( n14512 )  ;
assign n14514 =  ( n14513 ) ^ ( n9523 )  ;
assign n14515 =  ( n14514 ) ^ ( n9529 )  ;
assign n14516 = ~ ( n7779 ) ;
assign n14517 =  ( n7784 ) | ( n6524 )  ;
assign n14518 = ~ ( n14517 ) ;
assign n14519 =  ( n14516 ) | ( n14518 )  ;
assign n14520 = ~ ( n7801 ) ;
assign n14521 =  ( n14519 ) | ( n14520 )  ;
assign n14522 =  ( n14515 ) ^ ( n14521 )  ;
assign n14523 = ~ ( n7809 ) ;
assign n14524 = ~ ( n6553 ) ;
assign n14525 =  ( n14523 ) | ( n14524 )  ;
assign n14526 =  ( n14522 ) ^ ( n14525 )  ;
assign n14527 =  ( n14526 ) ^ ( n7455 )  ;
assign n14528 =  ( n6825 ) | ( n6834 )  ;
assign n14529 =  ( n14528 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14530 =  ( n14527 ) ^ ( n14529 )  ;
assign n14531 =  ( n6483 ) | ( n6492 )  ;
assign n14532 =  ( n14531 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14533 =  ( n14530 ) ^ ( n14532 )  ;
assign n14534 =  ( n6030 ) | ( n6039 )  ;
assign n14535 =  ( n14534 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14536 =  ( n14533 ) ^ ( n14535 )  ;
assign n14537 =  ( n5802 ) | ( n5811 )  ;
assign n14538 =  ( n14537 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14539 =  ( n14536 ) ^ ( n14538 )  ;
assign n14540 =  ( n5832 ) | ( n5841 )  ;
assign n14541 =  ( n14540 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n14542 =  ( n14539 ) ^ ( n14541 )  ;
assign n14543 =  ( n14542 ) ^ ( n11533 )  ;
assign n14544 = ~ ( n14543 ) ;
assign n14545 =  ( n14489 ) | ( n14544 )  ;
assign n14546 =  ( n5052 ) ^ ( n4889 )  ;
assign n14547 =  ( n14546 ) ^ ( n4561 )  ;
assign n14548 =  ( n14547 ) ^ ( n4571 )  ;
assign n14549 =  ( n14548 ) ^ ( n4274 )  ;
assign n14550 =  ( n14549 ) ^ ( n4290 )  ;
assign n14551 =  ( n14550 ) ^ ( n4307 )  ;
assign n14552 =  ( n14551 ) ^ ( n4324 )  ;
assign n14553 =  ( n14552 ) ^ ( n4353 )  ;
assign n14554 =  ( n14553 ) ^ ( n4602 )  ;
assign n14555 =  ( n14554 ) ^ ( n4590 )  ;
assign n14556 = ~ ( n5182 ) ;
assign n14557 =  ( n5000 ) ^ ( n4784 )  ;
assign n14558 =  ( n14557 ) ^ ( n4800 )  ;
assign n14559 =  ( n14558 ) ^ ( n4817 )  ;
assign n14560 =  ( n14559 ) ^ ( n4834 )  ;
assign n14561 =  ( n14560 ) ^ ( n4862 )  ;
assign n14562 =  ( n14561 ) ^ ( n4859 )  ;
assign n14563 = ~ ( n14562 ) ;
assign n14564 =  ( n14556 ) | ( n14563 )  ;
assign n14565 =  ( n14564 ) | ( n5201 )  ;
assign n14566 = ~ ( n14565 ) ;
assign n14567 =  ( n5248 ) | ( n5341 )  ;
assign n14568 =  ( n14567 ) | ( n10785 )  ;
assign n14569 =  ( n14568 ) | ( n11760 )  ;
assign n14570 =  ( n14569 ) | ( n11801 )  ;
assign n14571 = ~ ( n14570 ) ;
assign n14572 =  ( n5224 ) | ( n14571 )  ;
assign n14573 = ~ ( n14572 ) ;
assign n14574 =  ( n14566 ) | ( n14573 )  ;
assign n14575 =  ( n14555 ) ^ ( n14574 )  ;
assign n14576 = ~ ( n14575 ) ;
assign n14577 = ~ ( n10010 ) ;
assign n14578 = ~ ( n9798 ) ;
assign n14579 =  ( n9804 ) | ( n8179 )  ;
assign n14580 = ~ ( n14579 ) ;
assign n14581 =  ( n14578 ) | ( n14580 )  ;
assign n14582 =  ( n14577 ) ^ ( n14581 )  ;
assign n14583 = ~ ( n7779 ) ;
assign n14584 =  ( n7784 ) | ( n6524 )  ;
assign n14585 = ~ ( n14584 ) ;
assign n14586 =  ( n14583 ) | ( n14585 )  ;
assign n14587 = ~ ( n7801 ) ;
assign n14588 =  ( n14586 ) | ( n14587 )  ;
assign n14589 =  ( n14582 ) ^ ( n14588 )  ;
assign n14590 = ~ ( n7809 ) ;
assign n14591 = ~ ( n6553 ) ;
assign n14592 =  ( n14590 ) | ( n14591 )  ;
assign n14593 =  ( n14589 ) ^ ( n14592 )  ;
assign n14594 =  ( n14593 ) ^ ( n7455 )  ;
assign n14595 =  ( n6825 ) | ( n6834 )  ;
assign n14596 =  ( n14595 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14597 =  ( n14594 ) ^ ( n14596 )  ;
assign n14598 =  ( n6483 ) | ( n6492 )  ;
assign n14599 =  ( n14598 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14600 =  ( n14597 ) ^ ( n14599 )  ;
assign n14601 =  ( n6030 ) | ( n6039 )  ;
assign n14602 =  ( n14601 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14603 =  ( n14600 ) ^ ( n14602 )  ;
assign n14604 =  ( n5802 ) | ( n5811 )  ;
assign n14605 =  ( n14604 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14606 =  ( n14603 ) ^ ( n14605 )  ;
assign n14607 =  ( n14606 ) ^ ( n9471 )  ;
assign n14608 =  ( n14607 ) ^ ( n9468 )  ;
assign n14609 = ~ ( n10140 ) ;
assign n14610 =  ( n14609 ) | ( n10158 )  ;
assign n14611 =  ( n14610 ) | ( n10180 )  ;
assign n14612 = ~ ( n14611 ) ;
assign n14613 = ~ ( n10208 ) ;
assign n14614 = ~ ( n11992 ) ;
assign n14615 =  ( n14613 ) | ( n14614 )  ;
assign n14616 = ~ ( n14615 ) ;
assign n14617 =  ( n14612 ) | ( n14616 )  ;
assign n14618 =  ( n14608 ) ^ ( n14617 )  ;
assign n14619 = ~ ( n14618 ) ;
assign n14620 =  ( n14576 ) | ( n14619 )  ;
assign n14621 = ~ ( n14620 ) ;
assign n14622 =  ( n5052 ) ^ ( n4889 )  ;
assign n14623 =  ( n14622 ) ^ ( n4561 )  ;
assign n14624 =  ( n14623 ) ^ ( n4571 )  ;
assign n14625 =  ( n14624 ) ^ ( n4274 )  ;
assign n14626 =  ( n14625 ) ^ ( n4290 )  ;
assign n14627 =  ( n14626 ) ^ ( n4307 )  ;
assign n14628 =  ( n14627 ) ^ ( n4324 )  ;
assign n14629 =  ( n14628 ) ^ ( n4353 )  ;
assign n14630 =  ( n14629 ) ^ ( n4602 )  ;
assign n14631 =  ( n14630 ) ^ ( n4590 )  ;
assign n14632 =  ( n14566 ) | ( n14573 )  ;
assign n14633 =  ( n14631 ) ^ ( n14632 )  ;
assign n14634 = ~ ( n10010 ) ;
assign n14635 =  ( n14633 ) ^ ( n14634 )  ;
assign n14636 = ~ ( n9798 ) ;
assign n14637 =  ( n9804 ) | ( n8179 )  ;
assign n14638 = ~ ( n14637 ) ;
assign n14639 =  ( n14636 ) | ( n14638 )  ;
assign n14640 =  ( n14635 ) ^ ( n14639 )  ;
assign n14641 = ~ ( n7779 ) ;
assign n14642 =  ( n7784 ) | ( n6524 )  ;
assign n14643 = ~ ( n14642 ) ;
assign n14644 =  ( n14641 ) | ( n14643 )  ;
assign n14645 = ~ ( n7801 ) ;
assign n14646 =  ( n14644 ) | ( n14645 )  ;
assign n14647 =  ( n14640 ) ^ ( n14646 )  ;
assign n14648 = ~ ( n7809 ) ;
assign n14649 = ~ ( n6553 ) ;
assign n14650 =  ( n14648 ) | ( n14649 )  ;
assign n14651 =  ( n14647 ) ^ ( n14650 )  ;
assign n14652 =  ( n14651 ) ^ ( n7455 )  ;
assign n14653 =  ( n6825 ) | ( n6834 )  ;
assign n14654 =  ( n14653 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14655 =  ( n14652 ) ^ ( n14654 )  ;
assign n14656 =  ( n6483 ) | ( n6492 )  ;
assign n14657 =  ( n14656 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14658 =  ( n14655 ) ^ ( n14657 )  ;
assign n14659 =  ( n6030 ) | ( n6039 )  ;
assign n14660 =  ( n14659 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14661 =  ( n14658 ) ^ ( n14660 )  ;
assign n14662 =  ( n5802 ) | ( n5811 )  ;
assign n14663 =  ( n14662 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14664 =  ( n14661 ) ^ ( n14663 )  ;
assign n14665 =  ( n14664 ) ^ ( n9471 )  ;
assign n14666 =  ( n14665 ) ^ ( n9468 )  ;
assign n14667 =  ( n14666 ) ^ ( n14617 )  ;
assign n14668 = ~ ( n14667 ) ;
assign n14669 =  ( n5008 ) | ( n5019 )  ;
assign n14670 =  ( n5214 ) ^ ( n14669 )  ;
assign n14671 =  ( n14670 ) ^ ( n4866 )  ;
assign n14672 =  ( n14671 ) ^ ( n4876 )  ;
assign n14673 =  ( n14672 ) ^ ( n4478 )  ;
assign n14674 =  ( n14673 ) ^ ( n4494 )  ;
assign n14675 =  ( n14674 ) ^ ( n4511 )  ;
assign n14676 =  ( n14675 ) ^ ( n4528 )  ;
assign n14677 =  ( n14676 ) ^ ( n4557 )  ;
assign n14678 =  ( n5248 ) | ( n5341 )  ;
assign n14679 =  ( n14678 ) | ( n10785 )  ;
assign n14680 =  ( n14679 ) | ( n11760 )  ;
assign n14681 =  ( n14680 ) | ( n11801 )  ;
assign n14682 =  ( n14677 ) ^ ( n14681 )  ;
assign n14683 = ~ ( n14682 ) ;
assign n14684 =  ( n14668 ) | ( n14683 )  ;
assign n14685 = ~ ( n10140 ) ;
assign n14686 =  ( n14685 ) | ( n10158 )  ;
assign n14687 = ~ ( n14686 ) ;
assign n14688 = ~ ( n9931 ) ;
assign n14689 =  ( n14688 ) | ( n9952 )  ;
assign n14690 =  ( n14687 ) ^ ( n14689 )  ;
assign n14691 =  ( n14690 ) ^ ( n9792 )  ;
assign n14692 = ~ ( n7809 ) ;
assign n14693 = ~ ( n6553 ) ;
assign n14694 =  ( n14692 ) | ( n14693 )  ;
assign n14695 =  ( n14691 ) ^ ( n14694 )  ;
assign n14696 =  ( n14695 ) ^ ( n7455 )  ;
assign n14697 =  ( n6825 ) | ( n6834 )  ;
assign n14698 =  ( n14697 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14699 =  ( n14696 ) ^ ( n14698 )  ;
assign n14700 =  ( n6483 ) | ( n6492 )  ;
assign n14701 =  ( n14700 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14702 =  ( n14699 ) ^ ( n14701 )  ;
assign n14703 =  ( n6030 ) | ( n6039 )  ;
assign n14704 =  ( n14703 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14705 =  ( n14702 ) ^ ( n14704 )  ;
assign n14706 =  ( n5802 ) | ( n5811 )  ;
assign n14707 =  ( n14706 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14708 =  ( n14705 ) ^ ( n14707 )  ;
assign n14709 =  ( n14708 ) ^ ( n11992 )  ;
assign n14710 = ~ ( n14709 ) ;
assign n14711 =  ( n14684 ) | ( n14710 )  ;
assign n14712 = ~ ( n14711 ) ;
assign n14713 =  ( n14621 ) | ( n14712 )  ;
assign n14714 = ~ ( n14667 ) ;
assign n14715 =  ( n5008 ) | ( n5019 )  ;
assign n14716 =  ( n5214 ) ^ ( n14715 )  ;
assign n14717 =  ( n14716 ) ^ ( n4866 )  ;
assign n14718 =  ( n14717 ) ^ ( n4876 )  ;
assign n14719 =  ( n14718 ) ^ ( n4478 )  ;
assign n14720 =  ( n14719 ) ^ ( n4494 )  ;
assign n14721 =  ( n14720 ) ^ ( n4511 )  ;
assign n14722 =  ( n14721 ) ^ ( n4528 )  ;
assign n14723 =  ( n14722 ) ^ ( n4557 )  ;
assign n14724 =  ( n5248 ) | ( n5341 )  ;
assign n14725 =  ( n14724 ) | ( n10785 )  ;
assign n14726 =  ( n14725 ) | ( n11760 )  ;
assign n14727 =  ( n14726 ) | ( n11801 )  ;
assign n14728 =  ( n14723 ) ^ ( n14727 )  ;
assign n14729 = ~ ( n10140 ) ;
assign n14730 =  ( n14729 ) | ( n10158 )  ;
assign n14731 = ~ ( n14730 ) ;
assign n14732 =  ( n14728 ) ^ ( n14731 )  ;
assign n14733 = ~ ( n9931 ) ;
assign n14734 =  ( n14733 ) | ( n9952 )  ;
assign n14735 =  ( n14732 ) ^ ( n14734 )  ;
assign n14736 =  ( n14735 ) ^ ( n9792 )  ;
assign n14737 = ~ ( n7809 ) ;
assign n14738 = ~ ( n6553 ) ;
assign n14739 =  ( n14737 ) | ( n14738 )  ;
assign n14740 =  ( n14736 ) ^ ( n14739 )  ;
assign n14741 =  ( n14740 ) ^ ( n7455 )  ;
assign n14742 =  ( n6825 ) | ( n6834 )  ;
assign n14743 =  ( n14742 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14744 =  ( n14741 ) ^ ( n14743 )  ;
assign n14745 =  ( n6483 ) | ( n6492 )  ;
assign n14746 =  ( n14745 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14747 =  ( n14744 ) ^ ( n14746 )  ;
assign n14748 =  ( n6030 ) | ( n6039 )  ;
assign n14749 =  ( n14748 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14750 =  ( n14747 ) ^ ( n14749 )  ;
assign n14751 =  ( n5802 ) | ( n5811 )  ;
assign n14752 =  ( n14751 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n14753 =  ( n14750 ) ^ ( n14752 )  ;
assign n14754 =  ( n14753 ) ^ ( n11992 )  ;
assign n14755 = ~ ( n14754 ) ;
assign n14756 =  ( n14714 ) | ( n14755 )  ;
assign n14757 =  ( n5256 ) ^ ( n5182 )  ;
assign n14758 =  ( n14757 ) ^ ( n5000 )  ;
assign n14759 =  ( n14758 ) ^ ( n4784 )  ;
assign n14760 =  ( n14759 ) ^ ( n4800 )  ;
assign n14761 =  ( n14760 ) ^ ( n4817 )  ;
assign n14762 =  ( n14761 ) ^ ( n4834 )  ;
assign n14763 =  ( n14762 ) ^ ( n4862 )  ;
assign n14764 =  ( n14763 ) ^ ( n4859 )  ;
assign n14765 = ~ ( n5325 ) ;
assign n14766 =  ( n5083 ) ^ ( n5099 )  ;
assign n14767 =  ( n14766 ) ^ ( n5116 )  ;
assign n14768 =  ( n14767 ) ^ ( n5141 )  ;
assign n14769 =  ( n14768 ) ^ ( n5129 )  ;
assign n14770 = ~ ( n14769 ) ;
assign n14771 =  ( n14765 ) | ( n14770 )  ;
assign n14772 =  ( n5161 ) ^ ( n5171 )  ;
assign n14773 =  ( n14772 ) ^ ( n4960 )  ;
assign n14774 =  ( n14773 ) ^ ( n4976 )  ;
assign n14775 =  ( n14774 ) ^ ( n4996 )  ;
assign n14776 =  ( n14775 ) ^ ( n5236 )  ;
assign n14777 = ~ ( n14776 ) ;
assign n14778 =  ( n14771 ) | ( n14777 )  ;
assign n14779 = ~ ( n14778 ) ;
assign n14780 =  ( n5366 ) ^ ( n5161 )  ;
assign n14781 =  ( n14780 ) ^ ( n5171 )  ;
assign n14782 =  ( n14781 ) ^ ( n4960 )  ;
assign n14783 =  ( n14782 ) ^ ( n4976 )  ;
assign n14784 =  ( n14783 ) ^ ( n4996 )  ;
assign n14785 =  ( n14784 ) ^ ( n5236 )  ;
assign n14786 = ~ ( n14785 ) ;
assign n14787 =  ( n5446 ) | ( n5473 )  ;
assign n14788 =  ( n14787 ) | ( n5604 )  ;
assign n14789 =  ( n14788 ) | ( n5663 )  ;
assign n14790 = ~ ( n14789 ) ;
assign n14791 =  ( n14786 ) | ( n14790 )  ;
assign n14792 = ~ ( n14791 ) ;
assign n14793 =  ( n14779 ) | ( n14792 )  ;
assign n14794 =  ( n14764 ) ^ ( n14793 )  ;
assign n14795 = ~ ( n14794 ) ;
assign n14796 = ~ ( n10255 ) ;
assign n14797 =  ( n14796 ) ^ ( n10140 )  ;
assign n14798 = ~ ( n7809 ) ;
assign n14799 = ~ ( n9916 ) ;
assign n14800 =  ( n14798 ) | ( n14799 )  ;
assign n14801 =  ( n14797 ) ^ ( n14800 )  ;
assign n14802 =  ( n14801 ) ^ ( n7455 )  ;
assign n14803 =  ( n6825 ) | ( n6834 )  ;
assign n14804 =  ( n14803 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14805 =  ( n14802 ) ^ ( n14804 )  ;
assign n14806 =  ( n6483 ) | ( n6492 )  ;
assign n14807 =  ( n14806 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14808 =  ( n14805 ) ^ ( n14807 )  ;
assign n14809 =  ( n6030 ) | ( n6039 )  ;
assign n14810 =  ( n14809 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14811 =  ( n14808 ) ^ ( n14810 )  ;
assign n14812 =  ( n14811 ) ^ ( n9788 )  ;
assign n14813 =  ( n14812 ) ^ ( n9785 )  ;
assign n14814 = ~ ( n7809 ) ;
assign n14815 = ~ ( n9916 ) ;
assign n14816 =  ( n14814 ) | ( n14815 )  ;
assign n14817 = ~ ( n14816 ) ;
assign n14818 =  ( n14817 ) | ( n10288 )  ;
assign n14819 = ~ ( n10308 ) ;
assign n14820 =  ( n14818 ) | ( n14819 )  ;
assign n14821 = ~ ( n14820 ) ;
assign n14822 = ~ ( n10358 ) ;
assign n14823 = ~ ( n10571 ) ;
assign n14824 =  ( n14822 ) | ( n14823 )  ;
assign n14825 = ~ ( n14824 ) ;
assign n14826 =  ( n14821 ) | ( n14825 )  ;
assign n14827 =  ( n14813 ) ^ ( n14826 )  ;
assign n14828 = ~ ( n14827 ) ;
assign n14829 =  ( n14795 ) | ( n14828 )  ;
assign n14830 = ~ ( n14829 ) ;
assign n14831 =  ( n5256 ) ^ ( n5182 )  ;
assign n14832 =  ( n14831 ) ^ ( n5000 )  ;
assign n14833 =  ( n14832 ) ^ ( n4784 )  ;
assign n14834 =  ( n14833 ) ^ ( n4800 )  ;
assign n14835 =  ( n14834 ) ^ ( n4817 )  ;
assign n14836 =  ( n14835 ) ^ ( n4834 )  ;
assign n14837 =  ( n14836 ) ^ ( n4862 )  ;
assign n14838 =  ( n14837 ) ^ ( n4859 )  ;
assign n14839 =  ( n14779 ) | ( n14792 )  ;
assign n14840 =  ( n14838 ) ^ ( n14839 )  ;
assign n14841 = ~ ( n10255 ) ;
assign n14842 =  ( n14840 ) ^ ( n14841 )  ;
assign n14843 =  ( n14842 ) ^ ( n10140 )  ;
assign n14844 = ~ ( n7809 ) ;
assign n14845 = ~ ( n9916 ) ;
assign n14846 =  ( n14844 ) | ( n14845 )  ;
assign n14847 =  ( n14843 ) ^ ( n14846 )  ;
assign n14848 =  ( n14847 ) ^ ( n7455 )  ;
assign n14849 =  ( n6825 ) | ( n6834 )  ;
assign n14850 =  ( n14849 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14851 =  ( n14848 ) ^ ( n14850 )  ;
assign n14852 =  ( n6483 ) | ( n6492 )  ;
assign n14853 =  ( n14852 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14854 =  ( n14851 ) ^ ( n14853 )  ;
assign n14855 =  ( n6030 ) | ( n6039 )  ;
assign n14856 =  ( n14855 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14857 =  ( n14854 ) ^ ( n14856 )  ;
assign n14858 =  ( n14857 ) ^ ( n9788 )  ;
assign n14859 =  ( n14858 ) ^ ( n9785 )  ;
assign n14860 =  ( n14859 ) ^ ( n14826 )  ;
assign n14861 = ~ ( n14860 ) ;
assign n14862 =  ( n5366 ) ^ ( n5161 )  ;
assign n14863 =  ( n14862 ) ^ ( n5171 )  ;
assign n14864 =  ( n14863 ) ^ ( n4960 )  ;
assign n14865 =  ( n14864 ) ^ ( n4976 )  ;
assign n14866 =  ( n14865 ) ^ ( n4996 )  ;
assign n14867 =  ( n14866 ) ^ ( n5236 )  ;
assign n14868 =  ( n5446 ) | ( n5473 )  ;
assign n14869 =  ( n14868 ) | ( n5604 )  ;
assign n14870 =  ( n14869 ) | ( n5663 )  ;
assign n14871 =  ( n14867 ) ^ ( n14870 )  ;
assign n14872 = ~ ( n14871 ) ;
assign n14873 =  ( n14861 ) | ( n14872 )  ;
assign n14874 = ~ ( n10337 ) ;
assign n14875 = ~ ( n10086 ) ;
assign n14876 =  ( n7784 ) | ( n10091 )  ;
assign n14877 = ~ ( n14876 ) ;
assign n14878 =  ( n14875 ) | ( n14877 )  ;
assign n14879 =  ( n14878 ) | ( n10107 )  ;
assign n14880 =  ( n14874 ) ^ ( n14879 )  ;
assign n14881 = ~ ( n7809 ) ;
assign n14882 = ~ ( n10115 ) ;
assign n14883 =  ( n14881 ) | ( n14882 )  ;
assign n14884 =  ( n14880 ) ^ ( n14883 )  ;
assign n14885 =  ( n14884 ) ^ ( n7455 )  ;
assign n14886 =  ( n6825 ) | ( n6834 )  ;
assign n14887 =  ( n14886 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14888 =  ( n14885 ) ^ ( n14887 )  ;
assign n14889 =  ( n6483 ) | ( n6492 )  ;
assign n14890 =  ( n14889 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14891 =  ( n14888 ) ^ ( n14890 )  ;
assign n14892 =  ( n6030 ) | ( n6039 )  ;
assign n14893 =  ( n14892 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14894 =  ( n14891 ) ^ ( n14893 )  ;
assign n14895 =  ( n14894 ) ^ ( n10571 )  ;
assign n14896 = ~ ( n14895 ) ;
assign n14897 =  ( n14873 ) | ( n14896 )  ;
assign n14898 = ~ ( n14897 ) ;
assign n14899 =  ( n14830 ) | ( n14898 )  ;
assign n14900 = ~ ( n14899 ) ;
assign n14901 =  ( n14756 ) | ( n14900 )  ;
assign n14902 = ~ ( n14901 ) ;
assign n14903 =  ( n14713 ) | ( n14902 )  ;
assign n14904 = ~ ( n14903 ) ;
assign n14905 =  ( n14545 ) | ( n14904 )  ;
assign n14906 = ~ ( n14905 ) ;
assign n14907 =  ( n14484 ) | ( n14906 )  ;
assign n14908 = ~ ( n14169 ) ;
assign n14909 = ~ ( n14288 ) ;
assign n14910 =  ( n14908 ) | ( n14909 )  ;
assign n14911 = ~ ( n14420 ) ;
assign n14912 =  ( n14910 ) | ( n14911 )  ;
assign n14913 = ~ ( n14543 ) ;
assign n14914 =  ( n14912 ) | ( n14913 )  ;
assign n14915 = ~ ( n14667 ) ;
assign n14916 =  ( n14914 ) | ( n14915 )  ;
assign n14917 = ~ ( n14754 ) ;
assign n14918 =  ( n14916 ) | ( n14917 )  ;
assign n14919 =  ( n14918 ) | ( n14861 )  ;
assign n14920 =  ( n5366 ) ^ ( n5161 )  ;
assign n14921 =  ( n14920 ) ^ ( n5171 )  ;
assign n14922 =  ( n14921 ) ^ ( n4960 )  ;
assign n14923 =  ( n14922 ) ^ ( n4976 )  ;
assign n14924 =  ( n14923 ) ^ ( n4996 )  ;
assign n14925 =  ( n14924 ) ^ ( n5236 )  ;
assign n14926 =  ( n5446 ) | ( n5473 )  ;
assign n14927 =  ( n14926 ) | ( n5604 )  ;
assign n14928 =  ( n14927 ) | ( n5663 )  ;
assign n14929 =  ( n14925 ) ^ ( n14928 )  ;
assign n14930 = ~ ( n10337 ) ;
assign n14931 =  ( n14929 ) ^ ( n14930 )  ;
assign n14932 = ~ ( n10086 ) ;
assign n14933 =  ( n7784 ) | ( n10091 )  ;
assign n14934 = ~ ( n14933 ) ;
assign n14935 =  ( n14932 ) | ( n14934 )  ;
assign n14936 =  ( n14935 ) | ( n10107 )  ;
assign n14937 =  ( n14931 ) ^ ( n14936 )  ;
assign n14938 = ~ ( n7809 ) ;
assign n14939 = ~ ( n10115 ) ;
assign n14940 =  ( n14938 ) | ( n14939 )  ;
assign n14941 =  ( n14937 ) ^ ( n14940 )  ;
assign n14942 =  ( n14941 ) ^ ( n7455 )  ;
assign n14943 =  ( n6825 ) | ( n6834 )  ;
assign n14944 =  ( n14943 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14945 =  ( n14942 ) ^ ( n14944 )  ;
assign n14946 =  ( n6483 ) | ( n6492 )  ;
assign n14947 =  ( n14946 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n14948 =  ( n14945 ) ^ ( n14947 )  ;
assign n14949 =  ( n6030 ) | ( n6039 )  ;
assign n14950 =  ( n14949 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n14951 =  ( n14948 ) ^ ( n14950 )  ;
assign n14952 =  ( n14951 ) ^ ( n10571 )  ;
assign n14953 = ~ ( n14952 ) ;
assign n14954 =  ( n14919 ) | ( n14953 )  ;
assign n14955 =  ( n5452 ) ^ ( n5325 )  ;
assign n14956 =  ( n14955 ) ^ ( n5083 )  ;
assign n14957 =  ( n14956 ) ^ ( n5099 )  ;
assign n14958 =  ( n14957 ) ^ ( n5116 )  ;
assign n14959 =  ( n14958 ) ^ ( n5141 )  ;
assign n14960 =  ( n14959 ) ^ ( n5129 )  ;
assign n14961 =  ( n5394 ) ^ ( n5410 )  ;
assign n14962 =  ( n14961 ) ^ ( n5429 )  ;
assign n14963 = ~ ( n14962 ) ;
assign n14964 = ki[5:5] ;
assign n14965 = ~ ( n14964 ) ;
assign n14966 =  ( n14963 ) | ( n14965 )  ;
assign n14967 =  ( n14966 ) | ( n5424 )  ;
assign n14968 =  ( n5433 ) ^ ( n5285 )  ;
assign n14969 =  ( n14968 ) ^ ( n5301 )  ;
assign n14970 =  ( n14969 ) ^ ( n5321 )  ;
assign n14971 = ~ ( n14970 ) ;
assign n14972 =  ( n14967 ) | ( n14971 )  ;
assign n14973 = ~ ( n14972 ) ;
assign n14974 =  ( n5489 ) ^ ( n5433 )  ;
assign n14975 =  ( n14974 ) ^ ( n5285 )  ;
assign n14976 =  ( n14975 ) ^ ( n5301 )  ;
assign n14977 =  ( n14976 ) ^ ( n5321 )  ;
assign n14978 = ~ ( n14977 ) ;
assign n14979 =  ( n5539 ) | ( n5600 )  ;
assign n14980 =  ( n14979 ) | ( n10836 )  ;
assign n14981 = ~ ( n14980 ) ;
assign n14982 =  ( n14978 ) | ( n14981 )  ;
assign n14983 = ~ ( n14982 ) ;
assign n14984 =  ( n14973 ) | ( n14983 )  ;
assign n14985 =  ( n14960 ) ^ ( n14984 )  ;
assign n14986 = ~ ( n14985 ) ;
assign n14987 = ~ ( n10397 ) ;
assign n14988 =  ( n14987 ) | ( n10137 )  ;
assign n14989 = ~ ( n14988 ) ;
assign n14990 = ~ ( n7809 ) ;
assign n14991 = ~ ( n9916 ) ;
assign n14992 =  ( n14990 ) | ( n14991 )  ;
assign n14993 =  ( n14989 ) ^ ( n14992 )  ;
assign n14994 =  ( n14993 ) ^ ( n7455 )  ;
assign n14995 =  ( n6825 ) | ( n6834 )  ;
assign n14996 =  ( n14995 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n14997 =  ( n14994 ) ^ ( n14996 )  ;
assign n14998 =  ( n6483 ) | ( n6492 )  ;
assign n14999 =  ( n14998 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n15000 =  ( n14997 ) ^ ( n14999 )  ;
assign n15001 =  ( n15000 ) ^ ( n10084 )  ;
assign n15002 =  ( n15001 ) ^ ( n10081 )  ;
assign n15003 = kd[5:5] ;
assign n15004 = ~ ( n15003 ) ;
assign n15005 =  ( n10436 ) | ( n15004 )  ;
assign n15006 =  ( n15005 ) | ( n10388 )  ;
assign n15007 =  ( n15006 ) | ( n10449 )  ;
assign n15008 = ~ ( n15007 ) ;
assign n15009 = ~ ( n11086 ) ;
assign n15010 =  ( n10467 ) | ( n15009 )  ;
assign n15011 = ~ ( n15010 ) ;
assign n15012 =  ( n15008 ) | ( n15011 )  ;
assign n15013 =  ( n15002 ) ^ ( n15012 )  ;
assign n15014 = ~ ( n15013 ) ;
assign n15015 =  ( n14986 ) | ( n15014 )  ;
assign n15016 = ~ ( n15015 ) ;
assign n15017 =  ( n5452 ) ^ ( n5325 )  ;
assign n15018 =  ( n15017 ) ^ ( n5083 )  ;
assign n15019 =  ( n15018 ) ^ ( n5099 )  ;
assign n15020 =  ( n15019 ) ^ ( n5116 )  ;
assign n15021 =  ( n15020 ) ^ ( n5141 )  ;
assign n15022 =  ( n15021 ) ^ ( n5129 )  ;
assign n15023 =  ( n14973 ) | ( n14983 )  ;
assign n15024 =  ( n15022 ) ^ ( n15023 )  ;
assign n15025 = ~ ( n10397 ) ;
assign n15026 =  ( n15025 ) | ( n10137 )  ;
assign n15027 = ~ ( n15026 ) ;
assign n15028 =  ( n15024 ) ^ ( n15027 )  ;
assign n15029 = ~ ( n7809 ) ;
assign n15030 = ~ ( n9916 ) ;
assign n15031 =  ( n15029 ) | ( n15030 )  ;
assign n15032 =  ( n15028 ) ^ ( n15031 )  ;
assign n15033 =  ( n15032 ) ^ ( n7455 )  ;
assign n15034 =  ( n6825 ) | ( n6834 )  ;
assign n15035 =  ( n15034 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n15036 =  ( n15033 ) ^ ( n15035 )  ;
assign n15037 =  ( n6483 ) | ( n6492 )  ;
assign n15038 =  ( n15037 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n15039 =  ( n15036 ) ^ ( n15038 )  ;
assign n15040 =  ( n15039 ) ^ ( n10084 )  ;
assign n15041 =  ( n15040 ) ^ ( n10081 )  ;
assign n15042 =  ( n15041 ) ^ ( n15012 )  ;
assign n15043 = ~ ( n15042 ) ;
assign n15044 =  ( n5489 ) ^ ( n5433 )  ;
assign n15045 =  ( n15044 ) ^ ( n5285 )  ;
assign n15046 =  ( n15045 ) ^ ( n5301 )  ;
assign n15047 =  ( n15046 ) ^ ( n5321 )  ;
assign n15048 =  ( n5539 ) | ( n5600 )  ;
assign n15049 =  ( n15048 ) | ( n10836 )  ;
assign n15050 =  ( n15047 ) ^ ( n15049 )  ;
assign n15051 = ~ ( n15050 ) ;
assign n15052 =  ( n15043 ) | ( n15051 )  ;
assign n15053 =  ( n10458 ) ^ ( n10397 )  ;
assign n15054 =  ( n15053 ) ^ ( n7455 )  ;
assign n15055 =  ( n6825 ) | ( n6834 )  ;
assign n15056 =  ( n15055 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n15057 =  ( n15054 ) ^ ( n15056 )  ;
assign n15058 =  ( n6483 ) | ( n6492 )  ;
assign n15059 =  ( n15058 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n15060 =  ( n15057 ) ^ ( n15059 )  ;
assign n15061 =  ( n15060 ) ^ ( n11086 )  ;
assign n15062 = ~ ( n15061 ) ;
assign n15063 =  ( n15052 ) | ( n15062 )  ;
assign n15064 = ~ ( n15063 ) ;
assign n15065 =  ( n15016 ) | ( n15064 )  ;
assign n15066 = ~ ( n15042 ) ;
assign n15067 =  ( n5489 ) ^ ( n5433 )  ;
assign n15068 =  ( n15067 ) ^ ( n5285 )  ;
assign n15069 =  ( n15068 ) ^ ( n5301 )  ;
assign n15070 =  ( n15069 ) ^ ( n5321 )  ;
assign n15071 =  ( n5539 ) | ( n5600 )  ;
assign n15072 =  ( n15071 ) | ( n10836 )  ;
assign n15073 =  ( n15070 ) ^ ( n15072 )  ;
assign n15074 =  ( n15073 ) ^ ( n10458 )  ;
assign n15075 =  ( n15074 ) ^ ( n10397 )  ;
assign n15076 =  ( n15075 ) ^ ( n7455 )  ;
assign n15077 =  ( n6825 ) | ( n6834 )  ;
assign n15078 =  ( n15077 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n15079 =  ( n15076 ) ^ ( n15078 )  ;
assign n15080 =  ( n6483 ) | ( n6492 )  ;
assign n15081 =  ( n15080 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n15082 =  ( n15079 ) ^ ( n15081 )  ;
assign n15083 =  ( n15082 ) ^ ( n11086 )  ;
assign n15084 = ~ ( n15083 ) ;
assign n15085 =  ( n15066 ) | ( n15084 )  ;
assign n15086 = ~ ( n5515 ) ;
assign n15087 = ~ ( n5531 ) ;
assign n15088 =  ( n15086 ) | ( n15087 )  ;
assign n15089 = ~ ( n15088 ) ;
assign n15090 =  ( n15089 ) ^ ( n5394 )  ;
assign n15091 =  ( n15090 ) ^ ( n5410 )  ;
assign n15092 =  ( n15091 ) ^ ( n5429 )  ;
assign n15093 =  ( n15092 ) ^ ( n5426 )  ;
assign n15094 = ~ ( n5594 ) ;
assign n15095 =  ( n5515 ) ^ ( n5531 )  ;
assign n15096 = ~ ( n15095 ) ;
assign n15097 =  ( n15094 ) | ( n15096 )  ;
assign n15098 = ~ ( n15097 ) ;
assign n15099 =  ( n5594 ) ^ ( n5515 )  ;
assign n15100 =  ( n15099 ) ^ ( n5531 )  ;
assign n15101 = ~ ( n15100 ) ;
assign n15102 =  ( n5568 ) ^ ( n5583 )  ;
assign n15103 =  ( n15102 ) ^ ( n5580 )  ;
assign n15104 = ~ ( n15103 ) ;
assign n15105 =  ( n15101 ) | ( n15104 )  ;
assign n15106 = ~ ( n5648 ) ;
assign n15107 =  ( n15105 ) | ( n15106 )  ;
assign n15108 = ~ ( n5657 ) ;
assign n15109 =  ( n15107 ) | ( n15108 )  ;
assign n15110 = ki[1:1] ;
assign n15111 = ~ ( n15110 ) ;
assign n15112 =  ( n15109 ) | ( n15111 )  ;
assign n15113 = ~ ( n15112 ) ;
assign n15114 =  ( n15098 ) | ( n15113 )  ;
assign n15115 =  ( n15093 ) ^ ( n15114 )  ;
assign n15116 = ~ ( n15115 ) ;
assign n15117 = ~ ( n7809 ) ;
assign n15118 =  ( n15117 ) ^ ( n7455 )  ;
assign n15119 =  ( n6825 ) | ( n6834 )  ;
assign n15120 =  ( n15119 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n15121 =  ( n15118 ) ^ ( n15120 )  ;
assign n15122 =  ( n15121 ) ^ ( n10393 )  ;
assign n15123 =  ( n15122 ) ^ ( n10390 )  ;
assign n15124 = ~ ( n10533 ) ;
assign n15125 =  ( n15124 ) | ( n7784 )  ;
assign n15126 = ~ ( n15125 ) ;
assign n15127 =  ( n7455 ) ^ ( n10522 )  ;
assign n15128 =  ( n15127 ) ^ ( n10519 )  ;
assign n15129 = ~ ( n15128 ) ;
assign n15130 =  ( n10550 ) | ( n15129 )  ;
assign n15131 = ~ ( n7455 ) ;
assign n15132 =  ( n15130 ) | ( n15131 )  ;
assign n15133 = ~ ( n10564 ) ;
assign n15134 =  ( n15132 ) | ( n15133 )  ;
assign n15135 = kd[1:1] ;
assign n15136 = ~ ( n15135 ) ;
assign n15137 =  ( n15134 ) | ( n15136 )  ;
assign n15138 = ~ ( n15137 ) ;
assign n15139 =  ( n15126 ) | ( n15138 )  ;
assign n15140 =  ( n15123 ) ^ ( n15139 )  ;
assign n15141 = ~ ( n15140 ) ;
assign n15142 =  ( n15116 ) | ( n15141 )  ;
assign n15143 = ~ ( n15142 ) ;
assign n15144 = ~ ( n5515 ) ;
assign n15145 = ~ ( n5531 ) ;
assign n15146 =  ( n15144 ) | ( n15145 )  ;
assign n15147 = ~ ( n15146 ) ;
assign n15148 =  ( n15147 ) ^ ( n5394 )  ;
assign n15149 =  ( n15148 ) ^ ( n5410 )  ;
assign n15150 =  ( n15149 ) ^ ( n5429 )  ;
assign n15151 =  ( n15150 ) ^ ( n5426 )  ;
assign n15152 =  ( n15098 ) | ( n15113 )  ;
assign n15153 =  ( n15151 ) ^ ( n15152 )  ;
assign n15154 = ~ ( n7809 ) ;
assign n15155 =  ( n15153 ) ^ ( n15154 )  ;
assign n15156 =  ( n15155 ) ^ ( n7455 )  ;
assign n15157 =  ( n6825 ) | ( n6834 )  ;
assign n15158 =  ( n15157 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n15159 =  ( n15156 ) ^ ( n15158 )  ;
assign n15160 =  ( n15159 ) ^ ( n10393 )  ;
assign n15161 =  ( n15160 ) ^ ( n10390 )  ;
assign n15162 =  ( n15161 ) ^ ( n15139 )  ;
assign n15163 = ~ ( n15162 ) ;
assign n15164 =  ( n5594 ) ^ ( n5515 )  ;
assign n15165 =  ( n15164 ) ^ ( n5531 )  ;
assign n15166 =  ( n5568 ) ^ ( n5583 )  ;
assign n15167 =  ( n15166 ) ^ ( n5580 )  ;
assign n15168 = ~ ( n15167 ) ;
assign n15169 = ~ ( n5648 ) ;
assign n15170 =  ( n15168 ) | ( n15169 )  ;
assign n15171 = ~ ( n5657 ) ;
assign n15172 =  ( n15170 ) | ( n15171 )  ;
assign n15173 = ki[1:1] ;
assign n15174 = ~ ( n15173 ) ;
assign n15175 =  ( n15172 ) | ( n15174 )  ;
assign n15176 = ~ ( n15175 ) ;
assign n15177 =  ( n15165 ) ^ ( n15176 )  ;
assign n15178 = ~ ( n15177 ) ;
assign n15179 =  ( n15163 ) | ( n15178 )  ;
assign n15180 =  ( n10533 ) ^ ( n7455 )  ;
assign n15181 =  ( n6825 ) | ( n6834 )  ;
assign n15182 =  ( n15181 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n15183 =  ( n15180 ) ^ ( n15182 )  ;
assign n15184 =  ( n7455 ) ^ ( n10522 )  ;
assign n15185 =  ( n15184 ) ^ ( n10519 )  ;
assign n15186 = ~ ( n15185 ) ;
assign n15187 = ~ ( n7455 ) ;
assign n15188 =  ( n15186 ) | ( n15187 )  ;
assign n15189 = ~ ( n10564 ) ;
assign n15190 =  ( n15188 ) | ( n15189 )  ;
assign n15191 = kd[1:1] ;
assign n15192 = ~ ( n15191 ) ;
assign n15193 =  ( n15190 ) | ( n15192 )  ;
assign n15194 = ~ ( n15193 ) ;
assign n15195 =  ( n15183 ) ^ ( n15194 )  ;
assign n15196 = ~ ( n15195 ) ;
assign n15197 =  ( n15179 ) | ( n15196 )  ;
assign n15198 = ~ ( n15197 ) ;
assign n15199 =  ( n15143 ) | ( n15198 )  ;
assign n15200 = ~ ( n15199 ) ;
assign n15201 =  ( n15085 ) | ( n15200 )  ;
assign n15202 = ~ ( n15201 ) ;
assign n15203 =  ( n15065 ) | ( n15202 )  ;
assign n15204 = ~ ( n15042 ) ;
assign n15205 =  ( n15204 ) | ( n15084 )  ;
assign n15206 = ~ ( n15162 ) ;
assign n15207 =  ( n15205 ) | ( n15206 )  ;
assign n15208 =  ( n5594 ) ^ ( n5515 )  ;
assign n15209 =  ( n15208 ) ^ ( n5531 )  ;
assign n15210 =  ( n15209 ) ^ ( n15176 )  ;
assign n15211 =  ( n15210 ) ^ ( n10533 )  ;
assign n15212 =  ( n15211 ) ^ ( n7455 )  ;
assign n15213 =  ( n6825 ) | ( n6834 )  ;
assign n15214 =  ( n15213 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n15215 =  ( n15212 ) ^ ( n15214 )  ;
assign n15216 =  ( n15215 ) ^ ( n15194 )  ;
assign n15217 = ~ ( n15216 ) ;
assign n15218 =  ( n15207 ) | ( n15217 )  ;
assign n15219 =  ( n5568 ) ^ ( n5583 )  ;
assign n15220 =  ( n15219 ) ^ ( n5580 )  ;
assign n15221 = ~ ( n5648 ) ;
assign n15222 = ~ ( n5657 ) ;
assign n15223 =  ( n15221 ) | ( n15222 )  ;
assign n15224 = ki[1:1] ;
assign n15225 = ~ ( n15224 ) ;
assign n15226 =  ( n15223 ) | ( n15225 )  ;
assign n15227 = ~ ( n15226 ) ;
assign n15228 =  ( n15220 ) ^ ( n15227 )  ;
assign n15229 = ~ ( n15228 ) ;
assign n15230 =  ( n7455 ) ^ ( n10522 )  ;
assign n15231 =  ( n15230 ) ^ ( n10519 )  ;
assign n15232 = ~ ( n7455 ) ;
assign n15233 = ~ ( n10564 ) ;
assign n15234 =  ( n15232 ) | ( n15233 )  ;
assign n15235 = kd[1:1] ;
assign n15236 = ~ ( n15235 ) ;
assign n15237 =  ( n15234 ) | ( n15236 )  ;
assign n15238 = ~ ( n15237 ) ;
assign n15239 =  ( n15231 ) ^ ( n15238 )  ;
assign n15240 = ~ ( n15239 ) ;
assign n15241 =  ( n15229 ) | ( n15240 )  ;
assign n15242 = ~ ( n15241 ) ;
assign n15243 =  ( n5568 ) ^ ( n5583 )  ;
assign n15244 =  ( n15243 ) ^ ( n5580 )  ;
assign n15245 =  ( n15244 ) ^ ( n15227 )  ;
assign n15246 =  ( n15245 ) ^ ( n7455 )  ;
assign n15247 =  ( n15246 ) ^ ( n10522 )  ;
assign n15248 =  ( n15247 ) ^ ( n10519 )  ;
assign n15249 =  ( n15248 ) ^ ( n15238 )  ;
assign n15250 = ~ ( n15249 ) ;
assign n15251 = ~ ( n5657 ) ;
assign n15252 = ki[1:1] ;
assign n15253 = ~ ( n15252 ) ;
assign n15254 =  ( n15251 ) | ( n15253 )  ;
assign n15255 = ~ ( n15254 ) ;
assign n15256 =  ( n5648 ) ^ ( n15255 )  ;
assign n15257 = ~ ( n15256 ) ;
assign n15258 =  ( n15250 ) | ( n15257 )  ;
assign n15259 = ~ ( n10564 ) ;
assign n15260 = kd[1:1] ;
assign n15261 = ~ ( n15260 ) ;
assign n15262 =  ( n15259 ) | ( n15261 )  ;
assign n15263 = ~ ( n15262 ) ;
assign n15264 =  ( n7455 ) ^ ( n15263 )  ;
assign n15265 = ~ ( n15264 ) ;
assign n15266 =  ( n15258 ) | ( n15265 )  ;
assign n15267 = ~ ( n15266 ) ;
assign n15268 =  ( n15242 ) | ( n15267 )  ;
assign n15269 =  ( n5648 ) ^ ( n15255 )  ;
assign n15270 =  ( n15269 ) ^ ( n7455 )  ;
assign n15271 =  ( n15270 ) ^ ( n15263 )  ;
assign n15272 = ~ ( n15271 ) ;
assign n15273 =  ( n15250 ) | ( n15272 )  ;
assign n15274 = ki[1:1] ;
assign n15275 =  ( n5657 ) ^ ( n15274 )  ;
assign n15276 = ~ ( n15275 ) ;
assign n15277 =  ( n15273 ) | ( n15276 )  ;
assign n15278 = kd[1:1] ;
assign n15279 =  ( n10564 ) ^ ( n15278 )  ;
assign n15280 = ~ ( n15279 ) ;
assign n15281 =  ( n15277 ) | ( n15280 )  ;
assign n15282 = ~ ( n15281 ) ;
assign n15283 =  ( n15268 ) | ( n15282 )  ;
assign n15284 = ~ ( n15283 ) ;
assign n15285 =  ( n15218 ) | ( n15284 )  ;
assign n15286 = ~ ( n15285 ) ;
assign n15287 =  ( n15203 ) | ( n15286 )  ;
assign n15288 = ~ ( n15287 ) ;
assign n15289 =  ( n14954 ) | ( n15288 )  ;
assign n15290 = ~ ( n15289 ) ;
assign n15291 =  ( n14907 ) | ( n15290 )  ;
assign n15292 = ~ ( n15291 ) ;
assign n15293 =  ( n14021 ) | ( n15292 )  ;
assign n15294 = ~ ( n15293 ) ;
assign n15295 =  ( n13930 ) | ( n15294 )  ;
assign n15296 =  ( n10581 ) ^ ( n15295 )  ;
assign n15297 =  ( n373 ) | ( n382 )  ;
assign n15298 =  ( n15297 ) ? ( bv_1_0_n2 ) : ( n502 ) ;
assign n15299 = ~ ( n15298 ) ;
assign n15300 =  ( n509 ) ^ ( n15299 )  ;
assign n15301 =  ( n15300 ) ^ ( n10848 )  ;
assign n15302 =  ( n15301 ) ^ ( n5774 )  ;
assign n15303 =  ( n5713 ) | ( n5722 )  ;
assign n15304 =  ( n15303 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n15305 = ~ ( n15304 ) ;
assign n15306 =  ( n15302 ) ^ ( n15305 )  ;
assign n15307 = ~ ( n11094 ) ;
assign n15308 =  ( n5792 ) | ( n15307 )  ;
assign n15309 = ~ ( n15308 ) ;
assign n15310 =  ( n15306 ) ^ ( n15309 )  ;
assign n15311 =  ( bv_1_1_n5 ) ^ ( n488 )  ;
assign n15312 =  ( n15311 ) ^ ( n504 )  ;
assign n15313 =  ( n15312 ) ^ ( n10845 )  ;
assign n15314 = ~ ( n15313 ) ;
assign n15315 =  ( n15314 ) | ( n11130 )  ;
assign n15316 = ~ ( n15315 ) ;
assign n15317 = ~ ( n11340 ) ;
assign n15318 = ~ ( n11541 ) ;
assign n15319 =  ( n15317 ) | ( n15318 )  ;
assign n15320 = ~ ( n15319 ) ;
assign n15321 =  ( n15320 ) | ( n11593 )  ;
assign n15322 = ~ ( n11570 ) ;
assign n15323 =  ( n15322 ) | ( n11619 )  ;
assign n15324 = ~ ( n11810 ) ;
assign n15325 = ~ ( n12000 ) ;
assign n15326 =  ( n15324 ) | ( n15325 )  ;
assign n15327 = ~ ( n15326 ) ;
assign n15328 = ~ ( n12036 ) ;
assign n15329 =  ( n15328 ) | ( n12045 )  ;
assign n15330 =  ( n15329 ) | ( n12063 )  ;
assign n15331 = ~ ( n15330 ) ;
assign n15332 =  ( n15327 ) | ( n15331 )  ;
assign n15333 = ~ ( n15332 ) ;
assign n15334 =  ( n15323 ) | ( n15333 )  ;
assign n15335 = ~ ( n15334 ) ;
assign n15336 =  ( n15321 ) | ( n15335 )  ;
assign n15337 = ~ ( n11570 ) ;
assign n15338 =  ( n15337 ) | ( n11619 )  ;
assign n15339 = ~ ( n12036 ) ;
assign n15340 =  ( n15338 ) | ( n15339 )  ;
assign n15341 =  ( n15340 ) | ( n12090 )  ;
assign n15342 = ~ ( n12184 ) ;
assign n15343 = ~ ( n12301 ) ;
assign n15344 =  ( n15342 ) | ( n15343 )  ;
assign n15345 = ~ ( n15344 ) ;
assign n15346 = ~ ( n12343 ) ;
assign n15347 =  ( n15346 ) | ( n12354 )  ;
assign n15348 =  ( n15347 ) | ( n12376 )  ;
assign n15349 = ~ ( n15348 ) ;
assign n15350 =  ( n15345 ) | ( n15349 )  ;
assign n15351 = ~ ( n12343 ) ;
assign n15352 =  ( n15351 ) | ( n12426 )  ;
assign n15353 = ~ ( n12535 ) ;
assign n15354 = ~ ( n12665 ) ;
assign n15355 =  ( n15353 ) | ( n15354 )  ;
assign n15356 = ~ ( n15355 ) ;
assign n15357 = ~ ( n12722 ) ;
assign n15358 =  ( n15357 ) | ( n12735 )  ;
assign n15359 =  ( n15358 ) | ( n12761 )  ;
assign n15360 = ~ ( n15359 ) ;
assign n15361 =  ( n15356 ) | ( n15360 )  ;
assign n15362 = ~ ( n15361 ) ;
assign n15363 =  ( n15352 ) | ( n15362 )  ;
assign n15364 = ~ ( n15363 ) ;
assign n15365 =  ( n15350 ) | ( n15364 )  ;
assign n15366 = ~ ( n15365 ) ;
assign n15367 =  ( n15341 ) | ( n15366 )  ;
assign n15368 = ~ ( n15367 ) ;
assign n15369 =  ( n15336 ) | ( n15368 )  ;
assign n15370 = ~ ( n11570 ) ;
assign n15371 =  ( n15370 ) | ( n11619 )  ;
assign n15372 = ~ ( n12036 ) ;
assign n15373 =  ( n15371 ) | ( n15372 )  ;
assign n15374 =  ( n15373 ) | ( n12090 )  ;
assign n15375 = ~ ( n12343 ) ;
assign n15376 =  ( n15374 ) | ( n15375 )  ;
assign n15377 =  ( n15376 ) | ( n12426 )  ;
assign n15378 = ~ ( n12722 ) ;
assign n15379 =  ( n15377 ) | ( n15378 )  ;
assign n15380 =  ( n15379 ) | ( n12800 )  ;
assign n15381 = ~ ( n12912 ) ;
assign n15382 = ~ ( n13055 ) ;
assign n15383 =  ( n15381 ) | ( n15382 )  ;
assign n15384 = ~ ( n15383 ) ;
assign n15385 = ~ ( n13119 ) ;
assign n15386 =  ( n15385 ) | ( n13136 )  ;
assign n15387 =  ( n15386 ) | ( n13169 )  ;
assign n15388 = ~ ( n15387 ) ;
assign n15389 =  ( n15384 ) | ( n15388 )  ;
assign n15390 = ~ ( n13119 ) ;
assign n15391 =  ( n15390 ) | ( n13226 )  ;
assign n15392 = ~ ( n13334 ) ;
assign n15393 = ~ ( n13471 ) ;
assign n15394 =  ( n15392 ) | ( n15393 )  ;
assign n15395 = ~ ( n15394 ) ;
assign n15396 = ~ ( n13544 ) ;
assign n15397 =  ( n15396 ) | ( n13568 )  ;
assign n15398 = ~ ( n13613 ) ;
assign n15399 =  ( n15397 ) | ( n15398 )  ;
assign n15400 = ~ ( n15399 ) ;
assign n15401 =  ( n15395 ) | ( n15400 )  ;
assign n15402 = ~ ( n15401 ) ;
assign n15403 =  ( n15391 ) | ( n15402 )  ;
assign n15404 = ~ ( n15403 ) ;
assign n15405 =  ( n15389 ) | ( n15404 )  ;
assign n15406 = ~ ( n13119 ) ;
assign n15407 =  ( n15406 ) | ( n13226 )  ;
assign n15408 = ~ ( n13544 ) ;
assign n15409 =  ( n15407 ) | ( n15408 )  ;
assign n15410 = ~ ( n13683 ) ;
assign n15411 =  ( n15409 ) | ( n15410 )  ;
assign n15412 = ~ ( n13775 ) ;
assign n15413 =  ( n13717 ) | ( n15412 )  ;
assign n15414 = ~ ( n15413 ) ;
assign n15415 = ~ ( n13846 ) ;
assign n15416 =  ( n15415 ) | ( n13867 )  ;
assign n15417 = ~ ( n13914 ) ;
assign n15418 =  ( n15416 ) | ( n15417 )  ;
assign n15419 = ~ ( n15418 ) ;
assign n15420 =  ( n15414 ) | ( n15419 )  ;
assign n15421 = ~ ( n13846 ) ;
assign n15422 = ~ ( n14019 ) ;
assign n15423 =  ( n15421 ) | ( n15422 )  ;
assign n15424 = ~ ( n14106 ) ;
assign n15425 = ~ ( n14169 ) ;
assign n15426 =  ( n15425 ) | ( n14186 )  ;
assign n15427 = ~ ( n14227 ) ;
assign n15428 =  ( n15426 ) | ( n15427 )  ;
assign n15429 = ~ ( n15428 ) ;
assign n15430 =  ( n15424 ) | ( n15429 )  ;
assign n15431 = ~ ( n15430 ) ;
assign n15432 =  ( n15423 ) | ( n15431 )  ;
assign n15433 = ~ ( n15432 ) ;
assign n15434 =  ( n15420 ) | ( n15433 )  ;
assign n15435 = ~ ( n15434 ) ;
assign n15436 =  ( n15411 ) | ( n15435 )  ;
assign n15437 = ~ ( n15436 ) ;
assign n15438 =  ( n15405 ) | ( n15437 )  ;
assign n15439 = ~ ( n15438 ) ;
assign n15440 =  ( n15380 ) | ( n15439 )  ;
assign n15441 = ~ ( n15440 ) ;
assign n15442 =  ( n15369 ) | ( n15441 )  ;
assign n15443 = ~ ( n11570 ) ;
assign n15444 =  ( n15443 ) | ( n11619 )  ;
assign n15445 = ~ ( n12036 ) ;
assign n15446 =  ( n15444 ) | ( n15445 )  ;
assign n15447 =  ( n15446 ) | ( n12090 )  ;
assign n15448 = ~ ( n12343 ) ;
assign n15449 =  ( n15447 ) | ( n15448 )  ;
assign n15450 =  ( n15449 ) | ( n12426 )  ;
assign n15451 = ~ ( n12722 ) ;
assign n15452 =  ( n15450 ) | ( n15451 )  ;
assign n15453 =  ( n15452 ) | ( n12800 )  ;
assign n15454 = ~ ( n13119 ) ;
assign n15455 =  ( n15453 ) | ( n15454 )  ;
assign n15456 =  ( n15455 ) | ( n13226 )  ;
assign n15457 = ~ ( n13544 ) ;
assign n15458 =  ( n15456 ) | ( n15457 )  ;
assign n15459 = ~ ( n13683 ) ;
assign n15460 =  ( n15458 ) | ( n15459 )  ;
assign n15461 = ~ ( n13846 ) ;
assign n15462 =  ( n15460 ) | ( n15461 )  ;
assign n15463 = ~ ( n14019 ) ;
assign n15464 =  ( n15462 ) | ( n15463 )  ;
assign n15465 = ~ ( n14169 ) ;
assign n15466 =  ( n15464 ) | ( n15465 )  ;
assign n15467 = ~ ( n14288 ) ;
assign n15468 =  ( n15466 ) | ( n15467 )  ;
assign n15469 = ~ ( n14321 ) ;
assign n15470 = ~ ( n14365 ) ;
assign n15471 =  ( n15469 ) | ( n15470 )  ;
assign n15472 = ~ ( n15471 ) ;
assign n15473 = ~ ( n14420 ) ;
assign n15474 = ~ ( n14441 ) ;
assign n15475 =  ( n15473 ) | ( n15474 )  ;
assign n15476 = ~ ( n14476 ) ;
assign n15477 =  ( n15475 ) | ( n15476 )  ;
assign n15478 = ~ ( n15477 ) ;
assign n15479 =  ( n15472 ) | ( n15478 )  ;
assign n15480 = ~ ( n14420 ) ;
assign n15481 = ~ ( n14543 ) ;
assign n15482 =  ( n15480 ) | ( n15481 )  ;
assign n15483 = ~ ( n14620 ) ;
assign n15484 = ~ ( n14667 ) ;
assign n15485 =  ( n15484 ) | ( n14683 )  ;
assign n15486 = ~ ( n14709 ) ;
assign n15487 =  ( n15485 ) | ( n15486 )  ;
assign n15488 = ~ ( n15487 ) ;
assign n15489 =  ( n15483 ) | ( n15488 )  ;
assign n15490 = ~ ( n15489 ) ;
assign n15491 =  ( n15482 ) | ( n15490 )  ;
assign n15492 = ~ ( n15491 ) ;
assign n15493 =  ( n15479 ) | ( n15492 )  ;
assign n15494 = ~ ( n14420 ) ;
assign n15495 = ~ ( n14543 ) ;
assign n15496 =  ( n15494 ) | ( n15495 )  ;
assign n15497 = ~ ( n14667 ) ;
assign n15498 =  ( n15496 ) | ( n15497 )  ;
assign n15499 = ~ ( n14754 ) ;
assign n15500 =  ( n15498 ) | ( n15499 )  ;
assign n15501 = ~ ( n14829 ) ;
assign n15502 =  ( n14861 ) | ( n14872 )  ;
assign n15503 = ~ ( n14895 ) ;
assign n15504 =  ( n15502 ) | ( n15503 )  ;
assign n15505 = ~ ( n15504 ) ;
assign n15506 =  ( n15501 ) | ( n15505 )  ;
assign n15507 = ~ ( n14952 ) ;
assign n15508 =  ( n14861 ) | ( n15507 )  ;
assign n15509 = ~ ( n15015 ) ;
assign n15510 = ~ ( n15042 ) ;
assign n15511 =  ( n15510 ) | ( n15051 )  ;
assign n15512 =  ( n15511 ) | ( n15062 )  ;
assign n15513 = ~ ( n15512 ) ;
assign n15514 =  ( n15509 ) | ( n15513 )  ;
assign n15515 = ~ ( n15514 ) ;
assign n15516 =  ( n15508 ) | ( n15515 )  ;
assign n15517 = ~ ( n15516 ) ;
assign n15518 =  ( n15506 ) | ( n15517 )  ;
assign n15519 = ~ ( n15518 ) ;
assign n15520 =  ( n15500 ) | ( n15519 )  ;
assign n15521 = ~ ( n15520 ) ;
assign n15522 =  ( n15493 ) | ( n15521 )  ;
assign n15523 = ~ ( n14420 ) ;
assign n15524 = ~ ( n14543 ) ;
assign n15525 =  ( n15523 ) | ( n15524 )  ;
assign n15526 = ~ ( n14667 ) ;
assign n15527 =  ( n15525 ) | ( n15526 )  ;
assign n15528 = ~ ( n14754 ) ;
assign n15529 =  ( n15527 ) | ( n15528 )  ;
assign n15530 =  ( n15529 ) | ( n14861 )  ;
assign n15531 = ~ ( n14952 ) ;
assign n15532 =  ( n15530 ) | ( n15531 )  ;
assign n15533 = ~ ( n15042 ) ;
assign n15534 =  ( n15532 ) | ( n15533 )  ;
assign n15535 =  ( n15534 ) | ( n15084 )  ;
assign n15536 = ~ ( n15115 ) ;
assign n15537 =  ( n15536 ) | ( n15141 )  ;
assign n15538 = ~ ( n15537 ) ;
assign n15539 =  ( n15538 ) | ( n15198 )  ;
assign n15540 = ~ ( n15162 ) ;
assign n15541 =  ( n15540 ) | ( n15217 )  ;
assign n15542 =  ( n15242 ) | ( n15267 )  ;
assign n15543 = ~ ( n15542 ) ;
assign n15544 =  ( n15541 ) | ( n15543 )  ;
assign n15545 = ~ ( n15544 ) ;
assign n15546 =  ( n15539 ) | ( n15545 )  ;
assign n15547 = ~ ( n15162 ) ;
assign n15548 =  ( n15547 ) | ( n15217 )  ;
assign n15549 =  ( n15548 ) | ( n15250 )  ;
assign n15550 =  ( n5648 ) ^ ( n15255 )  ;
assign n15551 =  ( n15550 ) ^ ( n7455 )  ;
assign n15552 =  ( n15551 ) ^ ( n15263 )  ;
assign n15553 = ~ ( n15552 ) ;
assign n15554 =  ( n15549 ) | ( n15553 )  ;
assign n15555 = ki[1:1] ;
assign n15556 =  ( n5657 ) ^ ( n15555 )  ;
assign n15557 = ~ ( n15556 ) ;
assign n15558 =  ( n15554 ) | ( n15557 )  ;
assign n15559 = kd[1:1] ;
assign n15560 =  ( n10564 ) ^ ( n15559 )  ;
assign n15561 = ~ ( n15560 ) ;
assign n15562 =  ( n15558 ) | ( n15561 )  ;
assign n15563 = ~ ( n15562 ) ;
assign n15564 =  ( n15546 ) | ( n15563 )  ;
assign n15565 = ~ ( n15564 ) ;
assign n15566 =  ( n15535 ) | ( n15565 )  ;
assign n15567 = ~ ( n15566 ) ;
assign n15568 =  ( n15522 ) | ( n15567 )  ;
assign n15569 = ~ ( n15568 ) ;
assign n15570 =  ( n15468 ) | ( n15569 )  ;
assign n15571 = ~ ( n15570 ) ;
assign n15572 =  ( n15442 ) | ( n15571 )  ;
assign n15573 = ~ ( n15572 ) ;
assign n15574 =  ( n11145 ) | ( n15573 )  ;
assign n15575 = ~ ( n15574 ) ;
assign n15576 =  ( n15316 ) | ( n15575 )  ;
assign n15577 =  ( n15310 ) ^ ( n15576 )  ;
assign n15578 =  { ( n15296 ) , ( n15577 ) }  ;
assign n15579 =  ( n488 ) ^ ( n504 )  ;
assign n15580 =  ( n15579 ) ^ ( n10845 )  ;
assign n15581 = ~ ( n5747 ) ;
assign n15582 = ~ ( n5759 ) ;
assign n15583 =  ( n15581 ) | ( n15582 )  ;
assign n15584 =  ( n15580 ) ^ ( n15583 )  ;
assign n15585 =  ( n5713 ) | ( n5722 )  ;
assign n15586 =  ( n15585 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n15587 =  ( n15584 ) ^ ( n15586 )  ;
assign n15588 =  ( n15587 ) ^ ( n11094 )  ;
assign n15589 =  ( n15588 ) ^ ( n15572 )  ;
assign n15590 =  { ( n15578 ) , ( n15589 ) }  ;
assign n15591 =  ( n834 ) ^ ( n459 )  ;
assign n15592 =  ( n30 ) | ( n39 )  ;
assign n15593 =  ( n15592 ) ? ( bv_1_0_n2 ) : ( n342 ) ;
assign n15594 = ~ ( n15593 ) ;
assign n15595 =  ( n15591 ) ^ ( n15594 )  ;
assign n15596 =  ( n15595 ) ^ ( n484 )  ;
assign n15597 =  ( n15596 ) ^ ( n11339 )  ;
assign n15598 = ~ ( n5959 ) ;
assign n15599 =  ( n5965 ) | ( n5972 )  ;
assign n15600 = ~ ( n15599 ) ;
assign n15601 =  ( n15598 ) | ( n15600 )  ;
assign n15602 =  ( n15597 ) ^ ( n15601 )  ;
assign n15603 = ~ ( n5736 ) ;
assign n15604 =  ( n15603 ) | ( n5742 )  ;
assign n15605 =  ( n15602 ) ^ ( n15604 )  ;
assign n15606 =  ( n5682 ) | ( n5691 )  ;
assign n15607 =  ( n15606 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n15608 = ~ ( n15607 ) ;
assign n15609 =  ( n15605 ) ^ ( n15608 )  ;
assign n15610 =  ( n5713 ) | ( n5722 )  ;
assign n15611 =  ( n15610 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n15612 =  ( n15609 ) ^ ( n15611 )  ;
assign n15613 = ~ ( n11537 ) ;
assign n15614 =  ( n6020 ) | ( n15613 )  ;
assign n15615 = ~ ( n15614 ) ;
assign n15616 =  ( n15612 ) ^ ( n15615 )  ;
assign n15617 =  ( bv_1_1_n5 ) ^ ( n808 )  ;
assign n15618 =  ( n15617 ) ^ ( n823 )  ;
assign n15619 =  ( n15618 ) ^ ( n344 )  ;
assign n15620 =  ( n15619 ) ^ ( n454 )  ;
assign n15621 =  ( n15620 ) ^ ( n11336 )  ;
assign n15622 = ~ ( n15621 ) ;
assign n15623 =  ( n15622 ) | ( n11591 )  ;
assign n15624 = ~ ( n15623 ) ;
assign n15625 = ~ ( n11810 ) ;
assign n15626 = ~ ( n12000 ) ;
assign n15627 =  ( n15625 ) | ( n15626 )  ;
assign n15628 = ~ ( n15627 ) ;
assign n15629 = ~ ( n12036 ) ;
assign n15630 =  ( n15629 ) | ( n12045 )  ;
assign n15631 =  ( n15630 ) | ( n12063 )  ;
assign n15632 = ~ ( n15631 ) ;
assign n15633 =  ( n15628 ) | ( n15632 )  ;
assign n15634 = ~ ( n12036 ) ;
assign n15635 =  ( n15634 ) | ( n12090 )  ;
assign n15636 = ~ ( n12379 ) ;
assign n15637 =  ( n15635 ) | ( n15636 )  ;
assign n15638 = ~ ( n15637 ) ;
assign n15639 =  ( n15633 ) | ( n15638 )  ;
assign n15640 = ~ ( n12036 ) ;
assign n15641 =  ( n15640 ) | ( n12090 )  ;
assign n15642 = ~ ( n12343 ) ;
assign n15643 =  ( n15641 ) | ( n15642 )  ;
assign n15644 =  ( n15643 ) | ( n12426 )  ;
assign n15645 = ~ ( n12535 ) ;
assign n15646 = ~ ( n12665 ) ;
assign n15647 =  ( n15645 ) | ( n15646 )  ;
assign n15648 = ~ ( n15647 ) ;
assign n15649 = ~ ( n12722 ) ;
assign n15650 =  ( n15649 ) | ( n12735 )  ;
assign n15651 =  ( n15650 ) | ( n12761 )  ;
assign n15652 = ~ ( n15651 ) ;
assign n15653 =  ( n15648 ) | ( n15652 )  ;
assign n15654 = ~ ( n12722 ) ;
assign n15655 =  ( n15654 ) | ( n12800 )  ;
assign n15656 = ~ ( n13172 ) ;
assign n15657 =  ( n15655 ) | ( n15656 )  ;
assign n15658 = ~ ( n15657 ) ;
assign n15659 =  ( n15653 ) | ( n15658 )  ;
assign n15660 = ~ ( n15659 ) ;
assign n15661 =  ( n15644 ) | ( n15660 )  ;
assign n15662 = ~ ( n15661 ) ;
assign n15663 =  ( n15639 ) | ( n15662 )  ;
assign n15664 = ~ ( n12036 ) ;
assign n15665 =  ( n15664 ) | ( n12090 )  ;
assign n15666 = ~ ( n12343 ) ;
assign n15667 =  ( n15665 ) | ( n15666 )  ;
assign n15668 =  ( n15667 ) | ( n12426 )  ;
assign n15669 = ~ ( n12722 ) ;
assign n15670 =  ( n15668 ) | ( n15669 )  ;
assign n15671 =  ( n15670 ) | ( n12800 )  ;
assign n15672 = ~ ( n13119 ) ;
assign n15673 =  ( n15671 ) | ( n15672 )  ;
assign n15674 =  ( n15673 ) | ( n13226 )  ;
assign n15675 = ~ ( n13334 ) ;
assign n15676 = ~ ( n13471 ) ;
assign n15677 =  ( n15675 ) | ( n15676 )  ;
assign n15678 = ~ ( n15677 ) ;
assign n15679 = ~ ( n13544 ) ;
assign n15680 =  ( n15679 ) | ( n13568 )  ;
assign n15681 = ~ ( n13613 ) ;
assign n15682 =  ( n15680 ) | ( n15681 )  ;
assign n15683 = ~ ( n15682 ) ;
assign n15684 =  ( n15678 ) | ( n15683 )  ;
assign n15685 = ~ ( n13544 ) ;
assign n15686 = ~ ( n13683 ) ;
assign n15687 =  ( n15685 ) | ( n15686 )  ;
assign n15688 = ~ ( n13918 ) ;
assign n15689 =  ( n15687 ) | ( n15688 )  ;
assign n15690 = ~ ( n15689 ) ;
assign n15691 =  ( n15684 ) | ( n15690 )  ;
assign n15692 = ~ ( n13544 ) ;
assign n15693 = ~ ( n13683 ) ;
assign n15694 =  ( n15692 ) | ( n15693 )  ;
assign n15695 = ~ ( n13846 ) ;
assign n15696 =  ( n15694 ) | ( n15695 )  ;
assign n15697 = ~ ( n14019 ) ;
assign n15698 =  ( n15696 ) | ( n15697 )  ;
assign n15699 = ~ ( n14106 ) ;
assign n15700 = ~ ( n14169 ) ;
assign n15701 =  ( n15700 ) | ( n14186 )  ;
assign n15702 = ~ ( n14227 ) ;
assign n15703 =  ( n15701 ) | ( n15702 )  ;
assign n15704 = ~ ( n15703 ) ;
assign n15705 =  ( n15699 ) | ( n15704 )  ;
assign n15706 = ~ ( n14169 ) ;
assign n15707 = ~ ( n14288 ) ;
assign n15708 =  ( n15706 ) | ( n15707 )  ;
assign n15709 = ~ ( n14480 ) ;
assign n15710 =  ( n15708 ) | ( n15709 )  ;
assign n15711 = ~ ( n15710 ) ;
assign n15712 =  ( n15705 ) | ( n15711 )  ;
assign n15713 = ~ ( n15712 ) ;
assign n15714 =  ( n15698 ) | ( n15713 )  ;
assign n15715 = ~ ( n15714 ) ;
assign n15716 =  ( n15691 ) | ( n15715 )  ;
assign n15717 = ~ ( n15716 ) ;
assign n15718 =  ( n15674 ) | ( n15717 )  ;
assign n15719 = ~ ( n15718 ) ;
assign n15720 =  ( n15663 ) | ( n15719 )  ;
assign n15721 = ~ ( n12036 ) ;
assign n15722 =  ( n15721 ) | ( n12090 )  ;
assign n15723 = ~ ( n12343 ) ;
assign n15724 =  ( n15722 ) | ( n15723 )  ;
assign n15725 =  ( n15724 ) | ( n12426 )  ;
assign n15726 = ~ ( n12722 ) ;
assign n15727 =  ( n15725 ) | ( n15726 )  ;
assign n15728 =  ( n15727 ) | ( n12800 )  ;
assign n15729 = ~ ( n13119 ) ;
assign n15730 =  ( n15728 ) | ( n15729 )  ;
assign n15731 =  ( n15730 ) | ( n13226 )  ;
assign n15732 = ~ ( n13544 ) ;
assign n15733 =  ( n15731 ) | ( n15732 )  ;
assign n15734 = ~ ( n13683 ) ;
assign n15735 =  ( n15733 ) | ( n15734 )  ;
assign n15736 = ~ ( n13846 ) ;
assign n15737 =  ( n15735 ) | ( n15736 )  ;
assign n15738 = ~ ( n14019 ) ;
assign n15739 =  ( n15737 ) | ( n15738 )  ;
assign n15740 = ~ ( n14169 ) ;
assign n15741 =  ( n15739 ) | ( n15740 )  ;
assign n15742 = ~ ( n14288 ) ;
assign n15743 =  ( n15741 ) | ( n15742 )  ;
assign n15744 = ~ ( n14420 ) ;
assign n15745 =  ( n15743 ) | ( n15744 )  ;
assign n15746 = ~ ( n14543 ) ;
assign n15747 =  ( n15745 ) | ( n15746 )  ;
assign n15748 = ~ ( n14620 ) ;
assign n15749 = ~ ( n14667 ) ;
assign n15750 =  ( n15749 ) | ( n14683 )  ;
assign n15751 = ~ ( n14709 ) ;
assign n15752 =  ( n15750 ) | ( n15751 )  ;
assign n15753 = ~ ( n15752 ) ;
assign n15754 =  ( n15748 ) | ( n15753 )  ;
assign n15755 = ~ ( n14667 ) ;
assign n15756 = ~ ( n14754 ) ;
assign n15757 =  ( n15755 ) | ( n15756 )  ;
assign n15758 = ~ ( n14899 ) ;
assign n15759 =  ( n15757 ) | ( n15758 )  ;
assign n15760 = ~ ( n15759 ) ;
assign n15761 =  ( n15754 ) | ( n15760 )  ;
assign n15762 = ~ ( n14667 ) ;
assign n15763 = ~ ( n14754 ) ;
assign n15764 =  ( n15762 ) | ( n15763 )  ;
assign n15765 =  ( n15764 ) | ( n14861 )  ;
assign n15766 = ~ ( n14952 ) ;
assign n15767 =  ( n15765 ) | ( n15766 )  ;
assign n15768 = ~ ( n15015 ) ;
assign n15769 = ~ ( n15042 ) ;
assign n15770 =  ( n15769 ) | ( n15051 )  ;
assign n15771 =  ( n15770 ) | ( n15062 )  ;
assign n15772 = ~ ( n15771 ) ;
assign n15773 =  ( n15768 ) | ( n15772 )  ;
assign n15774 = ~ ( n15042 ) ;
assign n15775 =  ( n15774 ) | ( n15084 )  ;
assign n15776 = ~ ( n15199 ) ;
assign n15777 =  ( n15775 ) | ( n15776 )  ;
assign n15778 = ~ ( n15777 ) ;
assign n15779 =  ( n15773 ) | ( n15778 )  ;
assign n15780 = ~ ( n15779 ) ;
assign n15781 =  ( n15767 ) | ( n15780 )  ;
assign n15782 = ~ ( n15781 ) ;
assign n15783 =  ( n15761 ) | ( n15782 )  ;
assign n15784 = ~ ( n14667 ) ;
assign n15785 = ~ ( n14754 ) ;
assign n15786 =  ( n15784 ) | ( n15785 )  ;
assign n15787 =  ( n15786 ) | ( n14861 )  ;
assign n15788 = ~ ( n14952 ) ;
assign n15789 =  ( n15787 ) | ( n15788 )  ;
assign n15790 = ~ ( n15042 ) ;
assign n15791 =  ( n15789 ) | ( n15790 )  ;
assign n15792 =  ( n15791 ) | ( n15084 )  ;
assign n15793 = ~ ( n15162 ) ;
assign n15794 =  ( n15792 ) | ( n15793 )  ;
assign n15795 =  ( n15794 ) | ( n15217 )  ;
assign n15796 =  ( n15242 ) | ( n15267 )  ;
assign n15797 = ~ ( n15281 ) ;
assign n15798 =  ( n15796 ) | ( n15797 )  ;
assign n15799 = ~ ( n15798 ) ;
assign n15800 =  ( n15795 ) | ( n15799 )  ;
assign n15801 = ~ ( n15800 ) ;
assign n15802 =  ( n15783 ) | ( n15801 )  ;
assign n15803 = ~ ( n15802 ) ;
assign n15804 =  ( n15747 ) | ( n15803 )  ;
assign n15805 = ~ ( n15804 ) ;
assign n15806 =  ( n15720 ) | ( n15805 )  ;
assign n15807 = ~ ( n15806 ) ;
assign n15808 =  ( n11619 ) | ( n15807 )  ;
assign n15809 = ~ ( n15808 ) ;
assign n15810 =  ( n15624 ) | ( n15809 )  ;
assign n15811 =  ( n15616 ) ^ ( n15810 )  ;
assign n15812 =  { ( n15590 ) , ( n15811 ) }  ;
assign n15813 =  ( n808 ) ^ ( n823 )  ;
assign n15814 =  ( n15813 ) ^ ( n344 )  ;
assign n15815 =  ( n15814 ) ^ ( n454 )  ;
assign n15816 =  ( n15815 ) ^ ( n11336 )  ;
assign n15817 =  ( n15816 ) ^ ( n5936 )  ;
assign n15818 = ~ ( n5943 ) ;
assign n15819 = ~ ( n5955 ) ;
assign n15820 =  ( n15818 ) | ( n15819 )  ;
assign n15821 =  ( n15817 ) ^ ( n15820 )  ;
assign n15822 =  ( n5682 ) | ( n5691 )  ;
assign n15823 =  ( n15822 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n15824 =  ( n15821 ) ^ ( n15823 )  ;
assign n15825 =  ( n5713 ) | ( n5722 )  ;
assign n15826 =  ( n15825 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n15827 =  ( n15824 ) ^ ( n15826 )  ;
assign n15828 =  ( n15827 ) ^ ( n11537 )  ;
assign n15829 =  ( n15828 ) ^ ( n15806 )  ;
assign n15830 =  { ( n15812 ) , ( n15829 ) }  ;
assign n15831 =  ( n666 ) ^ ( n682 )  ;
assign n15832 =  ( n15831 ) ^ ( n697 )  ;
assign n15833 =  ( n15832 ) ^ ( n759 )  ;
assign n15834 =  ( n763 ) | ( n15833 )  ;
assign n15835 =  ( n1212 ) ^ ( n15834 )  ;
assign n15836 =  ( n15835 ) ^ ( n778 )  ;
assign n15837 =  ( n586 ) | ( n595 )  ;
assign n15838 =  ( n15837 ) ? ( bv_1_0_n2 ) : ( n680 ) ;
assign n15839 = ~ ( n15838 ) ;
assign n15840 =  ( n15836 ) ^ ( n15839 )  ;
assign n15841 =  ( n15840 ) ^ ( n796 )  ;
assign n15842 =  ( n15841 ) ^ ( n803 )  ;
assign n15843 =  ( n15842 ) ^ ( n11809 )  ;
assign n15844 =  ( n15843 ) ^ ( n6264 )  ;
assign n15845 =  ( n15844 ) ^ ( n5894 )  ;
assign n15846 = ~ ( n5902 ) ;
assign n15847 = ~ ( n5913 ) ;
assign n15848 =  ( n15846 ) | ( n15847 )  ;
assign n15849 =  ( n15845 ) ^ ( n15848 )  ;
assign n15850 =  ( n5832 ) | ( n5841 )  ;
assign n15851 =  ( n15850 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n15852 = ~ ( n15851 ) ;
assign n15853 =  ( n15849 ) ^ ( n15852 )  ;
assign n15854 =  ( n5682 ) | ( n5691 )  ;
assign n15855 =  ( n15854 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n15856 =  ( n15853 ) ^ ( n15855 )  ;
assign n15857 =  ( n5713 ) | ( n5722 )  ;
assign n15858 =  ( n15857 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n15859 =  ( n15856 ) ^ ( n15858 )  ;
assign n15860 = ~ ( n11996 ) ;
assign n15861 =  ( n6314 ) | ( n15860 )  ;
assign n15862 = ~ ( n15861 ) ;
assign n15863 =  ( n15859 ) ^ ( n15862 )  ;
assign n15864 =  ( n12045 ) | ( n12063 )  ;
assign n15865 = ~ ( n15864 ) ;
assign n15866 = ~ ( n12184 ) ;
assign n15867 = ~ ( n12301 ) ;
assign n15868 =  ( n15866 ) | ( n15867 )  ;
assign n15869 = ~ ( n15868 ) ;
assign n15870 = ~ ( n12343 ) ;
assign n15871 =  ( n15870 ) | ( n12354 )  ;
assign n15872 =  ( n15871 ) | ( n12376 )  ;
assign n15873 = ~ ( n15872 ) ;
assign n15874 =  ( n15869 ) | ( n15873 )  ;
assign n15875 = ~ ( n12343 ) ;
assign n15876 =  ( n15875 ) | ( n12426 )  ;
assign n15877 = ~ ( n15361 ) ;
assign n15878 =  ( n15876 ) | ( n15877 )  ;
assign n15879 = ~ ( n15878 ) ;
assign n15880 =  ( n15874 ) | ( n15879 )  ;
assign n15881 = ~ ( n12343 ) ;
assign n15882 =  ( n15881 ) | ( n12426 )  ;
assign n15883 = ~ ( n12722 ) ;
assign n15884 =  ( n15882 ) | ( n15883 )  ;
assign n15885 =  ( n15884 ) | ( n12800 )  ;
assign n15886 = ~ ( n12912 ) ;
assign n15887 = ~ ( n13055 ) ;
assign n15888 =  ( n15886 ) | ( n15887 )  ;
assign n15889 = ~ ( n15888 ) ;
assign n15890 = ~ ( n13119 ) ;
assign n15891 =  ( n15890 ) | ( n13136 )  ;
assign n15892 =  ( n15891 ) | ( n13169 )  ;
assign n15893 = ~ ( n15892 ) ;
assign n15894 =  ( n15889 ) | ( n15893 )  ;
assign n15895 = ~ ( n13119 ) ;
assign n15896 =  ( n15895 ) | ( n13226 )  ;
assign n15897 = ~ ( n15401 ) ;
assign n15898 =  ( n15896 ) | ( n15897 )  ;
assign n15899 = ~ ( n15898 ) ;
assign n15900 =  ( n15894 ) | ( n15899 )  ;
assign n15901 = ~ ( n15900 ) ;
assign n15902 =  ( n15885 ) | ( n15901 )  ;
assign n15903 = ~ ( n15902 ) ;
assign n15904 =  ( n15880 ) | ( n15903 )  ;
assign n15905 = ~ ( n12343 ) ;
assign n15906 =  ( n15905 ) | ( n12426 )  ;
assign n15907 = ~ ( n12722 ) ;
assign n15908 =  ( n15906 ) | ( n15907 )  ;
assign n15909 =  ( n15908 ) | ( n12800 )  ;
assign n15910 = ~ ( n13119 ) ;
assign n15911 =  ( n15909 ) | ( n15910 )  ;
assign n15912 =  ( n15911 ) | ( n13226 )  ;
assign n15913 = ~ ( n13544 ) ;
assign n15914 =  ( n15912 ) | ( n15913 )  ;
assign n15915 = ~ ( n13683 ) ;
assign n15916 =  ( n15914 ) | ( n15915 )  ;
assign n15917 = ~ ( n13775 ) ;
assign n15918 =  ( n13717 ) | ( n15917 )  ;
assign n15919 = ~ ( n15918 ) ;
assign n15920 = ~ ( n13846 ) ;
assign n15921 =  ( n15920 ) | ( n13867 )  ;
assign n15922 = ~ ( n13914 ) ;
assign n15923 =  ( n15921 ) | ( n15922 )  ;
assign n15924 = ~ ( n15923 ) ;
assign n15925 =  ( n15919 ) | ( n15924 )  ;
assign n15926 = ~ ( n13846 ) ;
assign n15927 = ~ ( n14019 ) ;
assign n15928 =  ( n15926 ) | ( n15927 )  ;
assign n15929 = ~ ( n15430 ) ;
assign n15930 =  ( n15928 ) | ( n15929 )  ;
assign n15931 = ~ ( n15930 ) ;
assign n15932 =  ( n15925 ) | ( n15931 )  ;
assign n15933 = ~ ( n13846 ) ;
assign n15934 = ~ ( n14019 ) ;
assign n15935 =  ( n15933 ) | ( n15934 )  ;
assign n15936 = ~ ( n14169 ) ;
assign n15937 =  ( n15935 ) | ( n15936 )  ;
assign n15938 = ~ ( n14288 ) ;
assign n15939 =  ( n15937 ) | ( n15938 )  ;
assign n15940 = ~ ( n14321 ) ;
assign n15941 = ~ ( n14365 ) ;
assign n15942 =  ( n15940 ) | ( n15941 )  ;
assign n15943 = ~ ( n15942 ) ;
assign n15944 = ~ ( n14420 ) ;
assign n15945 = ~ ( n14441 ) ;
assign n15946 =  ( n15944 ) | ( n15945 )  ;
assign n15947 = ~ ( n14476 ) ;
assign n15948 =  ( n15946 ) | ( n15947 )  ;
assign n15949 = ~ ( n15948 ) ;
assign n15950 =  ( n15943 ) | ( n15949 )  ;
assign n15951 = ~ ( n14420 ) ;
assign n15952 = ~ ( n14543 ) ;
assign n15953 =  ( n15951 ) | ( n15952 )  ;
assign n15954 = ~ ( n15489 ) ;
assign n15955 =  ( n15953 ) | ( n15954 )  ;
assign n15956 = ~ ( n15955 ) ;
assign n15957 =  ( n15950 ) | ( n15956 )  ;
assign n15958 = ~ ( n15957 ) ;
assign n15959 =  ( n15939 ) | ( n15958 )  ;
assign n15960 = ~ ( n15959 ) ;
assign n15961 =  ( n15932 ) | ( n15960 )  ;
assign n15962 = ~ ( n15961 ) ;
assign n15963 =  ( n15916 ) | ( n15962 )  ;
assign n15964 = ~ ( n15963 ) ;
assign n15965 =  ( n15904 ) | ( n15964 )  ;
assign n15966 = ~ ( n12343 ) ;
assign n15967 =  ( n15966 ) | ( n12426 )  ;
assign n15968 = ~ ( n12722 ) ;
assign n15969 =  ( n15967 ) | ( n15968 )  ;
assign n15970 =  ( n15969 ) | ( n12800 )  ;
assign n15971 = ~ ( n13119 ) ;
assign n15972 =  ( n15970 ) | ( n15971 )  ;
assign n15973 =  ( n15972 ) | ( n13226 )  ;
assign n15974 = ~ ( n13544 ) ;
assign n15975 =  ( n15973 ) | ( n15974 )  ;
assign n15976 = ~ ( n13683 ) ;
assign n15977 =  ( n15975 ) | ( n15976 )  ;
assign n15978 = ~ ( n13846 ) ;
assign n15979 =  ( n15977 ) | ( n15978 )  ;
assign n15980 = ~ ( n14019 ) ;
assign n15981 =  ( n15979 ) | ( n15980 )  ;
assign n15982 = ~ ( n14169 ) ;
assign n15983 =  ( n15981 ) | ( n15982 )  ;
assign n15984 = ~ ( n14288 ) ;
assign n15985 =  ( n15983 ) | ( n15984 )  ;
assign n15986 = ~ ( n14420 ) ;
assign n15987 =  ( n15985 ) | ( n15986 )  ;
assign n15988 = ~ ( n14543 ) ;
assign n15989 =  ( n15987 ) | ( n15988 )  ;
assign n15990 = ~ ( n14667 ) ;
assign n15991 =  ( n15989 ) | ( n15990 )  ;
assign n15992 = ~ ( n14754 ) ;
assign n15993 =  ( n15991 ) | ( n15992 )  ;
assign n15994 = ~ ( n14829 ) ;
assign n15995 =  ( n14861 ) | ( n14872 )  ;
assign n15996 = ~ ( n14895 ) ;
assign n15997 =  ( n15995 ) | ( n15996 )  ;
assign n15998 = ~ ( n15997 ) ;
assign n15999 =  ( n15994 ) | ( n15998 )  ;
assign n16000 = ~ ( n14952 ) ;
assign n16001 =  ( n14861 ) | ( n16000 )  ;
assign n16002 = ~ ( n15514 ) ;
assign n16003 =  ( n16001 ) | ( n16002 )  ;
assign n16004 = ~ ( n16003 ) ;
assign n16005 =  ( n15999 ) | ( n16004 )  ;
assign n16006 = ~ ( n14952 ) ;
assign n16007 =  ( n14861 ) | ( n16006 )  ;
assign n16008 = ~ ( n15042 ) ;
assign n16009 =  ( n16007 ) | ( n16008 )  ;
assign n16010 =  ( n16009 ) | ( n15084 )  ;
assign n16011 = ~ ( n15115 ) ;
assign n16012 =  ( n16011 ) | ( n15141 )  ;
assign n16013 = ~ ( n16012 ) ;
assign n16014 =  ( n16013 ) | ( n15198 )  ;
assign n16015 =  ( n16014 ) | ( n15545 )  ;
assign n16016 = ~ ( n16015 ) ;
assign n16017 =  ( n16010 ) | ( n16016 )  ;
assign n16018 = ~ ( n16017 ) ;
assign n16019 =  ( n16005 ) | ( n16018 )  ;
assign n16020 = ~ ( n14952 ) ;
assign n16021 =  ( n14861 ) | ( n16020 )  ;
assign n16022 = ~ ( n15042 ) ;
assign n16023 =  ( n16021 ) | ( n16022 )  ;
assign n16024 =  ( n16023 ) | ( n15084 )  ;
assign n16025 = ~ ( n15162 ) ;
assign n16026 =  ( n16024 ) | ( n16025 )  ;
assign n16027 =  ( n16026 ) | ( n15217 )  ;
assign n16028 =  ( n16027 ) | ( n15250 )  ;
assign n16029 =  ( n5648 ) ^ ( n15255 )  ;
assign n16030 =  ( n16029 ) ^ ( n7455 )  ;
assign n16031 =  ( n16030 ) ^ ( n15263 )  ;
assign n16032 = ~ ( n16031 ) ;
assign n16033 =  ( n16028 ) | ( n16032 )  ;
assign n16034 = ki[1:1] ;
assign n16035 =  ( n5657 ) ^ ( n16034 )  ;
assign n16036 = ~ ( n16035 ) ;
assign n16037 =  ( n16033 ) | ( n16036 )  ;
assign n16038 = kd[1:1] ;
assign n16039 =  ( n10564 ) ^ ( n16038 )  ;
assign n16040 = ~ ( n16039 ) ;
assign n16041 =  ( n16037 ) | ( n16040 )  ;
assign n16042 = ~ ( n16041 ) ;
assign n16043 =  ( n16019 ) | ( n16042 )  ;
assign n16044 = ~ ( n16043 ) ;
assign n16045 =  ( n15993 ) | ( n16044 )  ;
assign n16046 = ~ ( n16045 ) ;
assign n16047 =  ( n15965 ) | ( n16046 )  ;
assign n16048 = ~ ( n16047 ) ;
assign n16049 =  ( n12090 ) | ( n16048 )  ;
assign n16050 = ~ ( n16049 ) ;
assign n16051 =  ( n15865 ) | ( n16050 )  ;
assign n16052 =  ( n15863 ) ^ ( n16051 )  ;
assign n16053 =  { ( n15830 ) , ( n16052 ) }  ;
assign n16054 =  ( n1183 ) ^ ( n1199 )  ;
assign n16055 =  ( n16054 ) ^ ( n666 )  ;
assign n16056 =  ( n16055 ) ^ ( n682 )  ;
assign n16057 =  ( n16056 ) ^ ( n697 )  ;
assign n16058 =  ( n16057 ) ^ ( n759 )  ;
assign n16059 =  ( n16058 ) ^ ( n11806 )  ;
assign n16060 =  ( n16059 ) ^ ( n6216 )  ;
assign n16061 =  ( n16060 ) ^ ( n6242 )  ;
assign n16062 = ~ ( n5855 ) ;
assign n16063 = ~ ( n5867 ) ;
assign n16064 =  ( n16062 ) | ( n16063 )  ;
assign n16065 =  ( n16061 ) ^ ( n16064 )  ;
assign n16066 =  ( n5832 ) | ( n5841 )  ;
assign n16067 =  ( n16066 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16068 =  ( n16065 ) ^ ( n16067 )  ;
assign n16069 =  ( n5682 ) | ( n5691 )  ;
assign n16070 =  ( n16069 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16071 =  ( n16068 ) ^ ( n16070 )  ;
assign n16072 =  ( n5713 ) | ( n5722 )  ;
assign n16073 =  ( n16072 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16074 =  ( n16071 ) ^ ( n16073 )  ;
assign n16075 =  ( n16074 ) ^ ( n11996 )  ;
assign n16076 =  ( n16075 ) ^ ( n16047 )  ;
assign n16077 =  { ( n16053 ) , ( n16076 ) }  ;
assign n16078 =  ( n1436 ) ^ ( n1125 )  ;
assign n16079 =  ( n16078 ) ^ ( n1145 )  ;
assign n16080 =  ( n16079 ) ^ ( n1154 )  ;
assign n16081 =  ( n532 ) | ( n541 )  ;
assign n16082 =  ( n16081 ) ? ( bv_1_0_n2 ) : ( n557 ) ;
assign n16083 = ~ ( n16082 ) ;
assign n16084 =  ( n16080 ) ^ ( n16083 )  ;
assign n16085 =  ( n16084 ) ^ ( n624 )  ;
assign n16086 =  ( n16085 ) ^ ( n662 )  ;
assign n16087 =  ( n16086 ) ^ ( n1179 )  ;
assign n16088 =  ( n16087 ) ^ ( n12183 )  ;
assign n16089 = ~ ( n6402 ) ;
assign n16090 =  ( n16089 ) | ( n6421 )  ;
assign n16091 = ~ ( n16090 ) ;
assign n16092 =  ( n16088 ) ^ ( n16091 )  ;
assign n16093 = ~ ( n6105 ) ;
assign n16094 =  ( n6111 ) | ( n6124 )  ;
assign n16095 = ~ ( n16094 ) ;
assign n16096 =  ( n16093 ) | ( n16095 )  ;
assign n16097 =  ( n16092 ) ^ ( n16096 )  ;
assign n16098 =  ( n16097 ) ^ ( n6166 )  ;
assign n16099 = ~ ( n6173 ) ;
assign n16100 = ~ ( n5736 ) ;
assign n16101 =  ( n16099 ) | ( n16100 )  ;
assign n16102 =  ( n16098 ) ^ ( n16101 )  ;
assign n16103 =  ( n5802 ) | ( n5811 )  ;
assign n16104 =  ( n16103 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16105 = ~ ( n16104 ) ;
assign n16106 =  ( n16102 ) ^ ( n16105 )  ;
assign n16107 =  ( n5832 ) | ( n5841 )  ;
assign n16108 =  ( n16107 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16109 =  ( n16106 ) ^ ( n16108 )  ;
assign n16110 =  ( n5682 ) | ( n5691 )  ;
assign n16111 =  ( n16110 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16112 =  ( n16109 ) ^ ( n16111 )  ;
assign n16113 =  ( n5713 ) | ( n5722 )  ;
assign n16114 =  ( n16113 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16115 =  ( n16112 ) ^ ( n16114 )  ;
assign n16116 =  ( n16115 ) ^ ( n12300 )  ;
assign n16117 =  ( n12354 ) | ( n12376 )  ;
assign n16118 = ~ ( n16117 ) ;
assign n16119 = ~ ( n12535 ) ;
assign n16120 = ~ ( n12665 ) ;
assign n16121 =  ( n16119 ) | ( n16120 )  ;
assign n16122 = ~ ( n16121 ) ;
assign n16123 = ~ ( n12722 ) ;
assign n16124 =  ( n16123 ) | ( n12735 )  ;
assign n16125 =  ( n16124 ) | ( n12761 )  ;
assign n16126 = ~ ( n16125 ) ;
assign n16127 =  ( n16122 ) | ( n16126 )  ;
assign n16128 = ~ ( n12722 ) ;
assign n16129 =  ( n16128 ) | ( n12800 )  ;
assign n16130 = ~ ( n13172 ) ;
assign n16131 =  ( n16129 ) | ( n16130 )  ;
assign n16132 = ~ ( n16131 ) ;
assign n16133 =  ( n16127 ) | ( n16132 )  ;
assign n16134 =  ( n16133 ) | ( n13925 )  ;
assign n16135 = ~ ( n12722 ) ;
assign n16136 =  ( n16135 ) | ( n12800 )  ;
assign n16137 = ~ ( n13119 ) ;
assign n16138 =  ( n16136 ) | ( n16137 )  ;
assign n16139 =  ( n16138 ) | ( n13226 )  ;
assign n16140 = ~ ( n13544 ) ;
assign n16141 =  ( n16139 ) | ( n16140 )  ;
assign n16142 = ~ ( n13683 ) ;
assign n16143 =  ( n16141 ) | ( n16142 )  ;
assign n16144 = ~ ( n13846 ) ;
assign n16145 =  ( n16143 ) | ( n16144 )  ;
assign n16146 = ~ ( n14019 ) ;
assign n16147 =  ( n16145 ) | ( n16146 )  ;
assign n16148 = ~ ( n14106 ) ;
assign n16149 = ~ ( n14169 ) ;
assign n16150 =  ( n16149 ) | ( n14186 )  ;
assign n16151 = ~ ( n14227 ) ;
assign n16152 =  ( n16150 ) | ( n16151 )  ;
assign n16153 = ~ ( n16152 ) ;
assign n16154 =  ( n16148 ) | ( n16153 )  ;
assign n16155 = ~ ( n14169 ) ;
assign n16156 = ~ ( n14288 ) ;
assign n16157 =  ( n16155 ) | ( n16156 )  ;
assign n16158 = ~ ( n14480 ) ;
assign n16159 =  ( n16157 ) | ( n16158 )  ;
assign n16160 = ~ ( n16159 ) ;
assign n16161 =  ( n16154 ) | ( n16160 )  ;
assign n16162 =  ( n16161 ) | ( n14906 )  ;
assign n16163 = ~ ( n16162 ) ;
assign n16164 =  ( n16147 ) | ( n16163 )  ;
assign n16165 = ~ ( n16164 ) ;
assign n16166 =  ( n16134 ) | ( n16165 )  ;
assign n16167 = ~ ( n12722 ) ;
assign n16168 =  ( n16167 ) | ( n12800 )  ;
assign n16169 = ~ ( n13119 ) ;
assign n16170 =  ( n16168 ) | ( n16169 )  ;
assign n16171 =  ( n16170 ) | ( n13226 )  ;
assign n16172 = ~ ( n13544 ) ;
assign n16173 =  ( n16171 ) | ( n16172 )  ;
assign n16174 = ~ ( n13683 ) ;
assign n16175 =  ( n16173 ) | ( n16174 )  ;
assign n16176 = ~ ( n13846 ) ;
assign n16177 =  ( n16175 ) | ( n16176 )  ;
assign n16178 = ~ ( n14019 ) ;
assign n16179 =  ( n16177 ) | ( n16178 )  ;
assign n16180 = ~ ( n14169 ) ;
assign n16181 =  ( n16179 ) | ( n16180 )  ;
assign n16182 = ~ ( n14288 ) ;
assign n16183 =  ( n16181 ) | ( n16182 )  ;
assign n16184 = ~ ( n14420 ) ;
assign n16185 =  ( n16183 ) | ( n16184 )  ;
assign n16186 = ~ ( n14543 ) ;
assign n16187 =  ( n16185 ) | ( n16186 )  ;
assign n16188 = ~ ( n14667 ) ;
assign n16189 =  ( n16187 ) | ( n16188 )  ;
assign n16190 = ~ ( n14754 ) ;
assign n16191 =  ( n16189 ) | ( n16190 )  ;
assign n16192 =  ( n16191 ) | ( n14861 )  ;
assign n16193 = ~ ( n14952 ) ;
assign n16194 =  ( n16192 ) | ( n16193 )  ;
assign n16195 = ~ ( n15287 ) ;
assign n16196 =  ( n16194 ) | ( n16195 )  ;
assign n16197 = ~ ( n16196 ) ;
assign n16198 =  ( n16166 ) | ( n16197 )  ;
assign n16199 = ~ ( n16198 ) ;
assign n16200 =  ( n12426 ) | ( n16199 )  ;
assign n16201 = ~ ( n16200 ) ;
assign n16202 =  ( n16118 ) | ( n16201 )  ;
assign n16203 =  ( n16116 ) ^ ( n16202 )  ;
assign n16204 =  { ( n16077 ) , ( n16203 ) }  ;
assign n16205 =  ( n1773 ) ^ ( n1405 )  ;
assign n16206 =  ( n16205 ) ^ ( n1068 )  ;
assign n16207 =  ( n16206 ) ^ ( n1079 )  ;
assign n16208 =  ( n16207 ) ^ ( n1090 )  ;
assign n16209 =  ( n16208 ) ^ ( n1097 )  ;
assign n16210 =  ( n16209 ) ^ ( n1104 )  ;
assign n16211 =  ( n16210 ) ^ ( n1120 )  ;
assign n16212 =  ( n16211 ) ^ ( n12179 )  ;
assign n16213 =  ( n16212 ) ^ ( n6753 )  ;
assign n16214 =  ( n16213 ) ^ ( n6402 )  ;
assign n16215 =  ( n16214 ) ^ ( n6093 )  ;
assign n16216 = ~ ( n6100 ) ;
assign n16217 = ~ ( n5902 ) ;
assign n16218 =  ( n16216 ) | ( n16217 )  ;
assign n16219 =  ( n16215 ) ^ ( n16218 )  ;
assign n16220 =  ( n5802 ) | ( n5811 )  ;
assign n16221 =  ( n16220 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16222 =  ( n16219 ) ^ ( n16221 )  ;
assign n16223 =  ( n5832 ) | ( n5841 )  ;
assign n16224 =  ( n16223 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16225 =  ( n16222 ) ^ ( n16224 )  ;
assign n16226 =  ( n5682 ) | ( n5691 )  ;
assign n16227 =  ( n16226 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16228 =  ( n16225 ) ^ ( n16227 )  ;
assign n16229 =  ( n5713 ) | ( n5722 )  ;
assign n16230 =  ( n16229 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16231 =  ( n16228 ) ^ ( n16230 )  ;
assign n16232 =  ( n16231 ) ^ ( n12296 )  ;
assign n16233 =  ( n16232 ) ^ ( n16198 )  ;
assign n16234 =  { ( n16204 ) , ( n16233 ) }  ;
assign n16235 = ~ ( n2070 ) ;
assign n16236 =  ( n16235 ) | ( n2080 )  ;
assign n16237 = ~ ( n16236 ) ;
assign n16238 =  ( n16237 ) ^ ( n1740 )  ;
assign n16239 =  ( n16238 ) ^ ( n1755 )  ;
assign n16240 =  ( n16239 ) ^ ( n1379 )  ;
assign n16241 =  ( n16240 ) ^ ( n1389 )  ;
assign n16242 =  ( n873 ) | ( n882 )  ;
assign n16243 =  ( n16242 ) ? ( bv_1_0_n2 ) : ( n898 ) ;
assign n16244 = ~ ( n16243 ) ;
assign n16245 =  ( n16241 ) ^ ( n16244 )  ;
assign n16246 =  ( n16245 ) ^ ( n941 )  ;
assign n16247 =  ( n16246 ) ^ ( n967 )  ;
assign n16248 =  ( n16247 ) ^ ( n999 )  ;
assign n16249 =  ( n16248 ) ^ ( n1064 )  ;
assign n16250 =  ( n16249 ) ^ ( n12534 )  ;
assign n16251 = ~ ( n7022 ) ;
assign n16252 =  ( n16251 ) | ( n7045 )  ;
assign n16253 = ~ ( n16252 ) ;
assign n16254 =  ( n16250 ) ^ ( n16253 )  ;
assign n16255 =  ( n16254 ) ^ ( n6683 )  ;
assign n16256 = ~ ( n6690 ) ;
assign n16257 =  ( n6696 ) | ( n6711 )  ;
assign n16258 = ~ ( n16257 ) ;
assign n16259 =  ( n16256 ) | ( n16258 )  ;
assign n16260 =  ( n16255 ) ^ ( n16259 )  ;
assign n16261 = ~ ( n6330 ) ;
assign n16262 =  ( n6337 ) | ( n5909 )  ;
assign n16263 = ~ ( n16262 ) ;
assign n16264 =  ( n16261 ) | ( n16263 )  ;
assign n16265 = ~ ( n6356 ) ;
assign n16266 =  ( n16264 ) | ( n16265 )  ;
assign n16267 =  ( n16260 ) ^ ( n16266 )  ;
assign n16268 = ~ ( n6366 ) ;
assign n16269 = ~ ( n5902 ) ;
assign n16270 =  ( n16268 ) | ( n16269 )  ;
assign n16271 =  ( n16267 ) ^ ( n16270 )  ;
assign n16272 =  ( n6030 ) | ( n6039 )  ;
assign n16273 =  ( n16272 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16274 = ~ ( n16273 ) ;
assign n16275 =  ( n16271 ) ^ ( n16274 )  ;
assign n16276 =  ( n5802 ) | ( n5811 )  ;
assign n16277 =  ( n16276 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16278 =  ( n16275 ) ^ ( n16277 )  ;
assign n16279 =  ( n5832 ) | ( n5841 )  ;
assign n16280 =  ( n16279 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16281 =  ( n16278 ) ^ ( n16280 )  ;
assign n16282 =  ( n5682 ) | ( n5691 )  ;
assign n16283 =  ( n16282 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16284 =  ( n16281 ) ^ ( n16283 )  ;
assign n16285 =  ( n5713 ) | ( n5722 )  ;
assign n16286 =  ( n16285 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16287 =  ( n16284 ) ^ ( n16286 )  ;
assign n16288 =  ( n16287 ) ^ ( n12664 )  ;
assign n16289 =  ( n12735 ) | ( n12761 )  ;
assign n16290 = ~ ( n16289 ) ;
assign n16291 = ~ ( n12912 ) ;
assign n16292 = ~ ( n13055 ) ;
assign n16293 =  ( n16291 ) | ( n16292 )  ;
assign n16294 = ~ ( n16293 ) ;
assign n16295 = ~ ( n13119 ) ;
assign n16296 =  ( n16295 ) | ( n13136 )  ;
assign n16297 =  ( n16296 ) | ( n13169 )  ;
assign n16298 = ~ ( n16297 ) ;
assign n16299 =  ( n16294 ) | ( n16298 )  ;
assign n16300 = ~ ( n13119 ) ;
assign n16301 =  ( n16300 ) | ( n13226 )  ;
assign n16302 = ~ ( n15401 ) ;
assign n16303 =  ( n16301 ) | ( n16302 )  ;
assign n16304 = ~ ( n16303 ) ;
assign n16305 =  ( n16299 ) | ( n16304 )  ;
assign n16306 =  ( n16305 ) | ( n15437 )  ;
assign n16307 = ~ ( n13119 ) ;
assign n16308 =  ( n16307 ) | ( n13226 )  ;
assign n16309 = ~ ( n13544 ) ;
assign n16310 =  ( n16308 ) | ( n16309 )  ;
assign n16311 = ~ ( n13683 ) ;
assign n16312 =  ( n16310 ) | ( n16311 )  ;
assign n16313 = ~ ( n13846 ) ;
assign n16314 =  ( n16312 ) | ( n16313 )  ;
assign n16315 = ~ ( n14019 ) ;
assign n16316 =  ( n16314 ) | ( n16315 )  ;
assign n16317 = ~ ( n14169 ) ;
assign n16318 =  ( n16316 ) | ( n16317 )  ;
assign n16319 = ~ ( n14288 ) ;
assign n16320 =  ( n16318 ) | ( n16319 )  ;
assign n16321 = ~ ( n14321 ) ;
assign n16322 = ~ ( n14365 ) ;
assign n16323 =  ( n16321 ) | ( n16322 )  ;
assign n16324 = ~ ( n16323 ) ;
assign n16325 = ~ ( n14420 ) ;
assign n16326 = ~ ( n14441 ) ;
assign n16327 =  ( n16325 ) | ( n16326 )  ;
assign n16328 = ~ ( n14476 ) ;
assign n16329 =  ( n16327 ) | ( n16328 )  ;
assign n16330 = ~ ( n16329 ) ;
assign n16331 =  ( n16324 ) | ( n16330 )  ;
assign n16332 = ~ ( n14420 ) ;
assign n16333 = ~ ( n14543 ) ;
assign n16334 =  ( n16332 ) | ( n16333 )  ;
assign n16335 = ~ ( n15489 ) ;
assign n16336 =  ( n16334 ) | ( n16335 )  ;
assign n16337 = ~ ( n16336 ) ;
assign n16338 =  ( n16331 ) | ( n16337 )  ;
assign n16339 =  ( n16338 ) | ( n15521 )  ;
assign n16340 = ~ ( n16339 ) ;
assign n16341 =  ( n16320 ) | ( n16340 )  ;
assign n16342 = ~ ( n16341 ) ;
assign n16343 =  ( n16306 ) | ( n16342 )  ;
assign n16344 = ~ ( n13119 ) ;
assign n16345 =  ( n16344 ) | ( n13226 )  ;
assign n16346 = ~ ( n13544 ) ;
assign n16347 =  ( n16345 ) | ( n16346 )  ;
assign n16348 = ~ ( n13683 ) ;
assign n16349 =  ( n16347 ) | ( n16348 )  ;
assign n16350 = ~ ( n13846 ) ;
assign n16351 =  ( n16349 ) | ( n16350 )  ;
assign n16352 = ~ ( n14019 ) ;
assign n16353 =  ( n16351 ) | ( n16352 )  ;
assign n16354 = ~ ( n14169 ) ;
assign n16355 =  ( n16353 ) | ( n16354 )  ;
assign n16356 = ~ ( n14288 ) ;
assign n16357 =  ( n16355 ) | ( n16356 )  ;
assign n16358 = ~ ( n14420 ) ;
assign n16359 =  ( n16357 ) | ( n16358 )  ;
assign n16360 = ~ ( n14543 ) ;
assign n16361 =  ( n16359 ) | ( n16360 )  ;
assign n16362 = ~ ( n14667 ) ;
assign n16363 =  ( n16361 ) | ( n16362 )  ;
assign n16364 = ~ ( n14754 ) ;
assign n16365 =  ( n16363 ) | ( n16364 )  ;
assign n16366 =  ( n16365 ) | ( n14861 )  ;
assign n16367 = ~ ( n14952 ) ;
assign n16368 =  ( n16366 ) | ( n16367 )  ;
assign n16369 = ~ ( n15042 ) ;
assign n16370 =  ( n16368 ) | ( n16369 )  ;
assign n16371 =  ( n16370 ) | ( n15084 )  ;
assign n16372 = ~ ( n15564 ) ;
assign n16373 =  ( n16371 ) | ( n16372 )  ;
assign n16374 = ~ ( n16373 ) ;
assign n16375 =  ( n16343 ) | ( n16374 )  ;
assign n16376 = ~ ( n16375 ) ;
assign n16377 =  ( n12800 ) | ( n16376 )  ;
assign n16378 = ~ ( n16377 ) ;
assign n16379 =  ( n16290 ) | ( n16378 )  ;
assign n16380 =  ( n16288 ) ^ ( n16379 )  ;
assign n16381 =  { ( n16234 ) , ( n16380 ) }  ;
assign n16382 =  ( n2426 ) ^ ( n2070 )  ;
assign n16383 =  ( n16382 ) ^ ( n1682 )  ;
assign n16384 =  ( n16383 ) ^ ( n1713 )  ;
assign n16385 =  ( n16384 ) ^ ( n1723 )  ;
assign n16386 =  ( n16385 ) ^ ( n1281 )  ;
assign n16387 =  ( n16386 ) ^ ( n1297 )  ;
assign n16388 =  ( n16387 ) ^ ( n1314 )  ;
assign n16389 =  ( n16388 ) ^ ( n1331 )  ;
assign n16390 =  ( n16389 ) ^ ( n1375 )  ;
assign n16391 =  ( n16390 ) ^ ( n12530 )  ;
assign n16392 =  ( n16391 ) ^ ( n7392 )  ;
assign n16393 =  ( n16392 ) ^ ( n7022 )  ;
assign n16394 =  ( n16393 ) ^ ( n6589 )  ;
assign n16395 =  ( n16394 ) ^ ( n6634 )  ;
assign n16396 = ~ ( n6640 ) ;
assign n16397 = ~ ( n6173 ) ;
assign n16398 =  ( n16396 ) | ( n16397 )  ;
assign n16399 =  ( n16395 ) ^ ( n16398 )  ;
assign n16400 =  ( n6030 ) | ( n6039 )  ;
assign n16401 =  ( n16400 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16402 =  ( n16399 ) ^ ( n16401 )  ;
assign n16403 =  ( n5802 ) | ( n5811 )  ;
assign n16404 =  ( n16403 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16405 =  ( n16402 ) ^ ( n16404 )  ;
assign n16406 =  ( n5832 ) | ( n5841 )  ;
assign n16407 =  ( n16406 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16408 =  ( n16405 ) ^ ( n16407 )  ;
assign n16409 =  ( n5682 ) | ( n5691 )  ;
assign n16410 =  ( n16409 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16411 =  ( n16408 ) ^ ( n16410 )  ;
assign n16412 =  ( n5713 ) | ( n5722 )  ;
assign n16413 =  ( n16412 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16414 =  ( n16411 ) ^ ( n16413 )  ;
assign n16415 =  ( n16414 ) ^ ( n12660 )  ;
assign n16416 =  ( n16415 ) ^ ( n16375 )  ;
assign n16417 =  { ( n16381 ) , ( n16416 ) }  ;
assign n16418 = ~ ( n2727 ) ;
assign n16419 =  ( n16418 ) ^ ( n2388 )  ;
assign n16420 =  ( n16419 ) ^ ( n2038 )  ;
assign n16421 =  ( n16420 ) ^ ( n2052 )  ;
assign n16422 =  ( n16421 ) ^ ( n1632 )  ;
assign n16423 =  ( n16422 ) ^ ( n1642 )  ;
assign n16424 =  ( n1475 ) | ( n1484 )  ;
assign n16425 =  ( n16424 ) ? ( bv_1_0_n2 ) : ( n1511 ) ;
assign n16426 = ~ ( n16425 ) ;
assign n16427 =  ( n16423 ) ^ ( n16426 )  ;
assign n16428 =  ( n16427 ) ^ ( n1656 )  ;
assign n16429 =  ( n16428 ) ^ ( n1663 )  ;
assign n16430 =  ( n16429 ) ^ ( n1670 )  ;
assign n16431 =  ( n16430 ) ^ ( n1677 )  ;
assign n16432 =  ( n16431 ) ^ ( n2422 )  ;
assign n16433 =  ( n16432 ) ^ ( n12911 )  ;
assign n16434 = ~ ( n7649 ) ;
assign n16435 =  ( n16434 ) | ( n7679 )  ;
assign n16436 = ~ ( n16435 ) ;
assign n16437 =  ( n16433 ) ^ ( n16436 )  ;
assign n16438 = ~ ( n7281 ) ;
assign n16439 =  ( n7287 ) | ( n7311 )  ;
assign n16440 = ~ ( n16439 ) ;
assign n16441 =  ( n16438 ) | ( n16440 )  ;
assign n16442 =  ( n16437 ) ^ ( n16441 )  ;
assign n16443 =  ( n16442 ) ^ ( n6970 )  ;
assign n16444 = ~ ( n6977 ) ;
assign n16445 = ~ ( n6982 ) ;
assign n16446 =  ( n16444 ) | ( n16445 )  ;
assign n16447 =  ( n16443 ) ^ ( n16446 )  ;
assign n16448 = ~ ( n6517 ) ;
assign n16449 =  ( n6524 ) | ( n6150 )  ;
assign n16450 = ~ ( n16449 ) ;
assign n16451 =  ( n16448 ) | ( n16450 )  ;
assign n16452 = ~ ( n6543 ) ;
assign n16453 =  ( n16451 ) | ( n16452 )  ;
assign n16454 =  ( n16447 ) ^ ( n16453 )  ;
assign n16455 = ~ ( n6553 ) ;
assign n16456 = ~ ( n6173 ) ;
assign n16457 =  ( n16455 ) | ( n16456 )  ;
assign n16458 =  ( n16454 ) ^ ( n16457 )  ;
assign n16459 =  ( n6483 ) | ( n6492 )  ;
assign n16460 =  ( n16459 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n16461 = ~ ( n16460 ) ;
assign n16462 =  ( n16458 ) ^ ( n16461 )  ;
assign n16463 =  ( n6030 ) | ( n6039 )  ;
assign n16464 =  ( n16463 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16465 =  ( n16462 ) ^ ( n16464 )  ;
assign n16466 =  ( n5802 ) | ( n5811 )  ;
assign n16467 =  ( n16466 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16468 =  ( n16465 ) ^ ( n16467 )  ;
assign n16469 =  ( n5832 ) | ( n5841 )  ;
assign n16470 =  ( n16469 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16471 =  ( n16468 ) ^ ( n16470 )  ;
assign n16472 =  ( n5682 ) | ( n5691 )  ;
assign n16473 =  ( n16472 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16474 =  ( n16471 ) ^ ( n16473 )  ;
assign n16475 =  ( n5713 ) | ( n5722 )  ;
assign n16476 =  ( n16475 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16477 =  ( n16474 ) ^ ( n16476 )  ;
assign n16478 =  ( n16477 ) ^ ( n13054 )  ;
assign n16479 =  ( n13136 ) | ( n13169 )  ;
assign n16480 = ~ ( n16479 ) ;
assign n16481 = ~ ( n13334 ) ;
assign n16482 = ~ ( n13471 ) ;
assign n16483 =  ( n16481 ) | ( n16482 )  ;
assign n16484 = ~ ( n16483 ) ;
assign n16485 = ~ ( n13544 ) ;
assign n16486 =  ( n16485 ) | ( n13568 )  ;
assign n16487 = ~ ( n13613 ) ;
assign n16488 =  ( n16486 ) | ( n16487 )  ;
assign n16489 = ~ ( n16488 ) ;
assign n16490 =  ( n16484 ) | ( n16489 )  ;
assign n16491 = ~ ( n13544 ) ;
assign n16492 = ~ ( n13683 ) ;
assign n16493 =  ( n16491 ) | ( n16492 )  ;
assign n16494 = ~ ( n13918 ) ;
assign n16495 =  ( n16493 ) | ( n16494 )  ;
assign n16496 = ~ ( n16495 ) ;
assign n16497 =  ( n16490 ) | ( n16496 )  ;
assign n16498 =  ( n16497 ) | ( n15715 )  ;
assign n16499 = ~ ( n13544 ) ;
assign n16500 = ~ ( n13683 ) ;
assign n16501 =  ( n16499 ) | ( n16500 )  ;
assign n16502 = ~ ( n13846 ) ;
assign n16503 =  ( n16501 ) | ( n16502 )  ;
assign n16504 = ~ ( n14019 ) ;
assign n16505 =  ( n16503 ) | ( n16504 )  ;
assign n16506 = ~ ( n14169 ) ;
assign n16507 =  ( n16505 ) | ( n16506 )  ;
assign n16508 = ~ ( n14288 ) ;
assign n16509 =  ( n16507 ) | ( n16508 )  ;
assign n16510 = ~ ( n14420 ) ;
assign n16511 =  ( n16509 ) | ( n16510 )  ;
assign n16512 = ~ ( n14543 ) ;
assign n16513 =  ( n16511 ) | ( n16512 )  ;
assign n16514 = ~ ( n14620 ) ;
assign n16515 = ~ ( n14667 ) ;
assign n16516 =  ( n16515 ) | ( n14683 )  ;
assign n16517 = ~ ( n14709 ) ;
assign n16518 =  ( n16516 ) | ( n16517 )  ;
assign n16519 = ~ ( n16518 ) ;
assign n16520 =  ( n16514 ) | ( n16519 )  ;
assign n16521 = ~ ( n14667 ) ;
assign n16522 = ~ ( n14754 ) ;
assign n16523 =  ( n16521 ) | ( n16522 )  ;
assign n16524 = ~ ( n14899 ) ;
assign n16525 =  ( n16523 ) | ( n16524 )  ;
assign n16526 = ~ ( n16525 ) ;
assign n16527 =  ( n16520 ) | ( n16526 )  ;
assign n16528 =  ( n16527 ) | ( n15782 )  ;
assign n16529 = ~ ( n16528 ) ;
assign n16530 =  ( n16513 ) | ( n16529 )  ;
assign n16531 = ~ ( n16530 ) ;
assign n16532 =  ( n16498 ) | ( n16531 )  ;
assign n16533 = ~ ( n13544 ) ;
assign n16534 = ~ ( n13683 ) ;
assign n16535 =  ( n16533 ) | ( n16534 )  ;
assign n16536 = ~ ( n13846 ) ;
assign n16537 =  ( n16535 ) | ( n16536 )  ;
assign n16538 = ~ ( n14019 ) ;
assign n16539 =  ( n16537 ) | ( n16538 )  ;
assign n16540 = ~ ( n14169 ) ;
assign n16541 =  ( n16539 ) | ( n16540 )  ;
assign n16542 = ~ ( n14288 ) ;
assign n16543 =  ( n16541 ) | ( n16542 )  ;
assign n16544 = ~ ( n14420 ) ;
assign n16545 =  ( n16543 ) | ( n16544 )  ;
assign n16546 = ~ ( n14543 ) ;
assign n16547 =  ( n16545 ) | ( n16546 )  ;
assign n16548 = ~ ( n14667 ) ;
assign n16549 =  ( n16547 ) | ( n16548 )  ;
assign n16550 = ~ ( n14754 ) ;
assign n16551 =  ( n16549 ) | ( n16550 )  ;
assign n16552 =  ( n16551 ) | ( n14861 )  ;
assign n16553 = ~ ( n14952 ) ;
assign n16554 =  ( n16552 ) | ( n16553 )  ;
assign n16555 = ~ ( n15042 ) ;
assign n16556 =  ( n16554 ) | ( n16555 )  ;
assign n16557 =  ( n16556 ) | ( n15084 )  ;
assign n16558 = ~ ( n15162 ) ;
assign n16559 =  ( n16557 ) | ( n16558 )  ;
assign n16560 =  ( n16559 ) | ( n15217 )  ;
assign n16561 =  ( n15242 ) | ( n15267 )  ;
assign n16562 = ~ ( n15281 ) ;
assign n16563 =  ( n16561 ) | ( n16562 )  ;
assign n16564 = ~ ( n16563 ) ;
assign n16565 =  ( n16560 ) | ( n16564 )  ;
assign n16566 = ~ ( n16565 ) ;
assign n16567 =  ( n16532 ) | ( n16566 )  ;
assign n16568 = ~ ( n16567 ) ;
assign n16569 =  ( n13226 ) | ( n16568 )  ;
assign n16570 = ~ ( n16569 ) ;
assign n16571 =  ( n16480 ) | ( n16570 )  ;
assign n16572 =  ( n16478 ) ^ ( n16571 )  ;
assign n16573 =  { ( n16417 ) , ( n16572 ) }  ;
assign n16574 = ~ ( n2692 ) ;
assign n16575 =  ( n2675 ) | ( n16574 )  ;
assign n16576 =  ( n3043 ) ^ ( n16575 )  ;
assign n16577 =  ( n16576 ) ^ ( n2361 )  ;
assign n16578 =  ( n16577 ) ^ ( n2371 )  ;
assign n16579 =  ( n16578 ) ^ ( n1952 )  ;
assign n16580 =  ( n16579 ) ^ ( n1963 )  ;
assign n16581 =  ( n16580 ) ^ ( n1513 )  ;
assign n16582 =  ( n16581 ) ^ ( n1538 )  ;
assign n16583 =  ( n16582 ) ^ ( n1564 )  ;
assign n16584 =  ( n16583 ) ^ ( n1590 )  ;
assign n16585 =  ( n16584 ) ^ ( n1628 )  ;
assign n16586 =  ( n16585 ) ^ ( n2016 )  ;
assign n16587 =  ( n16586 ) ^ ( n12907 )  ;
assign n16588 =  ( n16587 ) ^ ( n8047 )  ;
assign n16589 =  ( n16588 ) ^ ( n7649 )  ;
assign n16590 =  ( n16589 ) ^ ( n7265 )  ;
assign n16591 = ~ ( n7271 ) ;
assign n16592 = ~ ( n7277 ) ;
assign n16593 =  ( n16591 ) | ( n16592 )  ;
assign n16594 =  ( n16590 ) ^ ( n16593 )  ;
assign n16595 =  ( n16594 ) ^ ( n6888 )  ;
assign n16596 = ~ ( n6895 ) ;
assign n16597 = ~ ( n6366 ) ;
assign n16598 =  ( n16596 ) | ( n16597 )  ;
assign n16599 =  ( n16595 ) ^ ( n16598 )  ;
assign n16600 =  ( n6483 ) | ( n6492 )  ;
assign n16601 =  ( n16600 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n16602 =  ( n16599 ) ^ ( n16601 )  ;
assign n16603 =  ( n6030 ) | ( n6039 )  ;
assign n16604 =  ( n16603 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16605 =  ( n16602 ) ^ ( n16604 )  ;
assign n16606 =  ( n5802 ) | ( n5811 )  ;
assign n16607 =  ( n16606 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16608 =  ( n16605 ) ^ ( n16607 )  ;
assign n16609 =  ( n5832 ) | ( n5841 )  ;
assign n16610 =  ( n16609 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16611 =  ( n16608 ) ^ ( n16610 )  ;
assign n16612 =  ( n5682 ) | ( n5691 )  ;
assign n16613 =  ( n16612 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16614 =  ( n16611 ) ^ ( n16613 )  ;
assign n16615 =  ( n5713 ) | ( n5722 )  ;
assign n16616 =  ( n16615 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16617 =  ( n16614 ) ^ ( n16616 )  ;
assign n16618 =  ( n16617 ) ^ ( n13050 )  ;
assign n16619 =  ( n16618 ) ^ ( n16567 )  ;
assign n16620 =  { ( n16573 ) , ( n16619 ) }  ;
assign n16621 = ~ ( n3371 ) ;
assign n16622 = ~ ( n2973 ) ;
assign n16623 =  ( n16622 ) | ( n2994 )  ;
assign n16624 =  ( n16621 ) ^ ( n16623 )  ;
assign n16625 =  ( n2633 ) | ( n2643 )  ;
assign n16626 =  ( n16625 ) | ( n2657 )  ;
assign n16627 =  ( n16624 ) ^ ( n16626 )  ;
assign n16628 =  ( n16627 ) ^ ( n2672 )  ;
assign n16629 =  ( n16628 ) ^ ( n2227 )  ;
assign n16630 =  ( n16629 ) ^ ( n2237 )  ;
assign n16631 =  ( n16630 ) ^ ( n2314 )  ;
assign n16632 =  ( n1838 ) | ( n1847 )  ;
assign n16633 =  ( n16632 ) ? ( bv_1_0_n2 ) : ( n1863 ) ;
assign n16634 = ~ ( n16633 ) ;
assign n16635 =  ( n16631 ) ^ ( n16634 )  ;
assign n16636 =  ( n16635 ) ^ ( n1879 )  ;
assign n16637 =  ( n16636 ) ^ ( n1896 )  ;
assign n16638 =  ( n16637 ) ^ ( n1913 )  ;
assign n16639 =  ( n16638 ) ^ ( n1948 )  ;
assign n16640 =  ( n16639 ) ^ ( n2357 )  ;
assign n16641 =  ( n16640 ) ^ ( n3039 )  ;
assign n16642 =  ( n16641 ) ^ ( n13333 )  ;
assign n16643 = ~ ( n8279 ) ;
assign n16644 = ~ ( n8321 ) ;
assign n16645 =  ( n16643 ) | ( n16644 )  ;
assign n16646 = ~ ( n16645 ) ;
assign n16647 =  ( n16642 ) ^ ( n16646 )  ;
assign n16648 =  ( n16647 ) ^ ( n7961 )  ;
assign n16649 =  ( n16648 ) ^ ( n7591 )  ;
assign n16650 = ~ ( n7597 ) ;
assign n16651 = ~ ( n7603 ) ;
assign n16652 =  ( n16650 ) | ( n16651 )  ;
assign n16653 =  ( n16649 ) ^ ( n16652 )  ;
assign n16654 = ~ ( n7133 ) ;
assign n16655 =  ( n7140 ) | ( n6337 )  ;
assign n16656 = ~ ( n16655 ) ;
assign n16657 =  ( n16654 ) | ( n16656 )  ;
assign n16658 = ~ ( n7159 ) ;
assign n16659 =  ( n16657 ) | ( n16658 )  ;
assign n16660 =  ( n16653 ) ^ ( n16659 )  ;
assign n16661 = ~ ( n7169 ) ;
assign n16662 = ~ ( n6366 ) ;
assign n16663 =  ( n16661 ) | ( n16662 )  ;
assign n16664 =  ( n16660 ) ^ ( n16663 )  ;
assign n16665 = ~ ( n5736 ) ;
assign n16666 =  ( n16665 ) | ( n5742 )  ;
assign n16667 =  ( n16664 ) ^ ( n16666 )  ;
assign n16668 =  ( n6825 ) | ( n6834 )  ;
assign n16669 =  ( n16668 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n16670 = ~ ( n16669 ) ;
assign n16671 =  ( n16667 ) ^ ( n16670 )  ;
assign n16672 =  ( n6483 ) | ( n6492 )  ;
assign n16673 =  ( n16672 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n16674 =  ( n16671 ) ^ ( n16673 )  ;
assign n16675 =  ( n6030 ) | ( n6039 )  ;
assign n16676 =  ( n16675 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16677 =  ( n16674 ) ^ ( n16676 )  ;
assign n16678 =  ( n5802 ) | ( n5811 )  ;
assign n16679 =  ( n16678 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16680 =  ( n16677 ) ^ ( n16679 )  ;
assign n16681 =  ( n5832 ) | ( n5841 )  ;
assign n16682 =  ( n16681 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16683 =  ( n16680 ) ^ ( n16682 )  ;
assign n16684 =  ( n5682 ) | ( n5691 )  ;
assign n16685 =  ( n16684 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16686 =  ( n16683 ) ^ ( n16685 )  ;
assign n16687 =  ( n5713 ) | ( n5722 )  ;
assign n16688 =  ( n16687 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16689 =  ( n16686 ) ^ ( n16688 )  ;
assign n16690 =  ( n16689 ) ^ ( n13470 )  ;
assign n16691 = ~ ( n13613 ) ;
assign n16692 =  ( n13568 ) | ( n16691 )  ;
assign n16693 = ~ ( n16692 ) ;
assign n16694 = ~ ( n13683 ) ;
assign n16695 = ~ ( n13775 ) ;
assign n16696 =  ( n13717 ) | ( n16695 )  ;
assign n16697 = ~ ( n16696 ) ;
assign n16698 = ~ ( n13846 ) ;
assign n16699 =  ( n16698 ) | ( n13867 )  ;
assign n16700 = ~ ( n13914 ) ;
assign n16701 =  ( n16699 ) | ( n16700 )  ;
assign n16702 = ~ ( n16701 ) ;
assign n16703 =  ( n16697 ) | ( n16702 )  ;
assign n16704 = ~ ( n13846 ) ;
assign n16705 = ~ ( n14019 ) ;
assign n16706 =  ( n16704 ) | ( n16705 )  ;
assign n16707 = ~ ( n15430 ) ;
assign n16708 =  ( n16706 ) | ( n16707 )  ;
assign n16709 = ~ ( n16708 ) ;
assign n16710 =  ( n16703 ) | ( n16709 )  ;
assign n16711 =  ( n16710 ) | ( n15960 )  ;
assign n16712 = ~ ( n13846 ) ;
assign n16713 = ~ ( n14019 ) ;
assign n16714 =  ( n16712 ) | ( n16713 )  ;
assign n16715 = ~ ( n14169 ) ;
assign n16716 =  ( n16714 ) | ( n16715 )  ;
assign n16717 = ~ ( n14288 ) ;
assign n16718 =  ( n16716 ) | ( n16717 )  ;
assign n16719 = ~ ( n14420 ) ;
assign n16720 =  ( n16718 ) | ( n16719 )  ;
assign n16721 = ~ ( n14543 ) ;
assign n16722 =  ( n16720 ) | ( n16721 )  ;
assign n16723 = ~ ( n14667 ) ;
assign n16724 =  ( n16722 ) | ( n16723 )  ;
assign n16725 = ~ ( n14754 ) ;
assign n16726 =  ( n16724 ) | ( n16725 )  ;
assign n16727 = ~ ( n14829 ) ;
assign n16728 =  ( n14861 ) | ( n14872 )  ;
assign n16729 = ~ ( n14895 ) ;
assign n16730 =  ( n16728 ) | ( n16729 )  ;
assign n16731 = ~ ( n16730 ) ;
assign n16732 =  ( n16727 ) | ( n16731 )  ;
assign n16733 = ~ ( n14952 ) ;
assign n16734 =  ( n14861 ) | ( n16733 )  ;
assign n16735 = ~ ( n15514 ) ;
assign n16736 =  ( n16734 ) | ( n16735 )  ;
assign n16737 = ~ ( n16736 ) ;
assign n16738 =  ( n16732 ) | ( n16737 )  ;
assign n16739 =  ( n16738 ) | ( n16018 )  ;
assign n16740 = ~ ( n16739 ) ;
assign n16741 =  ( n16726 ) | ( n16740 )  ;
assign n16742 = ~ ( n16741 ) ;
assign n16743 =  ( n16711 ) | ( n16742 )  ;
assign n16744 = ~ ( n13846 ) ;
assign n16745 = ~ ( n14019 ) ;
assign n16746 =  ( n16744 ) | ( n16745 )  ;
assign n16747 = ~ ( n14169 ) ;
assign n16748 =  ( n16746 ) | ( n16747 )  ;
assign n16749 = ~ ( n14288 ) ;
assign n16750 =  ( n16748 ) | ( n16749 )  ;
assign n16751 = ~ ( n14420 ) ;
assign n16752 =  ( n16750 ) | ( n16751 )  ;
assign n16753 = ~ ( n14543 ) ;
assign n16754 =  ( n16752 ) | ( n16753 )  ;
assign n16755 = ~ ( n14667 ) ;
assign n16756 =  ( n16754 ) | ( n16755 )  ;
assign n16757 = ~ ( n14754 ) ;
assign n16758 =  ( n16756 ) | ( n16757 )  ;
assign n16759 =  ( n16758 ) | ( n14861 )  ;
assign n16760 = ~ ( n14952 ) ;
assign n16761 =  ( n16759 ) | ( n16760 )  ;
assign n16762 = ~ ( n15042 ) ;
assign n16763 =  ( n16761 ) | ( n16762 )  ;
assign n16764 =  ( n16763 ) | ( n15084 )  ;
assign n16765 = ~ ( n15162 ) ;
assign n16766 =  ( n16764 ) | ( n16765 )  ;
assign n16767 =  ( n16766 ) | ( n15217 )  ;
assign n16768 =  ( n16767 ) | ( n15250 )  ;
assign n16769 =  ( n5648 ) ^ ( n15255 )  ;
assign n16770 =  ( n16769 ) ^ ( n7455 )  ;
assign n16771 =  ( n16770 ) ^ ( n15263 )  ;
assign n16772 = ~ ( n16771 ) ;
assign n16773 =  ( n16768 ) | ( n16772 )  ;
assign n16774 = ki[1:1] ;
assign n16775 =  ( n5657 ) ^ ( n16774 )  ;
assign n16776 = ~ ( n16775 ) ;
assign n16777 =  ( n16773 ) | ( n16776 )  ;
assign n16778 = kd[1:1] ;
assign n16779 =  ( n10564 ) ^ ( n16778 )  ;
assign n16780 = ~ ( n16779 ) ;
assign n16781 =  ( n16777 ) | ( n16780 )  ;
assign n16782 = ~ ( n16781 ) ;
assign n16783 =  ( n16743 ) | ( n16782 )  ;
assign n16784 = ~ ( n16783 ) ;
assign n16785 =  ( n16694 ) | ( n16784 )  ;
assign n16786 = ~ ( n16785 ) ;
assign n16787 =  ( n16693 ) | ( n16786 )  ;
assign n16788 =  ( n16690 ) ^ ( n16787 )  ;
assign n16789 =  { ( n16620 ) , ( n16788 ) }  ;
assign n16790 = ~ ( n3323 ) ;
assign n16791 =  ( n3306 ) | ( n16790 )  ;
assign n16792 =  ( n3623 ) ^ ( n16791 )  ;
assign n16793 = ~ ( n2928 ) ;
assign n16794 = ~ ( n2939 ) ;
assign n16795 =  ( n16793 ) | ( n16794 )  ;
assign n16796 = ~ ( n2954 ) ;
assign n16797 =  ( n16795 ) | ( n16796 )  ;
assign n16798 =  ( n16792 ) ^ ( n16797 )  ;
assign n16799 =  ( n16798 ) ^ ( n2971 )  ;
assign n16800 =  ( n16799 ) ^ ( n2552 )  ;
assign n16801 =  ( n16800 ) ^ ( n2561 )  ;
assign n16802 =  ( n16801 ) ^ ( n2624 )  ;
assign n16803 =  ( n16802 ) ^ ( n2144 )  ;
assign n16804 =  ( n16803 ) ^ ( n2160 )  ;
assign n16805 =  ( n16804 ) ^ ( n2177 )  ;
assign n16806 =  ( n16805 ) ^ ( n2194 )  ;
assign n16807 =  ( n16806 ) ^ ( n2223 )  ;
assign n16808 =  ( n16807 ) ^ ( n2263 )  ;
assign n16809 =  ( n16808 ) ^ ( n2309 )  ;
assign n16810 =  ( n16809 ) ^ ( n13329 )  ;
assign n16811 =  ( n16810 ) ^ ( n8625 )  ;
assign n16812 =  ( n16811 ) ^ ( n8279 )  ;
assign n16813 =  ( n16812 ) ^ ( n7899 )  ;
assign n16814 = ~ ( n7905 ) ;
assign n16815 = ~ ( n7911 ) ;
assign n16816 =  ( n16814 ) | ( n16815 )  ;
assign n16817 =  ( n16813 ) ^ ( n16816 )  ;
assign n16818 = ~ ( n7467 ) ;
assign n16819 =  ( n7473 ) | ( n6524 )  ;
assign n16820 = ~ ( n16819 ) ;
assign n16821 =  ( n16818 ) | ( n16820 )  ;
assign n16822 = ~ ( n7491 ) ;
assign n16823 =  ( n16821 ) | ( n16822 )  ;
assign n16824 =  ( n16817 ) ^ ( n16823 )  ;
assign n16825 = ~ ( n7498 ) ;
assign n16826 = ~ ( n6553 ) ;
assign n16827 =  ( n16825 ) | ( n16826 )  ;
assign n16828 =  ( n16824 ) ^ ( n16827 )  ;
assign n16829 = ~ ( n5902 ) ;
assign n16830 = ~ ( n5913 ) ;
assign n16831 =  ( n16829 ) | ( n16830 )  ;
assign n16832 =  ( n16828 ) ^ ( n16831 )  ;
assign n16833 =  ( n6825 ) | ( n6834 )  ;
assign n16834 =  ( n16833 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n16835 =  ( n16832 ) ^ ( n16834 )  ;
assign n16836 =  ( n6483 ) | ( n6492 )  ;
assign n16837 =  ( n16836 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n16838 =  ( n16835 ) ^ ( n16837 )  ;
assign n16839 =  ( n6030 ) | ( n6039 )  ;
assign n16840 =  ( n16839 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16841 =  ( n16838 ) ^ ( n16840 )  ;
assign n16842 =  ( n5802 ) | ( n5811 )  ;
assign n16843 =  ( n16842 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16844 =  ( n16841 ) ^ ( n16843 )  ;
assign n16845 =  ( n5832 ) | ( n5841 )  ;
assign n16846 =  ( n16845 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16847 =  ( n16844 ) ^ ( n16846 )  ;
assign n16848 =  ( n5682 ) | ( n5691 )  ;
assign n16849 =  ( n16848 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16850 =  ( n16847 ) ^ ( n16849 )  ;
assign n16851 =  ( n5713 ) | ( n5722 )  ;
assign n16852 =  ( n16851 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16853 =  ( n16850 ) ^ ( n16852 )  ;
assign n16854 =  ( n16853 ) ^ ( n13466 )  ;
assign n16855 =  ( n16854 ) ^ ( n16783 )  ;
assign n16856 =  { ( n16789 ) , ( n16855 ) }  ;
assign n16857 = ~ ( n3963 ) ;
assign n16858 = ~ ( n3583 ) ;
assign n16859 =  ( n3567 ) | ( n16858 )  ;
assign n16860 =  ( n16857 ) ^ ( n16859 )  ;
assign n16861 =  ( n3264 ) | ( n3274 )  ;
assign n16862 =  ( n16861 ) | ( n3288 )  ;
assign n16863 =  ( n16860 ) ^ ( n16862 )  ;
assign n16864 =  ( n16863 ) ^ ( n3303 )  ;
assign n16865 =  ( n16864 ) ^ ( n2846 )  ;
assign n16866 =  ( n16865 ) ^ ( n2856 )  ;
assign n16867 =  ( n16866 ) ^ ( n2919 )  ;
assign n16868 = ~ ( n2468 ) ;
assign n16869 =  ( n16867 ) ^ ( n16868 )  ;
assign n16870 =  ( n16869 ) ^ ( n2483 )  ;
assign n16871 =  ( n16870 ) ^ ( n2500 )  ;
assign n16872 =  ( n16871 ) ^ ( n2517 )  ;
assign n16873 =  ( n16872 ) ^ ( n2548 )  ;
assign n16874 =  ( n16873 ) ^ ( n2578 )  ;
assign n16875 =  ( n16874 ) ^ ( n2594 )  ;
assign n16876 =  ( n16875 ) ^ ( n2620 )  ;
assign n16877 =  ( n16876 ) ^ ( n13715 )  ;
assign n16878 = ~ ( n8880 ) ;
assign n16879 = ~ ( n8920 ) ;
assign n16880 =  ( n16878 ) | ( n16879 )  ;
assign n16881 = ~ ( n16880 ) ;
assign n16882 =  ( n16877 ) ^ ( n16881 )  ;
assign n16883 =  ( n16882 ) ^ ( n8541 )  ;
assign n16884 =  ( n16883 ) ^ ( n8227 )  ;
assign n16885 =  ( n16884 ) ^ ( n8233 )  ;
assign n16886 = ~ ( n7779 ) ;
assign n16887 =  ( n7784 ) | ( n6524 )  ;
assign n16888 = ~ ( n16887 ) ;
assign n16889 =  ( n16886 ) | ( n16888 )  ;
assign n16890 = ~ ( n7801 ) ;
assign n16891 =  ( n16889 ) | ( n16890 )  ;
assign n16892 =  ( n16885 ) ^ ( n16891 )  ;
assign n16893 = ~ ( n7809 ) ;
assign n16894 = ~ ( n6553 ) ;
assign n16895 =  ( n16893 ) | ( n16894 )  ;
assign n16896 =  ( n16892 ) ^ ( n16895 )  ;
assign n16897 = ~ ( n5902 ) ;
assign n16898 = ~ ( n5913 ) ;
assign n16899 =  ( n16897 ) | ( n16898 )  ;
assign n16900 =  ( n16896 ) ^ ( n16899 )  ;
assign n16901 = ~ ( n7455 ) ;
assign n16902 =  ( n16900 ) ^ ( n16901 )  ;
assign n16903 =  ( n6825 ) | ( n6834 )  ;
assign n16904 =  ( n16903 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n16905 =  ( n16902 ) ^ ( n16904 )  ;
assign n16906 =  ( n6483 ) | ( n6492 )  ;
assign n16907 =  ( n16906 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n16908 =  ( n16905 ) ^ ( n16907 )  ;
assign n16909 =  ( n6030 ) | ( n6039 )  ;
assign n16910 =  ( n16909 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16911 =  ( n16908 ) ^ ( n16910 )  ;
assign n16912 =  ( n5802 ) | ( n5811 )  ;
assign n16913 =  ( n16912 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16914 =  ( n16911 ) ^ ( n16913 )  ;
assign n16915 =  ( n5832 ) | ( n5841 )  ;
assign n16916 =  ( n16915 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16917 =  ( n16914 ) ^ ( n16916 )  ;
assign n16918 =  ( n5682 ) | ( n5691 )  ;
assign n16919 =  ( n16918 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16920 =  ( n16917 ) ^ ( n16919 )  ;
assign n16921 =  ( n5713 ) | ( n5722 )  ;
assign n16922 =  ( n16921 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16923 =  ( n16920 ) ^ ( n16922 )  ;
assign n16924 =  ( n16923 ) ^ ( n13774 )  ;
assign n16925 = ~ ( n13914 ) ;
assign n16926 =  ( n13867 ) | ( n16925 )  ;
assign n16927 = ~ ( n16926 ) ;
assign n16928 = ~ ( n14019 ) ;
assign n16929 = ~ ( n15291 ) ;
assign n16930 =  ( n16928 ) | ( n16929 )  ;
assign n16931 = ~ ( n16930 ) ;
assign n16932 =  ( n16927 ) | ( n16931 )  ;
assign n16933 =  ( n16924 ) ^ ( n16932 )  ;
assign n16934 =  { ( n16856 ) , ( n16933 ) }  ;
assign n16935 = ~ ( n3918 ) ;
assign n16936 =  ( n3902 ) | ( n16935 )  ;
assign n16937 =  ( n4234 ) ^ ( n16936 )  ;
assign n16938 =  ( n3519 ) | ( n3531 )  ;
assign n16939 =  ( n16938 ) | ( n3547 )  ;
assign n16940 =  ( n16937 ) ^ ( n16939 )  ;
assign n16941 =  ( n16940 ) ^ ( n3564 )  ;
assign n16942 =  ( n16941 ) ^ ( n3189 )  ;
assign n16943 =  ( n16942 ) ^ ( n3199 )  ;
assign n16944 =  ( n16943 ) ^ ( n3255 )  ;
assign n16945 =  ( n16944 ) ^ ( n2763 )  ;
assign n16946 =  ( n16945 ) ^ ( n2779 )  ;
assign n16947 =  ( n16946 ) ^ ( n2796 )  ;
assign n16948 =  ( n16947 ) ^ ( n2813 )  ;
assign n16949 =  ( n16948 ) ^ ( n2842 )  ;
assign n16950 =  ( n16949 ) ^ ( n2873 )  ;
assign n16951 =  ( n16950 ) ^ ( n2889 )  ;
assign n16952 =  ( n16951 ) ^ ( n2915 )  ;
assign n16953 =  ( n16952 ) ^ ( n5668 )  ;
assign n16954 = ~ ( n9088 ) ;
assign n16955 = ~ ( n9126 ) ;
assign n16956 =  ( n16954 ) | ( n16955 )  ;
assign n16957 = ~ ( n16956 ) ;
assign n16958 =  ( n16953 ) ^ ( n16957 )  ;
assign n16959 =  ( n16958 ) ^ ( n8880 )  ;
assign n16960 =  ( n16959 ) ^ ( n8490 )  ;
assign n16961 = ~ ( n7905 ) ;
assign n16962 =  ( n8179 ) | ( n8427 )  ;
assign n16963 = ~ ( n16962 ) ;
assign n16964 =  ( n16961 ) | ( n16963 )  ;
assign n16965 =  ( n16960 ) ^ ( n16964 )  ;
assign n16966 = ~ ( n7779 ) ;
assign n16967 =  ( n7784 ) | ( n6524 )  ;
assign n16968 = ~ ( n16967 ) ;
assign n16969 =  ( n16966 ) | ( n16968 )  ;
assign n16970 = ~ ( n7801 ) ;
assign n16971 =  ( n16969 ) | ( n16970 )  ;
assign n16972 =  ( n16965 ) ^ ( n16971 )  ;
assign n16973 = ~ ( n7809 ) ;
assign n16974 = ~ ( n6553 ) ;
assign n16975 =  ( n16973 ) | ( n16974 )  ;
assign n16976 =  ( n16972 ) ^ ( n16975 )  ;
assign n16977 =  ( n16976 ) ^ ( n8164 )  ;
assign n16978 =  ( n16977 ) ^ ( n7455 )  ;
assign n16979 =  ( n6825 ) | ( n6834 )  ;
assign n16980 =  ( n16979 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n16981 =  ( n16978 ) ^ ( n16980 )  ;
assign n16982 =  ( n6483 ) | ( n6492 )  ;
assign n16983 =  ( n16982 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n16984 =  ( n16981 ) ^ ( n16983 )  ;
assign n16985 =  ( n6030 ) | ( n6039 )  ;
assign n16986 =  ( n16985 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n16987 =  ( n16984 ) ^ ( n16986 )  ;
assign n16988 =  ( n5802 ) | ( n5811 )  ;
assign n16989 =  ( n16988 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n16990 =  ( n16987 ) ^ ( n16989 )  ;
assign n16991 =  ( n5832 ) | ( n5841 )  ;
assign n16992 =  ( n16991 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n16993 =  ( n16990 ) ^ ( n16992 )  ;
assign n16994 =  ( n5682 ) | ( n5691 )  ;
assign n16995 =  ( n16994 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n16996 =  ( n16993 ) ^ ( n16995 )  ;
assign n16997 =  ( n5713 ) | ( n5722 )  ;
assign n16998 =  ( n16997 ) ? ( bv_1_0_n2 ) : ( n5733 ) ;
assign n16999 =  ( n16996 ) ^ ( n16998 )  ;
assign n17000 =  ( n16999 ) ^ ( n10575 )  ;
assign n17001 =  ( n17000 ) ^ ( n15291 )  ;
assign n17002 =  { ( n16934 ) , ( n17001 ) }  ;
assign n17003 =  ( n4123 ) | ( n4142 )  ;
assign n17004 =  ( n4440 ) ^ ( n17003 )  ;
assign n17005 =  ( n3856 ) | ( n3866 )  ;
assign n17006 =  ( n17005 ) | ( n3884 )  ;
assign n17007 =  ( n17004 ) ^ ( n17006 )  ;
assign n17008 =  ( n17007 ) ^ ( n3899 )  ;
assign n17009 =  ( n17008 ) ^ ( n3496 )  ;
assign n17010 =  ( n17009 ) ^ ( n3506 )  ;
assign n17011 =  ( n17010 ) ^ ( n3106 )  ;
assign n17012 =  ( n17011 ) ^ ( n3122 )  ;
assign n17013 =  ( n17012 ) ^ ( n3139 )  ;
assign n17014 =  ( n17013 ) ^ ( n3156 )  ;
assign n17015 =  ( n17014 ) ^ ( n3185 )  ;
assign n17016 =  ( n17015 ) ^ ( n3216 )  ;
assign n17017 =  ( n17016 ) ^ ( n3232 )  ;
assign n17018 =  ( n17017 ) ^ ( n3251 )  ;
assign n17019 =  ( n17018 ) ^ ( n3248 )  ;
assign n17020 =  ( n17019 ) ^ ( n14048 )  ;
assign n17021 = ~ ( n9314 ) ;
assign n17022 = ~ ( n9348 ) ;
assign n17023 =  ( n17021 ) | ( n17022 )  ;
assign n17024 = ~ ( n17023 ) ;
assign n17025 =  ( n17020 ) ^ ( n17024 )  ;
assign n17026 =  ( n17025 ) ^ ( n9088 )  ;
assign n17027 =  ( n17026 ) ^ ( n8829 )  ;
assign n17028 = ~ ( n7905 ) ;
assign n17029 = ~ ( n8835 ) ;
assign n17030 =  ( n17028 ) | ( n17029 )  ;
assign n17031 =  ( n17027 ) ^ ( n17030 )  ;
assign n17032 = ~ ( n7779 ) ;
assign n17033 =  ( n7784 ) | ( n6524 )  ;
assign n17034 = ~ ( n17033 ) ;
assign n17035 =  ( n17032 ) | ( n17034 )  ;
assign n17036 = ~ ( n7801 ) ;
assign n17037 =  ( n17035 ) | ( n17036 )  ;
assign n17038 =  ( n17031 ) ^ ( n17037 )  ;
assign n17039 = ~ ( n7809 ) ;
assign n17040 = ~ ( n6553 ) ;
assign n17041 =  ( n17039 ) | ( n17040 )  ;
assign n17042 =  ( n17038 ) ^ ( n17041 )  ;
assign n17043 =  ( n17042 ) ^ ( n7455 )  ;
assign n17044 =  ( n6825 ) | ( n6834 )  ;
assign n17045 =  ( n17044 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17046 =  ( n17043 ) ^ ( n17045 )  ;
assign n17047 =  ( n6483 ) | ( n6492 )  ;
assign n17048 =  ( n17047 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17049 =  ( n17046 ) ^ ( n17048 )  ;
assign n17050 =  ( n6030 ) | ( n6039 )  ;
assign n17051 =  ( n17050 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17052 =  ( n17049 ) ^ ( n17051 )  ;
assign n17053 =  ( n5802 ) | ( n5811 )  ;
assign n17054 =  ( n17053 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n17055 =  ( n17052 ) ^ ( n17054 )  ;
assign n17056 =  ( n5832 ) | ( n5841 )  ;
assign n17057 =  ( n17056 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n17058 =  ( n17055 ) ^ ( n17057 )  ;
assign n17059 =  ( n5682 ) | ( n5691 )  ;
assign n17060 =  ( n17059 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n17061 =  ( n17058 ) ^ ( n17060 )  ;
assign n17062 =  ( n17061 ) ^ ( n8160 )  ;
assign n17063 =  ( n17062 ) ^ ( n8157 )  ;
assign n17064 =  ( n17063 ) ^ ( n14103 )  ;
assign n17065 = ~ ( n14227 ) ;
assign n17066 =  ( n14186 ) | ( n17065 )  ;
assign n17067 = ~ ( n17066 ) ;
assign n17068 = ~ ( n14288 ) ;
assign n17069 = ~ ( n15568 ) ;
assign n17070 =  ( n17068 ) | ( n17069 )  ;
assign n17071 = ~ ( n17070 ) ;
assign n17072 =  ( n17067 ) | ( n17071 )  ;
assign n17073 =  ( n17064 ) ^ ( n17072 )  ;
assign n17074 =  { ( n17002 ) , ( n17073 ) }  ;
assign n17075 = ~ ( n4695 ) ;
assign n17076 =  ( n4390 ) | ( n4403 )  ;
assign n17077 =  ( n17075 ) ^ ( n17076 )  ;
assign n17078 =  ( n17077 ) ^ ( n4111 )  ;
assign n17079 =  ( n17078 ) ^ ( n3776 )  ;
assign n17080 =  ( n17079 ) ^ ( n3786 )  ;
assign n17081 =  ( n17080 ) ^ ( n3847 )  ;
assign n17082 =  ( n17081 ) ^ ( n3413 )  ;
assign n17083 =  ( n17082 ) ^ ( n3429 )  ;
assign n17084 =  ( n17083 ) ^ ( n3446 )  ;
assign n17085 =  ( n17084 ) ^ ( n3463 )  ;
assign n17086 =  ( n17085 ) ^ ( n3492 )  ;
assign n17087 =  ( n17086 ) ^ ( n3881 )  ;
assign n17088 =  ( n17087 ) ^ ( n4139 )  ;
assign n17089 =  ( n17088 ) ^ ( n10841 )  ;
assign n17090 = ~ ( n9538 ) ;
assign n17091 = ~ ( n9569 ) ;
assign n17092 =  ( n17090 ) | ( n17091 )  ;
assign n17093 = ~ ( n17092 ) ;
assign n17094 =  ( n17089 ) ^ ( n17093 )  ;
assign n17095 =  ( n17094 ) ^ ( n9314 )  ;
assign n17096 =  ( n17095 ) ^ ( n9018 )  ;
assign n17097 = ~ ( n7779 ) ;
assign n17098 =  ( n7784 ) | ( n6524 )  ;
assign n17099 = ~ ( n17098 ) ;
assign n17100 =  ( n17097 ) | ( n17099 )  ;
assign n17101 = ~ ( n7801 ) ;
assign n17102 =  ( n17100 ) | ( n17101 )  ;
assign n17103 =  ( n17096 ) ^ ( n17102 )  ;
assign n17104 = ~ ( n7809 ) ;
assign n17105 = ~ ( n6553 ) ;
assign n17106 =  ( n17104 ) | ( n17105 )  ;
assign n17107 =  ( n17103 ) ^ ( n17106 )  ;
assign n17108 = ~ ( n8761 ) ;
assign n17109 =  ( n17108 ) | ( n8771 )  ;
assign n17110 =  ( n17107 ) ^ ( n17109 )  ;
assign n17111 =  ( n17110 ) ^ ( n7455 )  ;
assign n17112 =  ( n6825 ) | ( n6834 )  ;
assign n17113 =  ( n17112 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17114 =  ( n17111 ) ^ ( n17113 )  ;
assign n17115 =  ( n6483 ) | ( n6492 )  ;
assign n17116 =  ( n17115 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17117 =  ( n17114 ) ^ ( n17116 )  ;
assign n17118 =  ( n6030 ) | ( n6039 )  ;
assign n17119 =  ( n17118 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17120 =  ( n17117 ) ^ ( n17119 )  ;
assign n17121 =  ( n5802 ) | ( n5811 )  ;
assign n17122 =  ( n17121 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n17123 =  ( n17120 ) ^ ( n17122 )  ;
assign n17124 =  ( n5832 ) | ( n5841 )  ;
assign n17125 =  ( n17124 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n17126 =  ( n17123 ) ^ ( n17125 )  ;
assign n17127 =  ( n5682 ) | ( n5691 )  ;
assign n17128 =  ( n17127 ) ? ( bv_1_0_n2 ) : ( n5702 ) ;
assign n17129 =  ( n17126 ) ^ ( n17128 )  ;
assign n17130 =  ( n17129 ) ^ ( n11090 )  ;
assign n17131 =  ( n17130 ) ^ ( n15568 )  ;
assign n17132 =  { ( n17074 ) , ( n17131 ) }  ;
assign n17133 = ~ ( n4728 ) ;
assign n17134 =  ( n4722 ) | ( n17133 )  ;
assign n17135 = ~ ( n17134 ) ;
assign n17136 = ~ ( n4659 ) ;
assign n17137 =  ( n4647 ) | ( n17136 )  ;
assign n17138 =  ( n17135 ) ^ ( n17137 )  ;
assign n17139 =  ( n17138 ) ^ ( n4380 )  ;
assign n17140 =  ( n17139 ) ^ ( n4088 )  ;
assign n17141 =  ( n17140 ) ^ ( n4098 )  ;
assign n17142 =  ( n17141 ) ^ ( n3693 )  ;
assign n17143 =  ( n17142 ) ^ ( n3709 )  ;
assign n17144 =  ( n17143 ) ^ ( n3726 )  ;
assign n17145 =  ( n17144 ) ^ ( n3743 )  ;
assign n17146 =  ( n17145 ) ^ ( n3772 )  ;
assign n17147 =  ( n17146 ) ^ ( n3812 )  ;
assign n17148 =  ( n17147 ) ^ ( n3836 )  ;
assign n17149 =  ( n17148 ) ^ ( n3824 )  ;
assign n17150 =  ( n17149 ) ^ ( n14320 )  ;
assign n17151 = ~ ( n9719 ) ;
assign n17152 =  ( n17150 ) ^ ( n17151 )  ;
assign n17153 =  ( n17152 ) ^ ( n9538 )  ;
assign n17154 =  ( n17153 ) ^ ( n9018 )  ;
assign n17155 = ~ ( n7779 ) ;
assign n17156 =  ( n7784 ) | ( n6524 )  ;
assign n17157 = ~ ( n17156 ) ;
assign n17158 =  ( n17155 ) | ( n17157 )  ;
assign n17159 = ~ ( n7801 ) ;
assign n17160 =  ( n17158 ) | ( n17159 )  ;
assign n17161 =  ( n17154 ) ^ ( n17160 )  ;
assign n17162 = ~ ( n7809 ) ;
assign n17163 = ~ ( n6553 ) ;
assign n17164 =  ( n17162 ) | ( n17163 )  ;
assign n17165 =  ( n17161 ) ^ ( n17164 )  ;
assign n17166 =  ( n17165 ) ^ ( n7455 )  ;
assign n17167 =  ( n6825 ) | ( n6834 )  ;
assign n17168 =  ( n17167 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17169 =  ( n17166 ) ^ ( n17168 )  ;
assign n17170 =  ( n6483 ) | ( n6492 )  ;
assign n17171 =  ( n17170 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17172 =  ( n17169 ) ^ ( n17171 )  ;
assign n17173 =  ( n6030 ) | ( n6039 )  ;
assign n17174 =  ( n17173 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17175 =  ( n17172 ) ^ ( n17174 )  ;
assign n17176 =  ( n5802 ) | ( n5811 )  ;
assign n17177 =  ( n17176 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n17178 =  ( n17175 ) ^ ( n17177 )  ;
assign n17179 =  ( n5832 ) | ( n5841 )  ;
assign n17180 =  ( n17179 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n17181 =  ( n17178 ) ^ ( n17180 )  ;
assign n17182 =  ( n17181 ) ^ ( n8759 )  ;
assign n17183 =  ( n17182 ) ^ ( n8756 )  ;
assign n17184 =  ( n17183 ) ^ ( n14364 )  ;
assign n17185 = ~ ( n14441 ) ;
assign n17186 = ~ ( n14476 ) ;
assign n17187 =  ( n17185 ) | ( n17186 )  ;
assign n17188 = ~ ( n17187 ) ;
assign n17189 = ~ ( n14543 ) ;
assign n17190 = ~ ( n15802 ) ;
assign n17191 =  ( n17189 ) | ( n17190 )  ;
assign n17192 = ~ ( n17191 ) ;
assign n17193 =  ( n17188 ) | ( n17192 )  ;
assign n17194 =  ( n17184 ) ^ ( n17193 )  ;
assign n17195 =  { ( n17132 ) , ( n17194 ) }  ;
assign n17196 = ~ ( n4889 ) ;
assign n17197 =  ( n17196 ) | ( n4900 )  ;
assign n17198 = ~ ( n17197 ) ;
assign n17199 =  ( n4605 ) | ( n4615 )  ;
assign n17200 =  ( n17199 ) | ( n4629 )  ;
assign n17201 =  ( n17198 ) ^ ( n17200 )  ;
assign n17202 =  ( n17201 ) ^ ( n4644 )  ;
assign n17203 =  ( n17202 ) ^ ( n4357 )  ;
assign n17204 =  ( n17203 ) ^ ( n4367 )  ;
assign n17205 =  ( n17204 ) ^ ( n4005 )  ;
assign n17206 =  ( n17205 ) ^ ( n4021 )  ;
assign n17207 =  ( n17206 ) ^ ( n4038 )  ;
assign n17208 =  ( n17207 ) ^ ( n4055 )  ;
assign n17209 =  ( n17208 ) ^ ( n4084 )  ;
assign n17210 =  ( n17209 ) ^ ( n4728 )  ;
assign n17211 =  ( n5041 ) | ( n5203 )  ;
assign n17212 =  ( n17211 ) | ( n5345 )  ;
assign n17213 =  ( n17212 ) | ( n11288 )  ;
assign n17214 =  ( n17213 ) | ( n11331 )  ;
assign n17215 =  ( n17210 ) ^ ( n17214 )  ;
assign n17216 = ~ ( n9834 ) ;
assign n17217 =  ( n9808 ) | ( n17216 )  ;
assign n17218 = ~ ( n17217 ) ;
assign n17219 =  ( n17215 ) ^ ( n17218 )  ;
assign n17220 =  ( n17219 ) ^ ( n9523 )  ;
assign n17221 =  ( n17220 ) ^ ( n9529 )  ;
assign n17222 = ~ ( n7779 ) ;
assign n17223 =  ( n7784 ) | ( n6524 )  ;
assign n17224 = ~ ( n17223 ) ;
assign n17225 =  ( n17222 ) | ( n17224 )  ;
assign n17226 = ~ ( n7801 ) ;
assign n17227 =  ( n17225 ) | ( n17226 )  ;
assign n17228 =  ( n17221 ) ^ ( n17227 )  ;
assign n17229 = ~ ( n7809 ) ;
assign n17230 = ~ ( n6553 ) ;
assign n17231 =  ( n17229 ) | ( n17230 )  ;
assign n17232 =  ( n17228 ) ^ ( n17231 )  ;
assign n17233 =  ( n17232 ) ^ ( n7455 )  ;
assign n17234 =  ( n6825 ) | ( n6834 )  ;
assign n17235 =  ( n17234 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17236 =  ( n17233 ) ^ ( n17235 )  ;
assign n17237 =  ( n6483 ) | ( n6492 )  ;
assign n17238 =  ( n17237 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17239 =  ( n17236 ) ^ ( n17238 )  ;
assign n17240 =  ( n6030 ) | ( n6039 )  ;
assign n17241 =  ( n17240 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17242 =  ( n17239 ) ^ ( n17241 )  ;
assign n17243 =  ( n5802 ) | ( n5811 )  ;
assign n17244 =  ( n17243 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n17245 =  ( n17242 ) ^ ( n17244 )  ;
assign n17246 =  ( n5832 ) | ( n5841 )  ;
assign n17247 =  ( n17246 ) ? ( bv_1_0_n2 ) : ( n5852 ) ;
assign n17248 =  ( n17245 ) ^ ( n17247 )  ;
assign n17249 =  ( n17248 ) ^ ( n11533 )  ;
assign n17250 =  ( n17249 ) ^ ( n15802 )  ;
assign n17251 =  { ( n17195 ) , ( n17250 ) }  ;
assign n17252 =  ( n5052 ) ^ ( n4889 )  ;
assign n17253 =  ( n17252 ) ^ ( n4561 )  ;
assign n17254 =  ( n17253 ) ^ ( n4571 )  ;
assign n17255 =  ( n17254 ) ^ ( n4274 )  ;
assign n17256 =  ( n17255 ) ^ ( n4290 )  ;
assign n17257 =  ( n17256 ) ^ ( n4307 )  ;
assign n17258 =  ( n17257 ) ^ ( n4324 )  ;
assign n17259 =  ( n17258 ) ^ ( n4353 )  ;
assign n17260 =  ( n17259 ) ^ ( n4602 )  ;
assign n17261 =  ( n17260 ) ^ ( n4590 )  ;
assign n17262 =  ( n14566 ) | ( n14573 )  ;
assign n17263 =  ( n17261 ) ^ ( n17262 )  ;
assign n17264 = ~ ( n10010 ) ;
assign n17265 =  ( n17263 ) ^ ( n17264 )  ;
assign n17266 = ~ ( n9798 ) ;
assign n17267 =  ( n9804 ) | ( n8179 )  ;
assign n17268 = ~ ( n17267 ) ;
assign n17269 =  ( n17266 ) | ( n17268 )  ;
assign n17270 =  ( n17265 ) ^ ( n17269 )  ;
assign n17271 = ~ ( n7779 ) ;
assign n17272 =  ( n7784 ) | ( n6524 )  ;
assign n17273 = ~ ( n17272 ) ;
assign n17274 =  ( n17271 ) | ( n17273 )  ;
assign n17275 = ~ ( n7801 ) ;
assign n17276 =  ( n17274 ) | ( n17275 )  ;
assign n17277 =  ( n17270 ) ^ ( n17276 )  ;
assign n17278 = ~ ( n7809 ) ;
assign n17279 = ~ ( n6553 ) ;
assign n17280 =  ( n17278 ) | ( n17279 )  ;
assign n17281 =  ( n17277 ) ^ ( n17280 )  ;
assign n17282 =  ( n17281 ) ^ ( n7455 )  ;
assign n17283 =  ( n6825 ) | ( n6834 )  ;
assign n17284 =  ( n17283 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17285 =  ( n17282 ) ^ ( n17284 )  ;
assign n17286 =  ( n6483 ) | ( n6492 )  ;
assign n17287 =  ( n17286 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17288 =  ( n17285 ) ^ ( n17287 )  ;
assign n17289 =  ( n6030 ) | ( n6039 )  ;
assign n17290 =  ( n17289 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17291 =  ( n17288 ) ^ ( n17290 )  ;
assign n17292 =  ( n5802 ) | ( n5811 )  ;
assign n17293 =  ( n17292 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n17294 =  ( n17291 ) ^ ( n17293 )  ;
assign n17295 =  ( n17294 ) ^ ( n9471 )  ;
assign n17296 =  ( n17295 ) ^ ( n9468 )  ;
assign n17297 =  ( n17296 ) ^ ( n14617 )  ;
assign n17298 = ~ ( n14709 ) ;
assign n17299 =  ( n14683 ) | ( n17298 )  ;
assign n17300 = ~ ( n17299 ) ;
assign n17301 = ~ ( n14754 ) ;
assign n17302 = ~ ( n16043 ) ;
assign n17303 =  ( n17301 ) | ( n17302 )  ;
assign n17304 = ~ ( n17303 ) ;
assign n17305 =  ( n17300 ) | ( n17304 )  ;
assign n17306 =  ( n17297 ) ^ ( n17305 )  ;
assign n17307 =  { ( n17251 ) , ( n17306 ) }  ;
assign n17308 =  ( n5008 ) | ( n5019 )  ;
assign n17309 =  ( n5214 ) ^ ( n17308 )  ;
assign n17310 =  ( n17309 ) ^ ( n4866 )  ;
assign n17311 =  ( n17310 ) ^ ( n4876 )  ;
assign n17312 =  ( n17311 ) ^ ( n4478 )  ;
assign n17313 =  ( n17312 ) ^ ( n4494 )  ;
assign n17314 =  ( n17313 ) ^ ( n4511 )  ;
assign n17315 =  ( n17314 ) ^ ( n4528 )  ;
assign n17316 =  ( n17315 ) ^ ( n4557 )  ;
assign n17317 =  ( n5248 ) | ( n5341 )  ;
assign n17318 =  ( n17317 ) | ( n10785 )  ;
assign n17319 =  ( n17318 ) | ( n11760 )  ;
assign n17320 =  ( n17319 ) | ( n11801 )  ;
assign n17321 =  ( n17316 ) ^ ( n17320 )  ;
assign n17322 = ~ ( n10140 ) ;
assign n17323 =  ( n17322 ) | ( n10158 )  ;
assign n17324 = ~ ( n17323 ) ;
assign n17325 =  ( n17321 ) ^ ( n17324 )  ;
assign n17326 = ~ ( n9931 ) ;
assign n17327 =  ( n17326 ) | ( n9952 )  ;
assign n17328 =  ( n17325 ) ^ ( n17327 )  ;
assign n17329 =  ( n17328 ) ^ ( n9792 )  ;
assign n17330 = ~ ( n7809 ) ;
assign n17331 = ~ ( n6553 ) ;
assign n17332 =  ( n17330 ) | ( n17331 )  ;
assign n17333 =  ( n17329 ) ^ ( n17332 )  ;
assign n17334 =  ( n17333 ) ^ ( n7455 )  ;
assign n17335 =  ( n6825 ) | ( n6834 )  ;
assign n17336 =  ( n17335 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17337 =  ( n17334 ) ^ ( n17336 )  ;
assign n17338 =  ( n6483 ) | ( n6492 )  ;
assign n17339 =  ( n17338 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17340 =  ( n17337 ) ^ ( n17339 )  ;
assign n17341 =  ( n6030 ) | ( n6039 )  ;
assign n17342 =  ( n17341 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17343 =  ( n17340 ) ^ ( n17342 )  ;
assign n17344 =  ( n5802 ) | ( n5811 )  ;
assign n17345 =  ( n17344 ) ? ( bv_1_0_n2 ) : ( n5822 ) ;
assign n17346 =  ( n17343 ) ^ ( n17345 )  ;
assign n17347 =  ( n17346 ) ^ ( n11992 )  ;
assign n17348 =  ( n17347 ) ^ ( n16043 )  ;
assign n17349 =  { ( n17307 ) , ( n17348 ) }  ;
assign n17350 =  ( n5256 ) ^ ( n5182 )  ;
assign n17351 =  ( n17350 ) ^ ( n5000 )  ;
assign n17352 =  ( n17351 ) ^ ( n4784 )  ;
assign n17353 =  ( n17352 ) ^ ( n4800 )  ;
assign n17354 =  ( n17353 ) ^ ( n4817 )  ;
assign n17355 =  ( n17354 ) ^ ( n4834 )  ;
assign n17356 =  ( n17355 ) ^ ( n4862 )  ;
assign n17357 =  ( n17356 ) ^ ( n4859 )  ;
assign n17358 =  ( n14779 ) | ( n14792 )  ;
assign n17359 =  ( n17357 ) ^ ( n17358 )  ;
assign n17360 = ~ ( n10255 ) ;
assign n17361 =  ( n17359 ) ^ ( n17360 )  ;
assign n17362 =  ( n17361 ) ^ ( n10140 )  ;
assign n17363 = ~ ( n7809 ) ;
assign n17364 = ~ ( n9916 ) ;
assign n17365 =  ( n17363 ) | ( n17364 )  ;
assign n17366 =  ( n17362 ) ^ ( n17365 )  ;
assign n17367 =  ( n17366 ) ^ ( n7455 )  ;
assign n17368 =  ( n6825 ) | ( n6834 )  ;
assign n17369 =  ( n17368 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17370 =  ( n17367 ) ^ ( n17369 )  ;
assign n17371 =  ( n6483 ) | ( n6492 )  ;
assign n17372 =  ( n17371 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17373 =  ( n17370 ) ^ ( n17372 )  ;
assign n17374 =  ( n6030 ) | ( n6039 )  ;
assign n17375 =  ( n17374 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17376 =  ( n17373 ) ^ ( n17375 )  ;
assign n17377 =  ( n17376 ) ^ ( n9788 )  ;
assign n17378 =  ( n17377 ) ^ ( n9785 )  ;
assign n17379 =  ( n17378 ) ^ ( n14826 )  ;
assign n17380 = ~ ( n14895 ) ;
assign n17381 =  ( n14872 ) | ( n17380 )  ;
assign n17382 = ~ ( n17381 ) ;
assign n17383 = ~ ( n14952 ) ;
assign n17384 = ~ ( n15287 ) ;
assign n17385 =  ( n17383 ) | ( n17384 )  ;
assign n17386 = ~ ( n17385 ) ;
assign n17387 =  ( n17382 ) | ( n17386 )  ;
assign n17388 =  ( n17379 ) ^ ( n17387 )  ;
assign n17389 =  { ( n17349 ) , ( n17388 ) }  ;
assign n17390 =  ( n5366 ) ^ ( n5161 )  ;
assign n17391 =  ( n17390 ) ^ ( n5171 )  ;
assign n17392 =  ( n17391 ) ^ ( n4960 )  ;
assign n17393 =  ( n17392 ) ^ ( n4976 )  ;
assign n17394 =  ( n17393 ) ^ ( n4996 )  ;
assign n17395 =  ( n17394 ) ^ ( n5236 )  ;
assign n17396 =  ( n5446 ) | ( n5473 )  ;
assign n17397 =  ( n17396 ) | ( n5604 )  ;
assign n17398 =  ( n17397 ) | ( n5663 )  ;
assign n17399 =  ( n17395 ) ^ ( n17398 )  ;
assign n17400 = ~ ( n10337 ) ;
assign n17401 =  ( n17399 ) ^ ( n17400 )  ;
assign n17402 = ~ ( n10086 ) ;
assign n17403 =  ( n7784 ) | ( n10091 )  ;
assign n17404 = ~ ( n17403 ) ;
assign n17405 =  ( n17402 ) | ( n17404 )  ;
assign n17406 =  ( n17405 ) | ( n10107 )  ;
assign n17407 =  ( n17401 ) ^ ( n17406 )  ;
assign n17408 = ~ ( n7809 ) ;
assign n17409 = ~ ( n10115 ) ;
assign n17410 =  ( n17408 ) | ( n17409 )  ;
assign n17411 =  ( n17407 ) ^ ( n17410 )  ;
assign n17412 =  ( n17411 ) ^ ( n7455 )  ;
assign n17413 =  ( n6825 ) | ( n6834 )  ;
assign n17414 =  ( n17413 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17415 =  ( n17412 ) ^ ( n17414 )  ;
assign n17416 =  ( n6483 ) | ( n6492 )  ;
assign n17417 =  ( n17416 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17418 =  ( n17415 ) ^ ( n17417 )  ;
assign n17419 =  ( n6030 ) | ( n6039 )  ;
assign n17420 =  ( n17419 ) ? ( bv_1_0_n2 ) : ( n6050 ) ;
assign n17421 =  ( n17418 ) ^ ( n17420 )  ;
assign n17422 =  ( n17421 ) ^ ( n10571 )  ;
assign n17423 =  ( n17422 ) ^ ( n15287 )  ;
assign n17424 =  { ( n17389 ) , ( n17423 ) }  ;
assign n17425 =  ( n5452 ) ^ ( n5325 )  ;
assign n17426 =  ( n17425 ) ^ ( n5083 )  ;
assign n17427 =  ( n17426 ) ^ ( n5099 )  ;
assign n17428 =  ( n17427 ) ^ ( n5116 )  ;
assign n17429 =  ( n17428 ) ^ ( n5141 )  ;
assign n17430 =  ( n17429 ) ^ ( n5129 )  ;
assign n17431 =  ( n14973 ) | ( n14983 )  ;
assign n17432 =  ( n17430 ) ^ ( n17431 )  ;
assign n17433 = ~ ( n10397 ) ;
assign n17434 =  ( n17433 ) | ( n10137 )  ;
assign n17435 = ~ ( n17434 ) ;
assign n17436 =  ( n17432 ) ^ ( n17435 )  ;
assign n17437 = ~ ( n7809 ) ;
assign n17438 = ~ ( n9916 ) ;
assign n17439 =  ( n17437 ) | ( n17438 )  ;
assign n17440 =  ( n17436 ) ^ ( n17439 )  ;
assign n17441 =  ( n17440 ) ^ ( n7455 )  ;
assign n17442 =  ( n6825 ) | ( n6834 )  ;
assign n17443 =  ( n17442 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17444 =  ( n17441 ) ^ ( n17443 )  ;
assign n17445 =  ( n6483 ) | ( n6492 )  ;
assign n17446 =  ( n17445 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17447 =  ( n17444 ) ^ ( n17446 )  ;
assign n17448 =  ( n17447 ) ^ ( n10084 )  ;
assign n17449 =  ( n17448 ) ^ ( n10081 )  ;
assign n17450 =  ( n17449 ) ^ ( n15012 )  ;
assign n17451 =  ( n15051 ) | ( n15062 )  ;
assign n17452 = ~ ( n17451 ) ;
assign n17453 = ~ ( n15564 ) ;
assign n17454 =  ( n15084 ) | ( n17453 )  ;
assign n17455 = ~ ( n17454 ) ;
assign n17456 =  ( n17452 ) | ( n17455 )  ;
assign n17457 =  ( n17450 ) ^ ( n17456 )  ;
assign n17458 =  { ( n17424 ) , ( n17457 ) }  ;
assign n17459 =  ( n5489 ) ^ ( n5433 )  ;
assign n17460 =  ( n17459 ) ^ ( n5285 )  ;
assign n17461 =  ( n17460 ) ^ ( n5301 )  ;
assign n17462 =  ( n17461 ) ^ ( n5321 )  ;
assign n17463 =  ( n5539 ) | ( n5600 )  ;
assign n17464 =  ( n17463 ) | ( n10836 )  ;
assign n17465 =  ( n17462 ) ^ ( n17464 )  ;
assign n17466 =  ( n17465 ) ^ ( n10458 )  ;
assign n17467 =  ( n17466 ) ^ ( n10397 )  ;
assign n17468 =  ( n17467 ) ^ ( n7455 )  ;
assign n17469 =  ( n6825 ) | ( n6834 )  ;
assign n17470 =  ( n17469 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17471 =  ( n17468 ) ^ ( n17470 )  ;
assign n17472 =  ( n6483 ) | ( n6492 )  ;
assign n17473 =  ( n17472 ) ? ( bv_1_0_n2 ) : ( n6503 ) ;
assign n17474 =  ( n17471 ) ^ ( n17473 )  ;
assign n17475 =  ( n17474 ) ^ ( n11086 )  ;
assign n17476 =  ( n17475 ) ^ ( n15564 )  ;
assign n17477 =  { ( n17458 ) , ( n17476 ) }  ;
assign n17478 = ~ ( n5515 ) ;
assign n17479 = ~ ( n5531 ) ;
assign n17480 =  ( n17478 ) | ( n17479 )  ;
assign n17481 = ~ ( n17480 ) ;
assign n17482 =  ( n17481 ) ^ ( n5394 )  ;
assign n17483 =  ( n17482 ) ^ ( n5410 )  ;
assign n17484 =  ( n17483 ) ^ ( n5429 )  ;
assign n17485 =  ( n17484 ) ^ ( n5426 )  ;
assign n17486 =  ( n15098 ) | ( n15113 )  ;
assign n17487 =  ( n17485 ) ^ ( n17486 )  ;
assign n17488 = ~ ( n7809 ) ;
assign n17489 =  ( n17487 ) ^ ( n17488 )  ;
assign n17490 =  ( n17489 ) ^ ( n7455 )  ;
assign n17491 =  ( n6825 ) | ( n6834 )  ;
assign n17492 =  ( n17491 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17493 =  ( n17490 ) ^ ( n17492 )  ;
assign n17494 =  ( n17493 ) ^ ( n10393 )  ;
assign n17495 =  ( n17494 ) ^ ( n10390 )  ;
assign n17496 =  ( n17495 ) ^ ( n15139 )  ;
assign n17497 =  ( n5594 ) ^ ( n5515 )  ;
assign n17498 =  ( n17497 ) ^ ( n5531 )  ;
assign n17499 =  ( n17498 ) ^ ( n15176 )  ;
assign n17500 = ~ ( n17499 ) ;
assign n17501 =  ( n17500 ) | ( n15196 )  ;
assign n17502 = ~ ( n17501 ) ;
assign n17503 =  ( n15242 ) | ( n15267 )  ;
assign n17504 = ~ ( n15281 ) ;
assign n17505 =  ( n17503 ) | ( n17504 )  ;
assign n17506 = ~ ( n17505 ) ;
assign n17507 =  ( n15217 ) | ( n17506 )  ;
assign n17508 = ~ ( n17507 ) ;
assign n17509 =  ( n17502 ) | ( n17508 )  ;
assign n17510 =  ( n17496 ) ^ ( n17509 )  ;
assign n17511 =  { ( n17477 ) , ( n17510 ) }  ;
assign n17512 =  ( n5594 ) ^ ( n5515 )  ;
assign n17513 =  ( n17512 ) ^ ( n5531 )  ;
assign n17514 =  ( n17513 ) ^ ( n15176 )  ;
assign n17515 =  ( n17514 ) ^ ( n10533 )  ;
assign n17516 =  ( n17515 ) ^ ( n7455 )  ;
assign n17517 =  ( n6825 ) | ( n6834 )  ;
assign n17518 =  ( n17517 ) ? ( bv_1_0_n2 ) : ( n6845 ) ;
assign n17519 =  ( n17516 ) ^ ( n17518 )  ;
assign n17520 =  ( n17519 ) ^ ( n15194 )  ;
assign n17521 =  ( n15242 ) | ( n15267 )  ;
assign n17522 = ~ ( n15281 ) ;
assign n17523 =  ( n17521 ) | ( n17522 )  ;
assign n17524 =  ( n17520 ) ^ ( n17523 )  ;
assign n17525 =  { ( n17511 ) , ( n17524 ) }  ;
assign n17526 =  ( n5568 ) ^ ( n5583 )  ;
assign n17527 =  ( n17526 ) ^ ( n5580 )  ;
assign n17528 =  ( n17527 ) ^ ( n15227 )  ;
assign n17529 =  ( n17528 ) ^ ( n7455 )  ;
assign n17530 =  ( n17529 ) ^ ( n10522 )  ;
assign n17531 =  ( n17530 ) ^ ( n10519 )  ;
assign n17532 =  ( n17531 ) ^ ( n15238 )  ;
assign n17533 =  ( n5648 ) ^ ( n15255 )  ;
assign n17534 = ~ ( n17533 ) ;
assign n17535 =  ( n7455 ) ^ ( n15263 )  ;
assign n17536 = ~ ( n17535 ) ;
assign n17537 =  ( n17534 ) | ( n17536 )  ;
assign n17538 = ~ ( n17537 ) ;
assign n17539 =  ( n5648 ) ^ ( n15255 )  ;
assign n17540 =  ( n17539 ) ^ ( n7455 )  ;
assign n17541 =  ( n17540 ) ^ ( n15263 )  ;
assign n17542 = ~ ( n17541 ) ;
assign n17543 = ki[1:1] ;
assign n17544 =  ( n5657 ) ^ ( n17543 )  ;
assign n17545 = ~ ( n17544 ) ;
assign n17546 =  ( n17542 ) | ( n17545 )  ;
assign n17547 = kd[1:1] ;
assign n17548 =  ( n10564 ) ^ ( n17547 )  ;
assign n17549 = ~ ( n17548 ) ;
assign n17550 =  ( n17546 ) | ( n17549 )  ;
assign n17551 = ~ ( n17550 ) ;
assign n17552 =  ( n17538 ) | ( n17551 )  ;
assign n17553 =  ( n17532 ) ^ ( n17552 )  ;
assign n17554 =  { ( n17525 ) , ( n17553 ) }  ;
assign n17555 =  ( n5648 ) ^ ( n15255 )  ;
assign n17556 =  ( n17555 ) ^ ( n7455 )  ;
assign n17557 =  ( n17556 ) ^ ( n15263 )  ;
assign n17558 = ki[1:1] ;
assign n17559 =  ( n5657 ) ^ ( n17558 )  ;
assign n17560 = ~ ( n17559 ) ;
assign n17561 = kd[1:1] ;
assign n17562 =  ( n10564 ) ^ ( n17561 )  ;
assign n17563 = ~ ( n17562 ) ;
assign n17564 =  ( n17560 ) | ( n17563 )  ;
assign n17565 = ~ ( n17564 ) ;
assign n17566 =  ( n17557 ) ^ ( n17565 )  ;
assign n17567 =  { ( n17554 ) , ( n17566 ) }  ;
assign n17568 = ki[1:1] ;
assign n17569 =  ( n5657 ) ^ ( n17568 )  ;
assign n17570 =  ( n17569 ) ^ ( n10564 )  ;
assign n17571 = kd[1:1] ;
assign n17572 =  ( n17570 ) ^ ( n17571 )  ;
assign n17573 =  { ( n17567 ) , ( n17572 ) }  ;
always @(posedge clk) begin
   if(rst) begin
       __COUNTER_start__n0 <= 0;
   end
   else if(__ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           i_wb_data <= i_wb_data ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           kp <= kp ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           ki <= ki ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           kd <= kd ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           sp <= sp ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           pv <= pv ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           RS <= RS ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           un <= n17573 ;
       end
   end
end
endmodule
