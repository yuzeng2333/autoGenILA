module NV_BLKBOX_SRC0(Y);
  (* src = "./vmod/vlibs/NV_BLKBOX_SRC0.v:12" *)
  output Y;
  assign Y = 1'b0;
endmodule
