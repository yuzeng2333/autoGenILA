module SDP_Y_CORE_cfg_mul_prelu_rsc_triosy_obj_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:816" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:817" *)
  output outsig;
  assign outsig = in_0;
endmodule
