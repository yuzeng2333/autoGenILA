module color_to_memory(color_depth_i, color_i, x_lsb_i, mem_o, sel_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire [3:0] _13_;
  wire [3:0] _14_;
  wire [3:0] _15_;
  wire [3:0] _16_;
  wire [3:0] _17_;
  wire [31:0] _18_;
  wire [31:0] _19_;
  wire [31:0] _20_;
  wire [31:0] _21_;
  wire [31:0] _22_;
  input [1:0] color_depth_i;
  input [31:0] color_i;
  output [31:0] mem_o;
  output [3:0] sel_o;
  input [1:0] x_lsb_i;
  assign _00_ = ! color_depth_i;
  assign _01_ = ! x_lsb_i;
  assign _02_ = x_lsb_i == 1'b1;
  assign _03_ = x_lsb_i == 2'b10;
  assign _04_ = x_lsb_i == 2'b11;
  assign _05_ = color_depth_i == 1'b1;
  assign _06_ = ~ x_lsb_i[0];
  assign _07_ = _00_ && _01_;
  assign _08_ = _00_ && _02_;
  assign _09_ = _00_ && _03_;
  assign _10_ = _00_ && _04_;
  assign _11_ = _05_ && _06_;
  assign _12_ = _05_ && x_lsb_i[0];
  assign _13_ = _12_ ? 4'b0011 : 4'b1111;
  assign _14_ = _11_ ? 4'b1100 : _13_;
  assign _15_ = _10_ ? 4'b0001 : _14_;
  assign _16_ = _09_ ? 4'b0010 : _15_;
  assign _17_ = _08_ ? 4'b0100 : _16_;
  assign sel_o = _07_ ? 4'b1000 : _17_;
  assign _18_ = _12_ ? { 16'b0000000000000000, color_i[15:0] } : color_i;
  assign _19_ = _11_ ? { color_i[15:0], 16'b0000000000000000 } : _18_;
  assign _20_ = _10_ ? { 24'b000000000000000000000000, color_i[7:0] } : _19_;
  assign _21_ = _09_ ? { 16'b0000000000000000, color_i[7:0], 8'b00000000 } : _20_;
  assign _22_ = _08_ ? { 8'b00000000, color_i[7:0], 16'b0000000000000000 } : _21_;
  assign mem_o = _07_ ? { color_i[7:0], 24'b000000000000000000000000 } : _22_;
endmodule
