module SDP_X_X_trt_core(nvdla_core_clk, nvdla_core_rstn, chn_trt_in_rsc_slz, chn_trt_in_rsc_sz, chn_trt_in_rsc_z, chn_trt_in_rsc_vz, chn_trt_in_rsc_lz, cfg_mul_shift_value_rsc_triosy_lz, cfg_precision, chn_trt_out_rsc_z, chn_trt_out_rsc_vz, chn_trt_out_rsc_lz, chn_trt_in_rsci_oswt, chn_trt_in_rsci_oswt_unreg, cfg_mul_shift_value_rsci_d, chn_trt_out_rsci_oswt, cfg_mul_shift_value_rsc_triosy_obj_oswt, chn_trt_out_rsci_oswt_unreg_pff);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59652" *)
  wire [29:0] _0031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59084" *)
  wire _0032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59094" *)
  wire _0033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59102" *)
  wire _0034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59244" *)
  wire [29:0] _0035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59255" *)
  wire [29:0] _0038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59266" *)
  wire [29:0] _0041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59277" *)
  wire [29:0] _0044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59288" *)
  wire [29:0] _0047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59299" *)
  wire [29:0] _0050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59112" *)
  wire [29:0] _0053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59310" *)
  wire [29:0] _0054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59321" *)
  wire [29:0] _0059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59332" *)
  wire [29:0] _0062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59343" *)
  wire [29:0] _0065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59354" *)
  wire [29:0] _0068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59365" *)
  wire [29:0] _0071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59376" *)
  wire [29:0] _0074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59222" *)
  wire [29:0] _0076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59233" *)
  wire [29:0] _0079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59084" *)
  wire _0082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59387" *)
  wire _0083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59102" *)
  wire _0084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59123" *)
  wire _0115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59112" *)
  wire [29:0] _0116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59222" *)
  wire [29:0] _0117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59233" *)
  wire [29:0] _0118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59244" *)
  wire [29:0] _0119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59255" *)
  wire [29:0] _0120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59266" *)
  wire [29:0] _0121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59277" *)
  wire [29:0] _0122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59288" *)
  wire [29:0] _0123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59299" *)
  wire [29:0] _0124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59310" *)
  wire [29:0] _0125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59321" *)
  wire [29:0] _0126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59332" *)
  wire [29:0] _0127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59343" *)
  wire [29:0] _0128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59354" *)
  wire [29:0] _0129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59365" *)
  wire [29:0] _0130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59376" *)
  wire [29:0] _0131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58998" *)
  wire _0132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59008" *)
  wire _0133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59010" *)
  wire _0134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59013" *)
  wire _0135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59014" *)
  wire _0136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59015" *)
  wire _0137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59017" *)
  wire _0138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59019" *)
  wire _0139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59019" *)
  wire _0140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59020" *)
  wire _0141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59021" *)
  wire _0142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59023" *)
  wire _0143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59023" *)
  wire _0144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59024" *)
  wire _0145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59025" *)
  wire _0146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59027" *)
  wire _0147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59027" *)
  wire _0148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59028" *)
  wire _0149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59029" *)
  wire _0150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59031" *)
  wire _0151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59031" *)
  wire _0152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59032" *)
  wire _0153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59033" *)
  wire _0154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59035" *)
  wire _0155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59036" *)
  wire _0156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59037" *)
  wire _0157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59037" *)
  wire _0158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59039" *)
  wire _0159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59040" *)
  wire _0160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59041" *)
  wire _0161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59041" *)
  wire _0162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59043" *)
  wire _0163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59044" *)
  wire _0164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59045" *)
  wire _0165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59045" *)
  wire _0166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59047" *)
  wire _0167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59048" *)
  wire _0168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59049" *)
  wire _0169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59049" *)
  wire _0170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59051" *)
  wire _0171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59052" *)
  wire _0172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59053" *)
  wire _0173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59053" *)
  wire _0174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59055" *)
  wire _0175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59056" *)
  wire _0176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59057" *)
  wire _0177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59057" *)
  wire _0178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59059" *)
  wire _0179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59060" *)
  wire _0180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59061" *)
  wire _0181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59061" *)
  wire _0182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59063" *)
  wire _0183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59064" *)
  wire _0184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59065" *)
  wire _0185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59065" *)
  wire _0186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59067" *)
  wire _0187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59068" *)
  wire _0188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59069" *)
  wire _0189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59069" *)
  wire _0190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59071" *)
  wire _0191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59072" *)
  wire _0192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59073" *)
  wire _0193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59073" *)
  wire _0194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59075" *)
  wire _0195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59076" *)
  wire _0196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59077" *)
  wire _0197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59077" *)
  wire _0198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59079" *)
  wire _0199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59080" *)
  wire _0200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59081" *)
  wire _0201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59081" *)
  wire _0202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59090" *)
  wire _0203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59098" *)
  wire _0204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59106" *)
  wire _0205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59107" *)
  wire _0206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59116" *)
  wire _0207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *)
  wire _0208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *)
  wire _0209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *)
  wire _0210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *)
  wire _0211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59118" *)
  wire _0212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59227" *)
  wire _0213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59227" *)
  wire _0214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59227" *)
  wire _0215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59228" *)
  wire _0216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59238" *)
  wire _0217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59238" *)
  wire _0218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59238" *)
  wire _0219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59239" *)
  wire _0220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59249" *)
  wire _0221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59249" *)
  wire _0222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59249" *)
  wire _0223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59250" *)
  wire _0224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59260" *)
  wire _0225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59260" *)
  wire _0226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59260" *)
  wire _0227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59261" *)
  wire _0228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59271" *)
  wire _0229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59271" *)
  wire _0230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59271" *)
  wire _0231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59272" *)
  wire _0232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59282" *)
  wire _0233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59282" *)
  wire _0234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59282" *)
  wire _0235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59283" *)
  wire _0236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59293" *)
  wire _0237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59293" *)
  wire _0238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59293" *)
  wire _0239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59294" *)
  wire _0240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59304" *)
  wire _0241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59304" *)
  wire _0242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59304" *)
  wire _0243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59305" *)
  wire _0244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59315" *)
  wire _0245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59315" *)
  wire _0246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59315" *)
  wire _0247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59316" *)
  wire _0248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59326" *)
  wire _0249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59326" *)
  wire _0250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59326" *)
  wire _0251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59327" *)
  wire _0252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59337" *)
  wire _0253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59337" *)
  wire _0254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59337" *)
  wire _0255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59338" *)
  wire _0256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59348" *)
  wire _0257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59348" *)
  wire _0258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59348" *)
  wire _0259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59349" *)
  wire _0260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59359" *)
  wire _0261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59359" *)
  wire _0262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59359" *)
  wire _0263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59360" *)
  wire _0264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59370" *)
  wire _0265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59370" *)
  wire _0266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59370" *)
  wire _0267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59371" *)
  wire _0268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59381" *)
  wire _0269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59381" *)
  wire _0270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59381" *)
  wire _0271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59382" *)
  wire _0272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59391" *)
  wire _0273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58396" *)
  wire _0274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58436" *)
  wire _0275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58476" *)
  wire _0276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58516" *)
  wire _0277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58556" *)
  wire _0278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58596" *)
  wire _0279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58636" *)
  wire _0280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58676" *)
  wire _0281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58716" *)
  wire _0282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58756" *)
  wire _0283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58796" *)
  wire _0284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58836" *)
  wire _0285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58876" *)
  wire _0286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58916" *)
  wire _0287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58956" *)
  wire _0288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58996" *)
  wire _0289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58394" *)
  wire _0290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58434" *)
  wire _0291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58474" *)
  wire _0292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58514" *)
  wire _0293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58554" *)
  wire _0294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58594" *)
  wire _0295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58634" *)
  wire _0296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58674" *)
  wire _0297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58714" *)
  wire _0298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58754" *)
  wire _0299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58794" *)
  wire _0300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58834" *)
  wire _0301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58874" *)
  wire _0302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58914" *)
  wire _0303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58954" *)
  wire _0304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58994" *)
  wire _0305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58389" *)
  wire _0306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58394" *)
  wire _0307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58396" *)
  wire _0308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58429" *)
  wire _0309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58434" *)
  wire _0310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58436" *)
  wire _0311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58469" *)
  wire _0312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58474" *)
  wire _0313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58476" *)
  wire _0314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58509" *)
  wire _0315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58514" *)
  wire _0316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58516" *)
  wire _0317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58549" *)
  wire _0318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58554" *)
  wire _0319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58556" *)
  wire _0320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58589" *)
  wire _0321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58594" *)
  wire _0322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58596" *)
  wire _0323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58629" *)
  wire _0324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58634" *)
  wire _0325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58636" *)
  wire _0326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58669" *)
  wire _0327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58674" *)
  wire _0328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58676" *)
  wire _0329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58709" *)
  wire _0330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58714" *)
  wire _0331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58716" *)
  wire _0332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58749" *)
  wire _0333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58754" *)
  wire _0334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58756" *)
  wire _0335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58789" *)
  wire _0336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58794" *)
  wire _0337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58796" *)
  wire _0338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58829" *)
  wire _0339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58834" *)
  wire _0340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58836" *)
  wire _0341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58869" *)
  wire _0342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58874" *)
  wire _0343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58876" *)
  wire _0344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58909" *)
  wire _0345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58914" *)
  wire _0346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58916" *)
  wire _0347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58949" *)
  wire _0348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58954" *)
  wire _0349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58956" *)
  wire _0350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58989" *)
  wire _0351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58994" *)
  wire _0352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58996" *)
  wire _0353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58997" *)
  wire _0354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59008" *)
  wire _0355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59012" *)
  wire _0356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59090" *)
  wire _0357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59090" *)
  wire _0358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59116" *)
  wire _0359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59226" *)
  wire _0360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59237" *)
  wire _0361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59248" *)
  wire _0362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59259" *)
  wire _0363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59270" *)
  wire _0364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59281" *)
  wire _0365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59292" *)
  wire _0366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59303" *)
  wire _0367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59314" *)
  wire _0368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59325" *)
  wire _0369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59336" *)
  wire _0370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59347" *)
  wire _0371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59358" *)
  wire _0372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59369" *)
  wire _0373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59380" *)
  wire _0374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59392" *)
  wire _0375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59396" *)
  wire _0376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59406" *)
  wire _0377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59411" *)
  wire _0378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59416" *)
  wire _0379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59421" *)
  wire _0380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59426" *)
  wire _0381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59431" *)
  wire _0382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59436" *)
  wire _0383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59441" *)
  wire _0384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59446" *)
  wire _0385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59451" *)
  wire _0386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59456" *)
  wire _0387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59461" *)
  wire _0388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59466" *)
  wire _0389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59471" *)
  wire _0390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59476" *)
  wire _0391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59481" *)
  wire _0392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59486" *)
  wire _0393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59491" *)
  wire _0394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59496" *)
  wire _0395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59501" *)
  wire _0396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59506" *)
  wire _0397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59511" *)
  wire _0398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59516" *)
  wire _0399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59521" *)
  wire _0400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59526" *)
  wire _0401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59531" *)
  wire _0402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59536" *)
  wire _0403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59541" *)
  wire _0404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59546" *)
  wire _0405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59551" *)
  wire _0406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59556" *)
  wire _0407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58356" *)
  wire _0408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58359" *)
  wire _0409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58359" *)
  wire _0410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58360" *)
  wire _0411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58360" *)
  wire _0412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58361" *)
  wire _0413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58361" *)
  wire _0414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58362" *)
  wire _0415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58362" *)
  wire _0416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58363" *)
  wire _0417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58363" *)
  wire _0418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58364" *)
  wire _0419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58364" *)
  wire _0420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58365" *)
  wire _0421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58365" *)
  wire _0422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58366" *)
  wire _0423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58366" *)
  wire _0424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58367" *)
  wire _0425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58367" *)
  wire _0426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58368" *)
  wire _0427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58368" *)
  wire _0428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58369" *)
  wire _0429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58369" *)
  wire _0430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58370" *)
  wire _0431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58370" *)
  wire _0432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58371" *)
  wire _0433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58371" *)
  wire _0434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58372" *)
  wire _0435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58372" *)
  wire _0436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58373" *)
  wire _0437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58373" *)
  wire _0438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58374" *)
  wire _0439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58374" *)
  wire _0440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58375" *)
  wire _0441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58375" *)
  wire _0442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58376" *)
  wire _0443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58376" *)
  wire _0444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58377" *)
  wire _0445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58377" *)
  wire _0446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58378" *)
  wire _0447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58378" *)
  wire _0448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58379" *)
  wire _0449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58379" *)
  wire _0450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58380" *)
  wire _0451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58380" *)
  wire _0452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58381" *)
  wire _0453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58381" *)
  wire _0454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58382" *)
  wire _0455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58382" *)
  wire _0456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58383" *)
  wire _0457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58383" *)
  wire _0458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58384" *)
  wire _0459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58384" *)
  wire _0460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58385" *)
  wire _0461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58385" *)
  wire _0462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58386" *)
  wire _0463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58386" *)
  wire _0464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58387" *)
  wire _0465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58387" *)
  wire _0466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58388" *)
  wire _0467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58388" *)
  wire _0468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58389" *)
  wire _0469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58389" *)
  wire _0470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58394" *)
  wire _0471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58399" *)
  wire _0472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58399" *)
  wire _0473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58400" *)
  wire _0474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58400" *)
  wire _0475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58401" *)
  wire _0476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58401" *)
  wire _0477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58402" *)
  wire _0478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58402" *)
  wire _0479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58403" *)
  wire _0480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58403" *)
  wire _0481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58404" *)
  wire _0482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58404" *)
  wire _0483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58405" *)
  wire _0484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58405" *)
  wire _0485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58406" *)
  wire _0486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58406" *)
  wire _0487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58407" *)
  wire _0488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58407" *)
  wire _0489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58408" *)
  wire _0490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58408" *)
  wire _0491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58409" *)
  wire _0492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58409" *)
  wire _0493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58410" *)
  wire _0494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58410" *)
  wire _0495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58411" *)
  wire _0496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58411" *)
  wire _0497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58412" *)
  wire _0498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58412" *)
  wire _0499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58413" *)
  wire _0500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58413" *)
  wire _0501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58414" *)
  wire _0502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58414" *)
  wire _0503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58415" *)
  wire _0504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58415" *)
  wire _0505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58416" *)
  wire _0506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58416" *)
  wire _0507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58417" *)
  wire _0508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58417" *)
  wire _0509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58418" *)
  wire _0510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58418" *)
  wire _0511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58419" *)
  wire _0512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58419" *)
  wire _0513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58420" *)
  wire _0514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58420" *)
  wire _0515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58421" *)
  wire _0516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58421" *)
  wire _0517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58422" *)
  wire _0518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58422" *)
  wire _0519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58423" *)
  wire _0520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58423" *)
  wire _0521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58424" *)
  wire _0522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58424" *)
  wire _0523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58425" *)
  wire _0524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58425" *)
  wire _0525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58426" *)
  wire _0526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58426" *)
  wire _0527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58427" *)
  wire _0528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58427" *)
  wire _0529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58428" *)
  wire _0530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58428" *)
  wire _0531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58429" *)
  wire _0532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58429" *)
  wire _0533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58434" *)
  wire _0534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58439" *)
  wire _0535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58439" *)
  wire _0536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58440" *)
  wire _0537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58440" *)
  wire _0538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58441" *)
  wire _0539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58441" *)
  wire _0540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58442" *)
  wire _0541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58442" *)
  wire _0542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58443" *)
  wire _0543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58443" *)
  wire _0544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58444" *)
  wire _0545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58444" *)
  wire _0546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58445" *)
  wire _0547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58445" *)
  wire _0548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58446" *)
  wire _0549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58446" *)
  wire _0550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58447" *)
  wire _0551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58447" *)
  wire _0552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58448" *)
  wire _0553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58448" *)
  wire _0554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58449" *)
  wire _0555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58449" *)
  wire _0556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58450" *)
  wire _0557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58450" *)
  wire _0558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58451" *)
  wire _0559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58451" *)
  wire _0560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58452" *)
  wire _0561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58452" *)
  wire _0562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58453" *)
  wire _0563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58453" *)
  wire _0564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58454" *)
  wire _0565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58454" *)
  wire _0566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58455" *)
  wire _0567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58455" *)
  wire _0568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58456" *)
  wire _0569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58456" *)
  wire _0570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58457" *)
  wire _0571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58457" *)
  wire _0572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58458" *)
  wire _0573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58458" *)
  wire _0574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58459" *)
  wire _0575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58459" *)
  wire _0576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58460" *)
  wire _0577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58460" *)
  wire _0578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58461" *)
  wire _0579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58461" *)
  wire _0580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58462" *)
  wire _0581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58462" *)
  wire _0582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58463" *)
  wire _0583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58463" *)
  wire _0584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58464" *)
  wire _0585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58464" *)
  wire _0586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58465" *)
  wire _0587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58465" *)
  wire _0588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58466" *)
  wire _0589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58466" *)
  wire _0590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58467" *)
  wire _0591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58467" *)
  wire _0592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58468" *)
  wire _0593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58468" *)
  wire _0594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58469" *)
  wire _0595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58469" *)
  wire _0596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58474" *)
  wire _0597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58479" *)
  wire _0598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58479" *)
  wire _0599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58480" *)
  wire _0600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58480" *)
  wire _0601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58481" *)
  wire _0602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58481" *)
  wire _0603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58482" *)
  wire _0604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58482" *)
  wire _0605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58483" *)
  wire _0606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58483" *)
  wire _0607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58484" *)
  wire _0608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58484" *)
  wire _0609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58485" *)
  wire _0610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58485" *)
  wire _0611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58486" *)
  wire _0612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58486" *)
  wire _0613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58487" *)
  wire _0614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58487" *)
  wire _0615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58488" *)
  wire _0616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58488" *)
  wire _0617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58489" *)
  wire _0618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58489" *)
  wire _0619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58490" *)
  wire _0620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58490" *)
  wire _0621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58491" *)
  wire _0622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58491" *)
  wire _0623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58492" *)
  wire _0624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58492" *)
  wire _0625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58493" *)
  wire _0626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58493" *)
  wire _0627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58494" *)
  wire _0628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58494" *)
  wire _0629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58495" *)
  wire _0630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58495" *)
  wire _0631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58496" *)
  wire _0632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58496" *)
  wire _0633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58497" *)
  wire _0634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58497" *)
  wire _0635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58498" *)
  wire _0636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58498" *)
  wire _0637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58499" *)
  wire _0638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58499" *)
  wire _0639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58500" *)
  wire _0640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58500" *)
  wire _0641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58501" *)
  wire _0642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58501" *)
  wire _0643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58502" *)
  wire _0644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58502" *)
  wire _0645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58503" *)
  wire _0646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58503" *)
  wire _0647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58504" *)
  wire _0648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58504" *)
  wire _0649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58505" *)
  wire _0650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58505" *)
  wire _0651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58506" *)
  wire _0652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58506" *)
  wire _0653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58507" *)
  wire _0654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58507" *)
  wire _0655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58508" *)
  wire _0656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58508" *)
  wire _0657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58509" *)
  wire _0658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58509" *)
  wire _0659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58514" *)
  wire _0660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58519" *)
  wire _0661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58519" *)
  wire _0662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58520" *)
  wire _0663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58520" *)
  wire _0664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58521" *)
  wire _0665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58521" *)
  wire _0666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58522" *)
  wire _0667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58522" *)
  wire _0668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58523" *)
  wire _0669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58523" *)
  wire _0670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58524" *)
  wire _0671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58524" *)
  wire _0672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58525" *)
  wire _0673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58525" *)
  wire _0674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58526" *)
  wire _0675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58526" *)
  wire _0676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58527" *)
  wire _0677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58527" *)
  wire _0678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58528" *)
  wire _0679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58528" *)
  wire _0680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58529" *)
  wire _0681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58529" *)
  wire _0682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58530" *)
  wire _0683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58530" *)
  wire _0684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58531" *)
  wire _0685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58531" *)
  wire _0686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58532" *)
  wire _0687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58532" *)
  wire _0688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58533" *)
  wire _0689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58533" *)
  wire _0690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58534" *)
  wire _0691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58534" *)
  wire _0692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58535" *)
  wire _0693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58535" *)
  wire _0694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58536" *)
  wire _0695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58536" *)
  wire _0696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58537" *)
  wire _0697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58537" *)
  wire _0698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58538" *)
  wire _0699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58538" *)
  wire _0700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58539" *)
  wire _0701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58539" *)
  wire _0702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58540" *)
  wire _0703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58540" *)
  wire _0704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58541" *)
  wire _0705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58541" *)
  wire _0706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58542" *)
  wire _0707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58542" *)
  wire _0708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58543" *)
  wire _0709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58543" *)
  wire _0710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58544" *)
  wire _0711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58544" *)
  wire _0712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58545" *)
  wire _0713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58545" *)
  wire _0714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58546" *)
  wire _0715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58546" *)
  wire _0716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58547" *)
  wire _0717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58547" *)
  wire _0718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58548" *)
  wire _0719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58548" *)
  wire _0720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58549" *)
  wire _0721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58549" *)
  wire _0722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58554" *)
  wire _0723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58559" *)
  wire _0724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58559" *)
  wire _0725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58560" *)
  wire _0726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58560" *)
  wire _0727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58561" *)
  wire _0728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58561" *)
  wire _0729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58562" *)
  wire _0730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58562" *)
  wire _0731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58563" *)
  wire _0732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58563" *)
  wire _0733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58564" *)
  wire _0734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58564" *)
  wire _0735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58565" *)
  wire _0736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58565" *)
  wire _0737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58566" *)
  wire _0738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58566" *)
  wire _0739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58567" *)
  wire _0740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58567" *)
  wire _0741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58568" *)
  wire _0742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58568" *)
  wire _0743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58569" *)
  wire _0744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58569" *)
  wire _0745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58570" *)
  wire _0746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58570" *)
  wire _0747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58571" *)
  wire _0748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58571" *)
  wire _0749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58572" *)
  wire _0750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58572" *)
  wire _0751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58573" *)
  wire _0752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58573" *)
  wire _0753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58574" *)
  wire _0754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58574" *)
  wire _0755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58575" *)
  wire _0756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58575" *)
  wire _0757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58576" *)
  wire _0758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58576" *)
  wire _0759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58577" *)
  wire _0760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58577" *)
  wire _0761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58578" *)
  wire _0762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58578" *)
  wire _0763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58579" *)
  wire _0764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58579" *)
  wire _0765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58580" *)
  wire _0766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58580" *)
  wire _0767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58581" *)
  wire _0768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58581" *)
  wire _0769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58582" *)
  wire _0770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58582" *)
  wire _0771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58583" *)
  wire _0772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58583" *)
  wire _0773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58584" *)
  wire _0774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58584" *)
  wire _0775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58585" *)
  wire _0776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58585" *)
  wire _0777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58586" *)
  wire _0778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58586" *)
  wire _0779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58587" *)
  wire _0780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58587" *)
  wire _0781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58588" *)
  wire _0782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58588" *)
  wire _0783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58589" *)
  wire _0784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58589" *)
  wire _0785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58594" *)
  wire _0786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58599" *)
  wire _0787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58599" *)
  wire _0788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58600" *)
  wire _0789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58600" *)
  wire _0790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58601" *)
  wire _0791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58601" *)
  wire _0792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58602" *)
  wire _0793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58602" *)
  wire _0794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58603" *)
  wire _0795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58603" *)
  wire _0796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58604" *)
  wire _0797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58604" *)
  wire _0798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58605" *)
  wire _0799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58605" *)
  wire _0800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58606" *)
  wire _0801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58606" *)
  wire _0802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58607" *)
  wire _0803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58607" *)
  wire _0804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58608" *)
  wire _0805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58608" *)
  wire _0806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58609" *)
  wire _0807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58609" *)
  wire _0808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58610" *)
  wire _0809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58610" *)
  wire _0810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58611" *)
  wire _0811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58611" *)
  wire _0812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58612" *)
  wire _0813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58612" *)
  wire _0814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58613" *)
  wire _0815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58613" *)
  wire _0816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58614" *)
  wire _0817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58614" *)
  wire _0818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58615" *)
  wire _0819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58615" *)
  wire _0820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58616" *)
  wire _0821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58616" *)
  wire _0822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58617" *)
  wire _0823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58617" *)
  wire _0824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58618" *)
  wire _0825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58618" *)
  wire _0826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58619" *)
  wire _0827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58619" *)
  wire _0828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58620" *)
  wire _0829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58620" *)
  wire _0830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58621" *)
  wire _0831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58621" *)
  wire _0832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58622" *)
  wire _0833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58622" *)
  wire _0834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58623" *)
  wire _0835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58623" *)
  wire _0836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58624" *)
  wire _0837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58624" *)
  wire _0838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58625" *)
  wire _0839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58625" *)
  wire _0840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58626" *)
  wire _0841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58626" *)
  wire _0842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58627" *)
  wire _0843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58627" *)
  wire _0844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58628" *)
  wire _0845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58628" *)
  wire _0846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58629" *)
  wire _0847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58629" *)
  wire _0848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58634" *)
  wire _0849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58639" *)
  wire _0850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58639" *)
  wire _0851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58640" *)
  wire _0852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58640" *)
  wire _0853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58641" *)
  wire _0854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58641" *)
  wire _0855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58642" *)
  wire _0856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58642" *)
  wire _0857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58643" *)
  wire _0858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58643" *)
  wire _0859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58644" *)
  wire _0860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58644" *)
  wire _0861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58645" *)
  wire _0862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58645" *)
  wire _0863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58646" *)
  wire _0864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58646" *)
  wire _0865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58647" *)
  wire _0866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58647" *)
  wire _0867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58648" *)
  wire _0868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58648" *)
  wire _0869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58649" *)
  wire _0870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58649" *)
  wire _0871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58650" *)
  wire _0872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58650" *)
  wire _0873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58651" *)
  wire _0874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58651" *)
  wire _0875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58652" *)
  wire _0876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58652" *)
  wire _0877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58653" *)
  wire _0878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58653" *)
  wire _0879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58654" *)
  wire _0880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58654" *)
  wire _0881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58655" *)
  wire _0882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58655" *)
  wire _0883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58656" *)
  wire _0884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58656" *)
  wire _0885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58657" *)
  wire _0886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58657" *)
  wire _0887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58658" *)
  wire _0888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58658" *)
  wire _0889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58659" *)
  wire _0890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58659" *)
  wire _0891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58660" *)
  wire _0892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58660" *)
  wire _0893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58661" *)
  wire _0894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58661" *)
  wire _0895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58662" *)
  wire _0896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58662" *)
  wire _0897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58663" *)
  wire _0898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58663" *)
  wire _0899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58664" *)
  wire _0900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58664" *)
  wire _0901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58665" *)
  wire _0902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58665" *)
  wire _0903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58666" *)
  wire _0904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58666" *)
  wire _0905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58667" *)
  wire _0906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58667" *)
  wire _0907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58668" *)
  wire _0908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58668" *)
  wire _0909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58669" *)
  wire _0910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58669" *)
  wire _0911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58674" *)
  wire _0912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58679" *)
  wire _0913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58679" *)
  wire _0914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58680" *)
  wire _0915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58680" *)
  wire _0916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58681" *)
  wire _0917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58681" *)
  wire _0918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58682" *)
  wire _0919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58682" *)
  wire _0920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58683" *)
  wire _0921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58683" *)
  wire _0922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58684" *)
  wire _0923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58684" *)
  wire _0924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58685" *)
  wire _0925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58685" *)
  wire _0926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58686" *)
  wire _0927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58686" *)
  wire _0928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58687" *)
  wire _0929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58687" *)
  wire _0930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58688" *)
  wire _0931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58688" *)
  wire _0932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58689" *)
  wire _0933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58689" *)
  wire _0934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58690" *)
  wire _0935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58690" *)
  wire _0936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58691" *)
  wire _0937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58691" *)
  wire _0938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58692" *)
  wire _0939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58692" *)
  wire _0940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58693" *)
  wire _0941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58693" *)
  wire _0942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58694" *)
  wire _0943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58694" *)
  wire _0944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58695" *)
  wire _0945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58695" *)
  wire _0946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58696" *)
  wire _0947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58696" *)
  wire _0948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58697" *)
  wire _0949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58697" *)
  wire _0950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58698" *)
  wire _0951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58698" *)
  wire _0952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58699" *)
  wire _0953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58699" *)
  wire _0954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58700" *)
  wire _0955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58700" *)
  wire _0956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58701" *)
  wire _0957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58701" *)
  wire _0958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58702" *)
  wire _0959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58702" *)
  wire _0960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58703" *)
  wire _0961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58703" *)
  wire _0962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58704" *)
  wire _0963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58704" *)
  wire _0964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58705" *)
  wire _0965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58705" *)
  wire _0966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58706" *)
  wire _0967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58706" *)
  wire _0968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58707" *)
  wire _0969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58707" *)
  wire _0970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58708" *)
  wire _0971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58708" *)
  wire _0972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58709" *)
  wire _0973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58709" *)
  wire _0974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58714" *)
  wire _0975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58719" *)
  wire _0976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58719" *)
  wire _0977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58720" *)
  wire _0978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58720" *)
  wire _0979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58721" *)
  wire _0980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58721" *)
  wire _0981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58722" *)
  wire _0982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58722" *)
  wire _0983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58723" *)
  wire _0984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58723" *)
  wire _0985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58724" *)
  wire _0986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58724" *)
  wire _0987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58725" *)
  wire _0988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58725" *)
  wire _0989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58726" *)
  wire _0990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58726" *)
  wire _0991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58727" *)
  wire _0992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58727" *)
  wire _0993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58728" *)
  wire _0994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58728" *)
  wire _0995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58729" *)
  wire _0996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58729" *)
  wire _0997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58730" *)
  wire _0998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58730" *)
  wire _0999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58731" *)
  wire _1000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58731" *)
  wire _1001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58732" *)
  wire _1002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58732" *)
  wire _1003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58733" *)
  wire _1004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58733" *)
  wire _1005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58734" *)
  wire _1006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58734" *)
  wire _1007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58735" *)
  wire _1008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58735" *)
  wire _1009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58736" *)
  wire _1010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58736" *)
  wire _1011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58737" *)
  wire _1012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58737" *)
  wire _1013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58738" *)
  wire _1014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58738" *)
  wire _1015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58739" *)
  wire _1016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58739" *)
  wire _1017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58740" *)
  wire _1018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58740" *)
  wire _1019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58741" *)
  wire _1020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58741" *)
  wire _1021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58742" *)
  wire _1022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58742" *)
  wire _1023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58743" *)
  wire _1024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58743" *)
  wire _1025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58744" *)
  wire _1026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58744" *)
  wire _1027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58745" *)
  wire _1028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58745" *)
  wire _1029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58746" *)
  wire _1030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58746" *)
  wire _1031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58747" *)
  wire _1032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58747" *)
  wire _1033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58748" *)
  wire _1034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58748" *)
  wire _1035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58749" *)
  wire _1036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58749" *)
  wire _1037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58754" *)
  wire _1038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58759" *)
  wire _1039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58759" *)
  wire _1040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58760" *)
  wire _1041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58760" *)
  wire _1042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58761" *)
  wire _1043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58761" *)
  wire _1044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58762" *)
  wire _1045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58762" *)
  wire _1046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58763" *)
  wire _1047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58763" *)
  wire _1048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58764" *)
  wire _1049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58764" *)
  wire _1050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58765" *)
  wire _1051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58765" *)
  wire _1052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58766" *)
  wire _1053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58766" *)
  wire _1054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58767" *)
  wire _1055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58767" *)
  wire _1056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58768" *)
  wire _1057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58768" *)
  wire _1058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58769" *)
  wire _1059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58769" *)
  wire _1060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58770" *)
  wire _1061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58770" *)
  wire _1062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58771" *)
  wire _1063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58771" *)
  wire _1064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58772" *)
  wire _1065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58772" *)
  wire _1066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58773" *)
  wire _1067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58773" *)
  wire _1068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58774" *)
  wire _1069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58774" *)
  wire _1070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58775" *)
  wire _1071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58775" *)
  wire _1072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58776" *)
  wire _1073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58776" *)
  wire _1074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58777" *)
  wire _1075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58777" *)
  wire _1076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58778" *)
  wire _1077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58778" *)
  wire _1078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58779" *)
  wire _1079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58779" *)
  wire _1080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58780" *)
  wire _1081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58780" *)
  wire _1082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58781" *)
  wire _1083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58781" *)
  wire _1084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58782" *)
  wire _1085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58782" *)
  wire _1086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58783" *)
  wire _1087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58783" *)
  wire _1088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58784" *)
  wire _1089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58784" *)
  wire _1090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58785" *)
  wire _1091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58785" *)
  wire _1092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58786" *)
  wire _1093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58786" *)
  wire _1094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58787" *)
  wire _1095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58787" *)
  wire _1096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58788" *)
  wire _1097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58788" *)
  wire _1098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58789" *)
  wire _1099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58789" *)
  wire _1100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58794" *)
  wire _1101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58799" *)
  wire _1102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58799" *)
  wire _1103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58800" *)
  wire _1104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58800" *)
  wire _1105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58801" *)
  wire _1106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58801" *)
  wire _1107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58802" *)
  wire _1108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58802" *)
  wire _1109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58803" *)
  wire _1110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58803" *)
  wire _1111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58804" *)
  wire _1112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58804" *)
  wire _1113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58805" *)
  wire _1114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58805" *)
  wire _1115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58806" *)
  wire _1116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58806" *)
  wire _1117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58807" *)
  wire _1118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58807" *)
  wire _1119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58808" *)
  wire _1120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58808" *)
  wire _1121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58809" *)
  wire _1122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58809" *)
  wire _1123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58810" *)
  wire _1124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58810" *)
  wire _1125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58811" *)
  wire _1126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58811" *)
  wire _1127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58812" *)
  wire _1128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58812" *)
  wire _1129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58813" *)
  wire _1130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58813" *)
  wire _1131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58814" *)
  wire _1132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58814" *)
  wire _1133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58815" *)
  wire _1134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58815" *)
  wire _1135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58816" *)
  wire _1136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58816" *)
  wire _1137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58817" *)
  wire _1138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58817" *)
  wire _1139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58818" *)
  wire _1140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58818" *)
  wire _1141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58819" *)
  wire _1142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58819" *)
  wire _1143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58820" *)
  wire _1144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58820" *)
  wire _1145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58821" *)
  wire _1146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58821" *)
  wire _1147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58822" *)
  wire _1148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58822" *)
  wire _1149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58823" *)
  wire _1150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58823" *)
  wire _1151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58824" *)
  wire _1152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58824" *)
  wire _1153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58825" *)
  wire _1154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58825" *)
  wire _1155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58826" *)
  wire _1156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58826" *)
  wire _1157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58827" *)
  wire _1158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58827" *)
  wire _1159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58828" *)
  wire _1160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58828" *)
  wire _1161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58829" *)
  wire _1162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58829" *)
  wire _1163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58834" *)
  wire _1164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58839" *)
  wire _1165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58839" *)
  wire _1166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58840" *)
  wire _1167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58840" *)
  wire _1168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58841" *)
  wire _1169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58841" *)
  wire _1170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58842" *)
  wire _1171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58842" *)
  wire _1172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58843" *)
  wire _1173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58843" *)
  wire _1174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58844" *)
  wire _1175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58844" *)
  wire _1176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58845" *)
  wire _1177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58845" *)
  wire _1178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58846" *)
  wire _1179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58846" *)
  wire _1180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58847" *)
  wire _1181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58847" *)
  wire _1182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58848" *)
  wire _1183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58848" *)
  wire _1184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58849" *)
  wire _1185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58849" *)
  wire _1186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58850" *)
  wire _1187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58850" *)
  wire _1188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58851" *)
  wire _1189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58851" *)
  wire _1190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58852" *)
  wire _1191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58852" *)
  wire _1192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58853" *)
  wire _1193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58853" *)
  wire _1194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58854" *)
  wire _1195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58854" *)
  wire _1196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58855" *)
  wire _1197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58855" *)
  wire _1198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58856" *)
  wire _1199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58856" *)
  wire _1200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58857" *)
  wire _1201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58857" *)
  wire _1202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58858" *)
  wire _1203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58858" *)
  wire _1204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58859" *)
  wire _1205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58859" *)
  wire _1206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58860" *)
  wire _1207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58860" *)
  wire _1208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58861" *)
  wire _1209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58861" *)
  wire _1210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58862" *)
  wire _1211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58862" *)
  wire _1212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58863" *)
  wire _1213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58863" *)
  wire _1214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58864" *)
  wire _1215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58864" *)
  wire _1216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58865" *)
  wire _1217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58865" *)
  wire _1218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58866" *)
  wire _1219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58866" *)
  wire _1220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58867" *)
  wire _1221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58867" *)
  wire _1222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58868" *)
  wire _1223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58868" *)
  wire _1224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58869" *)
  wire _1225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58869" *)
  wire _1226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58874" *)
  wire _1227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58879" *)
  wire _1228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58879" *)
  wire _1229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58880" *)
  wire _1230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58880" *)
  wire _1231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58881" *)
  wire _1232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58881" *)
  wire _1233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58882" *)
  wire _1234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58882" *)
  wire _1235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58883" *)
  wire _1236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58883" *)
  wire _1237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58884" *)
  wire _1238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58884" *)
  wire _1239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58885" *)
  wire _1240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58885" *)
  wire _1241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58886" *)
  wire _1242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58886" *)
  wire _1243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58887" *)
  wire _1244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58887" *)
  wire _1245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58888" *)
  wire _1246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58888" *)
  wire _1247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58889" *)
  wire _1248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58889" *)
  wire _1249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58890" *)
  wire _1250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58890" *)
  wire _1251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58891" *)
  wire _1252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58891" *)
  wire _1253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58892" *)
  wire _1254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58892" *)
  wire _1255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58893" *)
  wire _1256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58893" *)
  wire _1257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58894" *)
  wire _1258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58894" *)
  wire _1259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58895" *)
  wire _1260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58895" *)
  wire _1261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58896" *)
  wire _1262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58896" *)
  wire _1263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58897" *)
  wire _1264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58897" *)
  wire _1265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58898" *)
  wire _1266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58898" *)
  wire _1267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58899" *)
  wire _1268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58899" *)
  wire _1269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58900" *)
  wire _1270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58900" *)
  wire _1271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58901" *)
  wire _1272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58901" *)
  wire _1273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58902" *)
  wire _1274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58902" *)
  wire _1275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58903" *)
  wire _1276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58903" *)
  wire _1277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58904" *)
  wire _1278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58904" *)
  wire _1279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58905" *)
  wire _1280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58905" *)
  wire _1281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58906" *)
  wire _1282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58906" *)
  wire _1283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58907" *)
  wire _1284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58907" *)
  wire _1285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58908" *)
  wire _1286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58908" *)
  wire _1287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58909" *)
  wire _1288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58909" *)
  wire _1289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58914" *)
  wire _1290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58919" *)
  wire _1291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58919" *)
  wire _1292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58920" *)
  wire _1293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58920" *)
  wire _1294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58921" *)
  wire _1295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58921" *)
  wire _1296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58922" *)
  wire _1297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58922" *)
  wire _1298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58923" *)
  wire _1299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58923" *)
  wire _1300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58924" *)
  wire _1301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58924" *)
  wire _1302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58925" *)
  wire _1303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58925" *)
  wire _1304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58926" *)
  wire _1305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58926" *)
  wire _1306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58927" *)
  wire _1307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58927" *)
  wire _1308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58928" *)
  wire _1309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58928" *)
  wire _1310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58929" *)
  wire _1311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58929" *)
  wire _1312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58930" *)
  wire _1313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58930" *)
  wire _1314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58931" *)
  wire _1315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58931" *)
  wire _1316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58932" *)
  wire _1317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58932" *)
  wire _1318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58933" *)
  wire _1319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58933" *)
  wire _1320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58934" *)
  wire _1321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58934" *)
  wire _1322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58935" *)
  wire _1323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58935" *)
  wire _1324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58936" *)
  wire _1325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58936" *)
  wire _1326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58937" *)
  wire _1327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58937" *)
  wire _1328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58938" *)
  wire _1329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58938" *)
  wire _1330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58939" *)
  wire _1331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58939" *)
  wire _1332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58940" *)
  wire _1333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58940" *)
  wire _1334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58941" *)
  wire _1335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58941" *)
  wire _1336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58942" *)
  wire _1337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58942" *)
  wire _1338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58943" *)
  wire _1339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58943" *)
  wire _1340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58944" *)
  wire _1341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58944" *)
  wire _1342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58945" *)
  wire _1343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58945" *)
  wire _1344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58946" *)
  wire _1345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58946" *)
  wire _1346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58947" *)
  wire _1347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58947" *)
  wire _1348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58948" *)
  wire _1349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58948" *)
  wire _1350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58949" *)
  wire _1351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58949" *)
  wire _1352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58954" *)
  wire _1353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58959" *)
  wire _1354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58959" *)
  wire _1355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58960" *)
  wire _1356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58960" *)
  wire _1357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58961" *)
  wire _1358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58961" *)
  wire _1359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58962" *)
  wire _1360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58962" *)
  wire _1361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58963" *)
  wire _1362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58963" *)
  wire _1363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58964" *)
  wire _1364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58964" *)
  wire _1365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58965" *)
  wire _1366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58965" *)
  wire _1367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58966" *)
  wire _1368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58966" *)
  wire _1369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58967" *)
  wire _1370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58967" *)
  wire _1371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58968" *)
  wire _1372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58968" *)
  wire _1373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58969" *)
  wire _1374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58969" *)
  wire _1375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58970" *)
  wire _1376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58970" *)
  wire _1377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58971" *)
  wire _1378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58971" *)
  wire _1379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58972" *)
  wire _1380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58972" *)
  wire _1381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58973" *)
  wire _1382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58973" *)
  wire _1383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58974" *)
  wire _1384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58974" *)
  wire _1385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58975" *)
  wire _1386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58975" *)
  wire _1387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58976" *)
  wire _1388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58976" *)
  wire _1389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58977" *)
  wire _1390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58977" *)
  wire _1391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58978" *)
  wire _1392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58978" *)
  wire _1393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58979" *)
  wire _1394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58979" *)
  wire _1395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58980" *)
  wire _1396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58980" *)
  wire _1397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58981" *)
  wire _1398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58981" *)
  wire _1399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58982" *)
  wire _1400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58982" *)
  wire _1401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58983" *)
  wire _1402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58983" *)
  wire _1403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58984" *)
  wire _1404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58984" *)
  wire _1405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58985" *)
  wire _1406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58985" *)
  wire _1407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58986" *)
  wire _1408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58986" *)
  wire _1409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58987" *)
  wire _1410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58987" *)
  wire _1411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58988" *)
  wire _1412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58988" *)
  wire _1413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58989" *)
  wire _1414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58989" *)
  wire _1415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58994" *)
  wire _1416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58997" *)
  wire _1417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58998" *)
  wire _1418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59008" *)
  wire _1419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59020" *)
  wire _1420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59024" *)
  wire _1421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59028" *)
  wire _1422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59032" *)
  wire _1423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59036" *)
  wire _1424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59040" *)
  wire _1425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59044" *)
  wire _1426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59048" *)
  wire _1427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59052" *)
  wire _1428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59056" *)
  wire _1429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59060" *)
  wire _1430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59064" *)
  wire _1431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59068" *)
  wire _1432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59072" *)
  wire _1433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59076" *)
  wire _1434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59080" *)
  wire _1435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59106" *)
  wire _1436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59106" *)
  wire _1437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59118" *)
  wire _1438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59118" *)
  wire _1439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59228" *)
  wire _1440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59228" *)
  wire _1441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59239" *)
  wire _1442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59239" *)
  wire _1443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59250" *)
  wire _1444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59250" *)
  wire _1445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59261" *)
  wire _1446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59261" *)
  wire _1447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59272" *)
  wire _1448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59272" *)
  wire _1449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59283" *)
  wire _1450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59283" *)
  wire _1451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59294" *)
  wire _1452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59294" *)
  wire _1453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59305" *)
  wire _1454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59305" *)
  wire _1455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59316" *)
  wire _1456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59316" *)
  wire _1457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59327" *)
  wire _1458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59327" *)
  wire _1459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59338" *)
  wire _1460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59338" *)
  wire _1461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59349" *)
  wire _1462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59349" *)
  wire _1463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59360" *)
  wire _1464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59360" *)
  wire _1465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59371" *)
  wire _1466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59371" *)
  wire _1467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59382" *)
  wire _1468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59382" *)
  wire _1469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59391" *)
  wire _1470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59396" *)
  wire _1471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59397" *)
  wire _1472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59406" *)
  wire _1473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59407" *)
  wire _1474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59411" *)
  wire _1475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59412" *)
  wire _1476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59416" *)
  wire _1477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59417" *)
  wire _1478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59421" *)
  wire _1479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59422" *)
  wire _1480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59426" *)
  wire _1481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59427" *)
  wire _1482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59431" *)
  wire _1483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59432" *)
  wire _1484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59436" *)
  wire _1485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59437" *)
  wire _1486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59441" *)
  wire _1487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59442" *)
  wire _1488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59446" *)
  wire _1489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59447" *)
  wire _1490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59451" *)
  wire _1491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59452" *)
  wire _1492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59456" *)
  wire _1493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59457" *)
  wire _1494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59461" *)
  wire _1495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59462" *)
  wire _1496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59466" *)
  wire _1497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59467" *)
  wire _1498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59471" *)
  wire _1499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59472" *)
  wire _1500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59476" *)
  wire _1501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59477" *)
  wire _1502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59481" *)
  wire _1503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59482" *)
  wire _1504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59486" *)
  wire _1505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59487" *)
  wire _1506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59491" *)
  wire _1507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59492" *)
  wire _1508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59496" *)
  wire _1509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59497" *)
  wire _1510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59501" *)
  wire _1511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59502" *)
  wire _1512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59506" *)
  wire _1513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59507" *)
  wire _1514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59511" *)
  wire _1515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59512" *)
  wire _1516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59516" *)
  wire _1517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59517" *)
  wire _1518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59521" *)
  wire _1519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59522" *)
  wire _1520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59526" *)
  wire _1521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59527" *)
  wire _1522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59531" *)
  wire _1523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59532" *)
  wire _1524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59536" *)
  wire _1525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59537" *)
  wire _1526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59541" *)
  wire _1527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59542" *)
  wire _1528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59546" *)
  wire _1529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59547" *)
  wire _1530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59551" *)
  wire _1531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59552" *)
  wire _1532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59556" *)
  wire _1533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59557" *)
  wire _1534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57874" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57873" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57872" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57871" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57870" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57869" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57883" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57882" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57881" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57880" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57879" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57878" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57877" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57876" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57875" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57868" *)
  wire [111:0] IntShiftRight_49U_6U_32U_mbits_fixed_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57896" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57894" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57892" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57890" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57888" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57886" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57914" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57912" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57910" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57908" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57906" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57904" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57902" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57900" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57898" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57884" *)
  wire [49:0] IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57956" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57958" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57960" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57962" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57964" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57966" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57938" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57940" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57942" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57944" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57946" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57948" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57950" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57952" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57954" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57968" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57955" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57957" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57959" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57961" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57963" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57965" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57937" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57939" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57941" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57943" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57945" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57947" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57949" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57951" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57953" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57967" *)
  wire IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57865" *)
  wire and_148_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57866" *)
  wire and_150_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57867" *)
  wire and_4_mdf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57851" *)
  wire and_dcpl_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57856" *)
  wire and_dcpl_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57863" *)
  wire and_dcpl_134;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57857" *)
  wire and_dcpl_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57858" *)
  wire and_dcpl_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57859" *)
  wire and_dcpl_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57861" *)
  wire and_dcpl_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57862" *)
  wire and_dcpl_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57853" *)
  wire and_dcpl_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57855" *)
  wire and_dcpl_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57780" *)
  output cfg_mul_shift_value_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57801" *)
  wire cfg_mul_shift_value_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57789" *)
  input cfg_mul_shift_value_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57787" *)
  input [5:0] cfg_mul_shift_value_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57781" *)
  input [1:0] cfg_precision;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57779" *)
  output chn_trt_in_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57775" *)
  output chn_trt_in_rsc_slz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57776" *)
  input chn_trt_in_rsc_sz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57778" *)
  input chn_trt_in_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57777" *)
  input [799:0] chn_trt_in_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57794" *)
  wire chn_trt_in_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57797" *)
  wire [799:0] chn_trt_in_rsci_d_mxwt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57793" *)
  reg chn_trt_in_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57796" *)
  reg chn_trt_in_rsci_ld_core_psct;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57919" *)
  wire chn_trt_in_rsci_ld_core_psct_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57785" *)
  input chn_trt_in_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57786" *)
  output chn_trt_in_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57795" *)
  wire chn_trt_in_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57916" *)
  wire chn_trt_out_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57784" *)
  output chn_trt_out_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57783" *)
  input chn_trt_out_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57782" *)
  output [511:0] chn_trt_out_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57799" *)
  wire chn_trt_out_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57849" *)
  reg chn_trt_out_rsci_d_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57920" *)
  wire chn_trt_out_rsci_d_0_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57839" *)
  reg [29:0] chn_trt_out_rsci_d_126_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57924" *)
  wire chn_trt_out_rsci_d_126_97_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57838" *)
  reg chn_trt_out_rsci_d_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57837" *)
  reg chn_trt_out_rsci_d_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57836" *)
  reg [29:0] chn_trt_out_rsci_d_158_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57925" *)
  wire chn_trt_out_rsci_d_158_129_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57835" *)
  reg chn_trt_out_rsci_d_159;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57834" *)
  reg chn_trt_out_rsci_d_160;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57833" *)
  reg [29:0] chn_trt_out_rsci_d_190_161;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57926" *)
  wire chn_trt_out_rsci_d_190_161_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57832" *)
  reg chn_trt_out_rsci_d_191;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57831" *)
  reg chn_trt_out_rsci_d_192;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57830" *)
  reg [29:0] chn_trt_out_rsci_d_222_193;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57927" *)
  wire chn_trt_out_rsci_d_222_193_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57829" *)
  reg chn_trt_out_rsci_d_223;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57828" *)
  reg chn_trt_out_rsci_d_224;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57827" *)
  reg [29:0] chn_trt_out_rsci_d_254_225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57928" *)
  wire chn_trt_out_rsci_d_254_225_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57826" *)
  reg chn_trt_out_rsci_d_255;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57825" *)
  reg chn_trt_out_rsci_d_256;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57824" *)
  reg [29:0] chn_trt_out_rsci_d_286_257;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57929" *)
  wire chn_trt_out_rsci_d_286_257_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57823" *)
  reg chn_trt_out_rsci_d_287;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57822" *)
  reg chn_trt_out_rsci_d_288;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57848" *)
  reg [29:0] chn_trt_out_rsci_d_30_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57921" *)
  wire chn_trt_out_rsci_d_30_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57847" *)
  reg chn_trt_out_rsci_d_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57821" *)
  reg [29:0] chn_trt_out_rsci_d_318_289;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57930" *)
  wire chn_trt_out_rsci_d_318_289_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57820" *)
  reg chn_trt_out_rsci_d_319;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57846" *)
  reg chn_trt_out_rsci_d_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57819" *)
  reg chn_trt_out_rsci_d_320;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57818" *)
  reg [29:0] chn_trt_out_rsci_d_350_321;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57931" *)
  wire chn_trt_out_rsci_d_350_321_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57817" *)
  reg chn_trt_out_rsci_d_351;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57816" *)
  reg chn_trt_out_rsci_d_352;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57815" *)
  reg [29:0] chn_trt_out_rsci_d_382_353;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57932" *)
  wire chn_trt_out_rsci_d_382_353_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57814" *)
  reg chn_trt_out_rsci_d_383;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57813" *)
  reg chn_trt_out_rsci_d_384;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57812" *)
  reg [29:0] chn_trt_out_rsci_d_414_385;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57933" *)
  wire chn_trt_out_rsci_d_414_385_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57811" *)
  reg chn_trt_out_rsci_d_415;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57810" *)
  reg chn_trt_out_rsci_d_416;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57809" *)
  reg [29:0] chn_trt_out_rsci_d_446_417;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57934" *)
  wire chn_trt_out_rsci_d_446_417_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57808" *)
  reg chn_trt_out_rsci_d_447;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57807" *)
  reg chn_trt_out_rsci_d_448;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57806" *)
  reg [29:0] chn_trt_out_rsci_d_478_449;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57935" *)
  wire chn_trt_out_rsci_d_478_449_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57805" *)
  reg chn_trt_out_rsci_d_479;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57804" *)
  reg chn_trt_out_rsci_d_480;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57803" *)
  reg [29:0] chn_trt_out_rsci_d_510_481;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57936" *)
  wire chn_trt_out_rsci_d_510_481_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57802" *)
  reg chn_trt_out_rsci_d_511;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57845" *)
  reg [29:0] chn_trt_out_rsci_d_62_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57922" *)
  wire chn_trt_out_rsci_d_62_33_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57844" *)
  reg chn_trt_out_rsci_d_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57843" *)
  reg chn_trt_out_rsci_d_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57842" *)
  reg [29:0] chn_trt_out_rsci_d_94_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57923" *)
  wire chn_trt_out_rsci_d_94_65_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57841" *)
  reg chn_trt_out_rsci_d_95;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57840" *)
  reg chn_trt_out_rsci_d_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57788" *)
  input chn_trt_out_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57790" *)
  output chn_trt_out_rsci_oswt_unreg_pff;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57800" *)
  wire chn_trt_out_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57792" *)
  wire core_wen;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57798" *)
  wire core_wten;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57850" *)
  wire [1:0] fsm_output;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58087" *)
  wire mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58088" *)
  wire mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58089" *)
  wire mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58090" *)
  wire mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58091" *)
  wire mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58092" *)
  wire mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58093" *)
  wire mux_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58094" *)
  wire mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58095" *)
  wire mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58096" *)
  wire mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58081" *)
  wire mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58082" *)
  wire mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58083" *)
  wire mux_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58084" *)
  wire mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58085" *)
  wire mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58086" *)
  wire mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57897" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57895" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57893" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57891" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57889" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57887" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57915" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57913" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57911" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57909" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57907" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57905" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57903" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57901" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57899" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57885" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58146" *)
  wire [511:0] nl_X_trt_core_chn_trt_out_rsci_inst_chn_trt_out_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58125" *)
  wire [111:0] nl_trt_loop_10_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58128" *)
  wire [111:0] nl_trt_loop_11_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58131" *)
  wire [111:0] nl_trt_loop_12_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58134" *)
  wire [111:0] nl_trt_loop_13_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58137" *)
  wire [111:0] nl_trt_loop_14_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58140" *)
  wire [111:0] nl_trt_loop_15_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58143" *)
  wire [111:0] nl_trt_loop_16_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58098" *)
  wire [111:0] nl_trt_loop_1_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58101" *)
  wire [111:0] nl_trt_loop_2_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58104" *)
  wire [111:0] nl_trt_loop_3_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58107" *)
  wire [111:0] nl_trt_loop_4_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58110" *)
  wire [111:0] nl_trt_loop_5_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58113" *)
  wire [111:0] nl_trt_loop_6_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58116" *)
  wire [111:0] nl_trt_loop_7_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58119" *)
  wire [111:0] nl_trt_loop_8_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58122" *)
  wire [111:0] nl_trt_loop_9_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57860" *)
  wire not_tmp_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57773" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57774" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57852" *)
  wire or_dcpl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57854" *)
  wire or_dcpl_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57864" *)
  wire or_tmp_150;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57917" *)
  reg reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57918" *)
  reg reg_chn_trt_out_rsci_ld_core_psct_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58024" *)
  wire trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58028" *)
  wire trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58025" *)
  wire [29:0] trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58074" *)
  wire trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58026" *)
  wire [29:0] trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58030" *)
  wire trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58034" *)
  wire trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58031" *)
  wire [29:0] trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58075" *)
  wire trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58032" *)
  wire [29:0] trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58036" *)
  wire trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58040" *)
  wire trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58037" *)
  wire [29:0] trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58076" *)
  wire trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58038" *)
  wire [29:0] trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58042" *)
  wire trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58046" *)
  wire trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58043" *)
  wire [29:0] trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58077" *)
  wire trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58044" *)
  wire [29:0] trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58048" *)
  wire trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58052" *)
  wire trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58049" *)
  wire [29:0] trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58078" *)
  wire trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58050" *)
  wire [29:0] trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58054" *)
  wire trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58058" *)
  wire trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58055" *)
  wire [29:0] trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58079" *)
  wire trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58056" *)
  wire [29:0] trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58060" *)
  wire trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58064" *)
  wire trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58061" *)
  wire [29:0] trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58080" *)
  wire trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58062" *)
  wire [29:0] trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57970" *)
  wire trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57974" *)
  wire trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57971" *)
  wire [29:0] trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58065" *)
  wire trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57972" *)
  wire [29:0] trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57976" *)
  wire trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57980" *)
  wire trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57977" *)
  wire [29:0] trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58066" *)
  wire trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57978" *)
  wire [29:0] trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57982" *)
  wire trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57986" *)
  wire trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57983" *)
  wire [29:0] trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58067" *)
  wire trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57984" *)
  wire [29:0] trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57988" *)
  wire trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57992" *)
  wire trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57989" *)
  wire [29:0] trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58068" *)
  wire trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57990" *)
  wire [29:0] trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57994" *)
  wire trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57998" *)
  wire trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57995" *)
  wire [29:0] trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58069" *)
  wire trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57996" *)
  wire [29:0] trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58000" *)
  wire trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58004" *)
  wire trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58001" *)
  wire [29:0] trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58070" *)
  wire trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58002" *)
  wire [29:0] trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58006" *)
  wire trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58010" *)
  wire trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58007" *)
  wire [29:0] trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58071" *)
  wire trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58008" *)
  wire [29:0] trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58012" *)
  wire trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58016" *)
  wire trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58013" *)
  wire [29:0] trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58072" *)
  wire trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58014" *)
  wire [29:0] trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58018" *)
  wire trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58022" *)
  wire trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58019" *)
  wire [29:0] trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58073" *)
  wire trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58020" *)
  wire [29:0] trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57969" *)
  wire trt_loop_else_mux_112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57973" *)
  wire trt_loop_else_mux_113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57975" *)
  wire trt_loop_else_mux_114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57979" *)
  wire trt_loop_else_mux_115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57981" *)
  wire trt_loop_else_mux_116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57985" *)
  wire trt_loop_else_mux_117_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57987" *)
  wire trt_loop_else_mux_118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57991" *)
  wire trt_loop_else_mux_119_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57993" *)
  wire trt_loop_else_mux_120_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57997" *)
  wire trt_loop_else_mux_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:57999" *)
  wire trt_loop_else_mux_122_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58003" *)
  wire trt_loop_else_mux_123_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58005" *)
  wire trt_loop_else_mux_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58009" *)
  wire trt_loop_else_mux_125_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58011" *)
  wire trt_loop_else_mux_126_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58015" *)
  wire trt_loop_else_mux_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58017" *)
  wire trt_loop_else_mux_128_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58021" *)
  wire trt_loop_else_mux_129_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58023" *)
  wire trt_loop_else_mux_130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58027" *)
  wire trt_loop_else_mux_131_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58029" *)
  wire trt_loop_else_mux_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58033" *)
  wire trt_loop_else_mux_133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58035" *)
  wire trt_loop_else_mux_134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58039" *)
  wire trt_loop_else_mux_135_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58041" *)
  wire trt_loop_else_mux_136_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58045" *)
  wire trt_loop_else_mux_137_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58047" *)
  wire trt_loop_else_mux_138_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58051" *)
  wire trt_loop_else_mux_139_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58053" *)
  wire trt_loop_else_mux_140_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58057" *)
  wire trt_loop_else_mux_141_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58059" *)
  wire trt_loop_else_mux_142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58063" *)
  wire trt_loop_else_mux_143_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58391" *) trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58431" *) trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58471" *) trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58511" *) trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58551" *) trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58591" *) trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58631" *) trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58671" *) trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58711" *) trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58751" *) trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58791" *) trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58831" *) trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58871" *) trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58911" *) trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58951" *) trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva = { IntShiftRight_49U_6U_32U_mbits_fixed_sva[111], IntShiftRight_49U_6U_32U_mbits_fixed_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58991" *) trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_and_nl;
  assign chn_trt_out_and_2_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58356" *) _0408_;
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58389" *) _0470_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58396" *) _0308_;
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58429" *) _0533_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58436" *) _0311_;
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58469" *) _0596_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58476" *) _0314_;
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58509" *) _0659_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58516" *) _0317_;
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58549" *) _0722_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58556" *) _0320_;
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58589" *) _0785_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58596" *) _0323_;
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58629" *) _0848_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58636" *) _0326_;
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58669" *) _0911_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58676" *) _0329_;
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58709" *) _0974_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58716" *) _0332_;
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58749" *) _1037_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58756" *) _0335_;
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58789" *) _1100_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58796" *) _0338_;
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58829" *) _1163_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58836" *) _0341_;
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58869" *) _1226_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58876" *) _0344_;
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58909" *) _1289_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58916" *) _0347_;
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58949" *) _1352_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58956" *) _0350_;
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_and_nl = IntShiftRight_49U_6U_32U_mbits_fixed_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58989" *) _1415_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58996" *) _0353_;
  assign _0132_ = chn_trt_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58998" *) _1417_;
  assign and_4_mdf = _0132_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58998" *) _1418_;
  assign and_dcpl_1 = chn_trt_out_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58999" *) cfg_mul_shift_value_rsc_triosy_obj_bawt;
  assign and_dcpl_3 = and_dcpl_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59001" *) reg_chn_trt_out_rsci_ld_core_psct_cse;
  assign and_dcpl_7 = or_dcpl_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59003" *) chn_trt_in_rsci_bawt;
  assign and_dcpl_11 = chn_trt_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59004" *) and_dcpl_24;
  assign and_dcpl_15 = or_dcpl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59005" *) or_dcpl_3;
  assign and_dcpl_17 = reg_chn_trt_out_rsci_ld_core_psct_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59006" *) chn_trt_in_rsci_bawt;
  assign and_dcpl_19 = and_dcpl_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59007" *) or_dcpl_3;
  assign _0133_ = cfg_precision[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59008" *) or_dcpl;
  assign _0134_ = cfg_mul_shift_value_rsc_triosy_obj_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59010" *) reg_chn_trt_out_rsci_ld_core_psct_cse;
  assign and_dcpl_23 = _0134_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59010" *) chn_trt_in_rsci_bawt;
  assign and_dcpl_134 = and_dcpl_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59012" *) _0356_;
  assign _0135_ = or_dcpl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59013" *) and_dcpl_7;
  assign and_148_cse = _0135_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59013" *) fsm_output[1];
  assign _0136_ = or_dcpl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59014" *) and_dcpl_11;
  assign and_150_cse = _0136_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59014" *) fsm_output[1];
  assign _0137_ = or_dcpl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59015" *) chn_trt_in_rsci_bawt;
  assign or_tmp_150 = _0137_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59015" *) fsm_output[1];
  assign _0138_ = and_dcpl_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59017" *) and_dcpl_11;
  assign _0139_ = mux_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59019" *) chn_trt_in_rsci_bawt;
  assign _0140_ = _0139_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59019" *) fsm_output[1];
  assign _0141_ = _1420_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59020" *) chn_trt_out_rsci_bawt;
  assign _0142_ = _0141_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59021" *) and_dcpl_23;
  assign _0143_ = mux_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59023" *) chn_trt_in_rsci_bawt;
  assign _0144_ = _0143_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59023" *) fsm_output[1];
  assign _0145_ = _1421_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59024" *) chn_trt_out_rsci_bawt;
  assign _0146_ = _0145_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59025" *) and_dcpl_23;
  assign _0147_ = mux_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59027" *) chn_trt_in_rsci_bawt;
  assign _0148_ = _0147_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59027" *) fsm_output[1];
  assign _0149_ = _1422_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59028" *) chn_trt_out_rsci_bawt;
  assign _0150_ = _0149_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59029" *) and_dcpl_23;
  assign _0151_ = mux_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59031" *) chn_trt_in_rsci_bawt;
  assign _0152_ = _0151_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59031" *) fsm_output[1];
  assign _0153_ = _1423_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59032" *) chn_trt_out_rsci_bawt;
  assign _0154_ = _0153_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59033" *) and_dcpl_23;
  assign _0155_ = mux_8_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59035" *) chn_trt_in_rsci_bawt;
  assign _0156_ = _0155_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59036" *) fsm_output[1];
  assign _0157_ = _1424_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59037" *) chn_trt_out_rsci_bawt;
  assign _0158_ = _0157_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59037" *) and_dcpl_23;
  assign _0159_ = mux_9_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59039" *) chn_trt_in_rsci_bawt;
  assign _0160_ = _0159_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59040" *) fsm_output[1];
  assign _0161_ = _1425_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59041" *) chn_trt_out_rsci_bawt;
  assign _0162_ = _0161_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59041" *) and_dcpl_23;
  assign _0163_ = mux_10_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59043" *) chn_trt_in_rsci_bawt;
  assign _0164_ = _0163_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59044" *) fsm_output[1];
  assign _0165_ = _1426_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59045" *) chn_trt_out_rsci_bawt;
  assign _0166_ = _0165_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59045" *) and_dcpl_23;
  assign _0167_ = mux_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59047" *) chn_trt_in_rsci_bawt;
  assign _0168_ = _0167_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59048" *) fsm_output[1];
  assign _0169_ = _1427_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59049" *) chn_trt_out_rsci_bawt;
  assign _0170_ = _0169_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59049" *) and_dcpl_23;
  assign _0171_ = mux_12_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59051" *) chn_trt_in_rsci_bawt;
  assign _0172_ = _0171_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59052" *) fsm_output[1];
  assign _0173_ = _1428_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59053" *) chn_trt_out_rsci_bawt;
  assign _0174_ = _0173_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59053" *) and_dcpl_23;
  assign _0175_ = mux_13_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59055" *) chn_trt_in_rsci_bawt;
  assign _0176_ = _0175_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59056" *) fsm_output[1];
  assign _0177_ = _1429_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59057" *) chn_trt_out_rsci_bawt;
  assign _0178_ = _0177_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59057" *) and_dcpl_23;
  assign _0179_ = mux_14_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59059" *) chn_trt_in_rsci_bawt;
  assign _0180_ = _0179_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59060" *) fsm_output[1];
  assign _0181_ = _1430_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59061" *) chn_trt_out_rsci_bawt;
  assign _0182_ = _0181_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59061" *) and_dcpl_23;
  assign _0183_ = mux_15_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59063" *) chn_trt_in_rsci_bawt;
  assign _0184_ = _0183_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59064" *) fsm_output[1];
  assign _0185_ = _1431_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59065" *) chn_trt_out_rsci_bawt;
  assign _0186_ = _0185_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59065" *) and_dcpl_23;
  assign _0187_ = mux_16_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59067" *) chn_trt_in_rsci_bawt;
  assign _0188_ = _0187_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59068" *) fsm_output[1];
  assign _0189_ = _1432_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59069" *) chn_trt_out_rsci_bawt;
  assign _0190_ = _0189_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59069" *) and_dcpl_23;
  assign _0191_ = mux_17_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59071" *) chn_trt_in_rsci_bawt;
  assign _0192_ = _0191_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59072" *) fsm_output[1];
  assign _0193_ = _1433_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59073" *) chn_trt_out_rsci_bawt;
  assign _0194_ = _0193_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59073" *) and_dcpl_23;
  assign _0195_ = mux_18_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59075" *) chn_trt_in_rsci_bawt;
  assign _0196_ = _0195_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59076" *) fsm_output[1];
  assign _0197_ = _1434_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59077" *) chn_trt_out_rsci_bawt;
  assign _0198_ = _0197_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59077" *) and_dcpl_23;
  assign _0199_ = mux_19_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59079" *) chn_trt_in_rsci_bawt;
  assign _0200_ = _0199_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59080" *) fsm_output[1];
  assign _0201_ = _1435_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59081" *) chn_trt_out_rsci_bawt;
  assign _0202_ = _0201_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59081" *) and_dcpl_23;
  assign _0203_ = _0357_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59090" *) fsm_output[1];
  assign _0204_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59098" *) chn_trt_in_rsci_ld_core_psct_mx0c0;
  assign _0205_ = and_dcpl_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59106" *) and_dcpl_7;
  assign _0206_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59107" *) _1437_;
  assign _0207_ = and_dcpl_15 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59116" *) chn_trt_in_rsci_bawt;
  assign _0208_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *) _0359_;
  assign _0209_ = _0208_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *) fsm_output[1];
  assign _0210_ = and_dcpl_19 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *) and_dcpl_17;
  assign _0211_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59117" *) _0359_;
  assign _0212_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59118" *) _1439_;
  assign _0213_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59227" *) _0360_;
  assign _0214_ = _0213_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59227" *) fsm_output[1];
  assign _0215_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59227" *) _0360_;
  assign _0216_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59228" *) _1441_;
  assign _0217_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59238" *) _0361_;
  assign _0218_ = _0217_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59238" *) fsm_output[1];
  assign _0219_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59238" *) _0361_;
  assign _0220_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59239" *) _1443_;
  assign _0221_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59249" *) _0362_;
  assign _0222_ = _0221_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59249" *) fsm_output[1];
  assign _0223_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59249" *) _0362_;
  assign _0224_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59250" *) _1445_;
  assign _0225_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59260" *) _0363_;
  assign _0226_ = _0225_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59260" *) fsm_output[1];
  assign _0227_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59260" *) _0363_;
  assign _0228_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59261" *) _1447_;
  assign _0229_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59271" *) _0364_;
  assign _0230_ = _0229_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59271" *) fsm_output[1];
  assign _0231_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59271" *) _0364_;
  assign _0232_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59272" *) _1449_;
  assign _0233_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59282" *) _0365_;
  assign _0234_ = _0233_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59282" *) fsm_output[1];
  assign _0235_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59282" *) _0365_;
  assign _0236_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59283" *) _1451_;
  assign _0237_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59293" *) _0366_;
  assign _0238_ = _0237_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59293" *) fsm_output[1];
  assign _0239_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59293" *) _0366_;
  assign _0240_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59294" *) _1453_;
  assign _0241_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59304" *) _0367_;
  assign _0242_ = _0241_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59304" *) fsm_output[1];
  assign _0243_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59304" *) _0367_;
  assign _0244_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59305" *) _1455_;
  assign _0245_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59315" *) _0368_;
  assign _0246_ = _0245_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59315" *) fsm_output[1];
  assign _0247_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59315" *) _0368_;
  assign _0248_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59316" *) _1457_;
  assign _0249_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59326" *) _0369_;
  assign _0250_ = _0249_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59326" *) fsm_output[1];
  assign _0251_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59326" *) _0369_;
  assign _0252_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59327" *) _1459_;
  assign _0253_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59337" *) _0370_;
  assign _0254_ = _0253_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59337" *) fsm_output[1];
  assign _0255_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59337" *) _0370_;
  assign _0256_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59338" *) _1461_;
  assign _0257_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59348" *) _0371_;
  assign _0258_ = _0257_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59348" *) fsm_output[1];
  assign _0259_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59348" *) _0371_;
  assign _0260_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59349" *) _1463_;
  assign _0261_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59359" *) _0372_;
  assign _0262_ = _0261_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59359" *) fsm_output[1];
  assign _0263_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59359" *) _0372_;
  assign _0264_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59360" *) _1465_;
  assign _0265_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59370" *) _0373_;
  assign _0266_ = _0265_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59370" *) fsm_output[1];
  assign _0267_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59370" *) _0373_;
  assign _0268_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59371" *) _1467_;
  assign _0269_ = _0207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59381" *) _0374_;
  assign _0270_ = _0269_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59381" *) fsm_output[1];
  assign _0271_ = _0210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59381" *) _0374_;
  assign _0272_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59382" *) _1469_;
  assign _0273_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59391" *) _1470_;
  assign _0274_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58396" *) 18'b111111111111111111;
  assign _0275_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58436" *) 18'b111111111111111111;
  assign _0276_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58476" *) 18'b111111111111111111;
  assign _0277_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58516" *) 18'b111111111111111111;
  assign _0278_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58556" *) 18'b111111111111111111;
  assign _0279_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58596" *) 18'b111111111111111111;
  assign _0280_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58636" *) 18'b111111111111111111;
  assign _0281_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58676" *) 18'b111111111111111111;
  assign _0282_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58716" *) 18'b111111111111111111;
  assign _0283_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58756" *) 18'b111111111111111111;
  assign _0284_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58796" *) 18'b111111111111111111;
  assign _0285_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58836" *) 18'b111111111111111111;
  assign _0286_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58876" *) 18'b111111111111111111;
  assign _0287_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58916" *) 18'b111111111111111111;
  assign _0288_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58956" *) 18'b111111111111111111;
  assign _0289_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[48:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58996" *) 18'b111111111111111111;
  assign and_dcpl_24 = cfg_precision == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59004" *) 2'b10;
  assign _0290_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58394" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[48:31];
  assign _0291_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58434" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[48:31];
  assign _0292_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58474" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[48:31];
  assign _0293_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58514" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[48:31];
  assign _0294_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58554" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[48:31];
  assign _0295_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58594" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[48:31];
  assign _0296_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58634" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[48:31];
  assign _0297_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58674" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[48:31];
  assign _0298_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58714" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[48:31];
  assign _0299_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58754" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[48:31];
  assign _0300_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58794" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[48:31];
  assign _0301_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58834" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[48:31];
  assign _0302_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58874" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[48:31];
  assign _0303_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58914" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[48:31];
  assign _0304_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58954" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[48:31];
  assign _0305_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58994" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[48:31];
  assign or_dcpl_3 = cfg_precision != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59002" *) 2'b10;
  assign _0306_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58389" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[111];
  assign _0307_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58394" *) _0290_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58394" *) _0471_;
  assign _0308_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58396" *) _0274_;
  assign _0309_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58429" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[111];
  assign _0310_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58434" *) _0291_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58434" *) _0534_;
  assign _0311_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58436" *) _0275_;
  assign _0312_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58469" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[111];
  assign _0313_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58474" *) _0292_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58474" *) _0597_;
  assign _0314_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58476" *) _0276_;
  assign _0315_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58509" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[111];
  assign _0316_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58514" *) _0293_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58514" *) _0660_;
  assign _0317_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58516" *) _0277_;
  assign _0318_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58549" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[111];
  assign _0319_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58554" *) _0294_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58554" *) _0723_;
  assign _0320_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58556" *) _0278_;
  assign _0321_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58589" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[111];
  assign _0322_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58594" *) _0295_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58594" *) _0786_;
  assign _0323_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58596" *) _0279_;
  assign _0324_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58629" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[111];
  assign _0325_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58634" *) _0296_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58634" *) _0849_;
  assign _0326_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58636" *) _0280_;
  assign _0327_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58669" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[111];
  assign _0328_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58674" *) _0297_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58674" *) _0912_;
  assign _0329_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58676" *) _0281_;
  assign _0330_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58709" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[111];
  assign _0331_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58714" *) _0298_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58714" *) _0975_;
  assign _0332_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58716" *) _0282_;
  assign _0333_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58749" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[111];
  assign _0334_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58754" *) _0299_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58754" *) _1038_;
  assign _0335_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58756" *) _0283_;
  assign _0336_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58789" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[111];
  assign _0337_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58794" *) _0300_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58794" *) _1101_;
  assign _0338_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58796" *) _0284_;
  assign _0339_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58829" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[111];
  assign _0340_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58834" *) _0301_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58834" *) _1164_;
  assign _0341_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58836" *) _0285_;
  assign _0342_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58869" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[111];
  assign _0343_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58874" *) _0302_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58874" *) _1227_;
  assign _0344_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58876" *) _0286_;
  assign _0345_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58909" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[111];
  assign _0346_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58914" *) _0303_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58914" *) _1290_;
  assign _0347_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58916" *) _0287_;
  assign _0348_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58949" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[111];
  assign _0349_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58954" *) _0304_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58954" *) _1353_;
  assign _0350_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58956" *) _0288_;
  assign _0351_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58989" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[111];
  assign _0352_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58994" *) _0305_;
  assign IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58994" *) _1416_;
  assign _0353_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58996" *) _0289_;
  assign _0354_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58997" *) reg_chn_trt_out_rsci_ld_core_psct_cse;
  assign _0355_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59008" *) _0133_;
  assign not_tmp_9 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59008" *) _1419_;
  assign _0356_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59012" *) chn_trt_in_rsci_bawt;
  assign _0357_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59090" *) and_4_mdf;
  assign _0358_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59090" *) _0203_;
  assign _0359_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59116" *) chn_trt_in_rsci_d_mxwt[784];
  assign _0360_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59226" *) chn_trt_in_rsci_d_mxwt[785];
  assign _0361_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59237" *) chn_trt_in_rsci_d_mxwt[786];
  assign _0362_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59248" *) chn_trt_in_rsci_d_mxwt[787];
  assign _0363_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59259" *) chn_trt_in_rsci_d_mxwt[788];
  assign _0364_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59270" *) chn_trt_in_rsci_d_mxwt[789];
  assign _0365_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59281" *) chn_trt_in_rsci_d_mxwt[790];
  assign _0366_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59292" *) chn_trt_in_rsci_d_mxwt[791];
  assign _0367_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59303" *) chn_trt_in_rsci_d_mxwt[792];
  assign _0368_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59314" *) chn_trt_in_rsci_d_mxwt[793];
  assign _0369_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59325" *) chn_trt_in_rsci_d_mxwt[794];
  assign _0370_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59336" *) chn_trt_in_rsci_d_mxwt[795];
  assign _0371_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59347" *) chn_trt_in_rsci_d_mxwt[796];
  assign _0372_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59358" *) chn_trt_in_rsci_d_mxwt[797];
  assign _0373_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59369" *) chn_trt_in_rsci_d_mxwt[798];
  assign _0374_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59380" *) chn_trt_in_rsci_d_mxwt[799];
  assign _0375_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59392" *) and_dcpl_134;
  assign _0376_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59396" *) _1471_;
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59397" *) _1472_;
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59401" *) _0000_;
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59404" *) _0001_;
  assign _0377_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59406" *) _1473_;
  assign trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59407" *) _1474_;
  assign _0378_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59411" *) _1475_;
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59412" *) _1476_;
  assign _0379_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59416" *) _1477_;
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59417" *) _1478_;
  assign _0380_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59421" *) _1479_;
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59422" *) _1480_;
  assign _0381_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59426" *) _1481_;
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59427" *) _1482_;
  assign _0382_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59431" *) _1483_;
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59432" *) _1484_;
  assign _0383_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59436" *) _1485_;
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59437" *) _1486_;
  assign _0384_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59441" *) _1487_;
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59442" *) _1488_;
  assign _0385_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59446" *) _1489_;
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59447" *) _1490_;
  assign _0386_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59451" *) _1491_;
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59452" *) _1492_;
  assign _0387_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59456" *) _1493_;
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59457" *) _1494_;
  assign _0388_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59461" *) _1495_;
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59462" *) _1496_;
  assign _0389_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59466" *) _1497_;
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59467" *) _1498_;
  assign _0390_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59471" *) _1499_;
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59472" *) _1500_;
  assign _0391_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59476" *) _1501_;
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59477" *) _1502_;
  assign _0392_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59481" *) _1503_;
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59482" *) _1504_;
  assign _0393_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59486" *) _1505_;
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59487" *) _1506_;
  assign _0394_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59491" *) _1507_;
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59492" *) _1508_;
  assign _0395_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59496" *) _1509_;
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59497" *) _1510_;
  assign _0396_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59501" *) _1511_;
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59502" *) _1512_;
  assign _0397_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59506" *) _1513_;
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59507" *) _1514_;
  assign _0398_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59511" *) _1515_;
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59512" *) _1516_;
  assign _0399_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59516" *) _1517_;
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59517" *) _1518_;
  assign _0400_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59521" *) _1519_;
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59522" *) _1520_;
  assign _0401_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59526" *) _1521_;
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59527" *) _1522_;
  assign _0402_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59531" *) _1523_;
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59532" *) _1524_;
  assign _0403_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59536" *) _1525_;
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59537" *) _1526_;
  assign _0404_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59541" *) _1527_;
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59542" *) _1528_;
  assign _0405_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59546" *) _1529_;
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59547" *) _1530_;
  assign _0406_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59551" *) _1531_;
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59552" *) _1532_;
  assign _0407_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59556" *) _1533_;
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59557" *) _1534_;
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59561" *) _0002_;
  assign trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59564" *) _0003_;
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59566" *) _0004_;
  assign trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59569" *) _0005_;
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59571" *) _0006_;
  assign trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59574" *) _0007_;
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59576" *) _0008_;
  assign trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59579" *) _0009_;
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59581" *) _0010_;
  assign trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59584" *) _0011_;
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59586" *) _0012_;
  assign trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59589" *) _0013_;
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59591" *) _0014_;
  assign trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59594" *) _0015_;
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59596" *) _0016_;
  assign trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59599" *) _0017_;
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59601" *) _0018_;
  assign trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59604" *) _0019_;
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59606" *) _0020_;
  assign trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59609" *) _0021_;
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59611" *) _0022_;
  assign trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59614" *) _0023_;
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59616" *) _0024_;
  assign trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59619" *) _0025_;
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59621" *) _0026_;
  assign trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59624" *) _0027_;
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59626" *) _0028_;
  assign trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59629" *) _0029_;
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59631" *) _0030_;
  assign trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59634" *) _0031_;
  assign _0408_ = and_148_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58356" *) and_150_cse;
  assign _0409_ = IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58359" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[1];
  assign _0410_ = _0409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58359" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[2];
  assign _0411_ = _0410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58360" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[3];
  assign _0412_ = _0411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58360" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[4];
  assign _0413_ = _0412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58361" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[5];
  assign _0414_ = _0413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58361" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[6];
  assign _0415_ = _0414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58362" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[7];
  assign _0416_ = _0415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58362" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[8];
  assign _0417_ = _0416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58363" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[9];
  assign _0418_ = _0417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58363" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[10];
  assign _0419_ = _0418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58364" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[11];
  assign _0420_ = _0419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58364" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[12];
  assign _0421_ = _0420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58365" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[13];
  assign _0422_ = _0421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58365" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[14];
  assign _0423_ = _0422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58366" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[15];
  assign _0424_ = _0423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58366" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[16];
  assign _0425_ = _0424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58367" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[17];
  assign _0426_ = _0425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58367" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[18];
  assign _0427_ = _0426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58368" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[19];
  assign _0428_ = _0427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58368" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[20];
  assign _0429_ = _0428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58369" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[21];
  assign _0430_ = _0429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58369" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[22];
  assign _0431_ = _0430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58370" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[23];
  assign _0432_ = _0431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58370" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[24];
  assign _0433_ = _0432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58371" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[25];
  assign _0434_ = _0433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58371" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[26];
  assign _0435_ = _0434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58372" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[27];
  assign _0436_ = _0435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58372" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[28];
  assign _0437_ = _0436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58373" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[29];
  assign _0438_ = _0437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58373" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[30];
  assign _0439_ = _0438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58374" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[31];
  assign _0440_ = _0439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58374" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[32];
  assign _0441_ = _0440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58375" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[33];
  assign _0442_ = _0441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58375" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[34];
  assign _0443_ = _0442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58376" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[35];
  assign _0444_ = _0443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58376" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[36];
  assign _0445_ = _0444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58377" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[37];
  assign _0446_ = _0445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58377" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[38];
  assign _0447_ = _0446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58378" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[39];
  assign _0448_ = _0447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58378" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[40];
  assign _0449_ = _0448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58379" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[41];
  assign _0450_ = _0449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58379" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[42];
  assign _0451_ = _0450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58380" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[43];
  assign _0452_ = _0451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58380" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[44];
  assign _0453_ = _0452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58381" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[45];
  assign _0454_ = _0453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58381" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[46];
  assign _0455_ = _0454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58382" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[47];
  assign _0456_ = _0455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58382" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[48];
  assign _0457_ = _0456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58383" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[49];
  assign _0458_ = _0457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58383" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[50];
  assign _0459_ = _0458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58384" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[51];
  assign _0460_ = _0459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58384" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[52];
  assign _0461_ = _0460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58385" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[53];
  assign _0462_ = _0461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58385" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[54];
  assign _0463_ = _0462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58386" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[55];
  assign _0464_ = _0463_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58386" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[56];
  assign _0465_ = _0464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58387" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[57];
  assign _0466_ = _0465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58387" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[58];
  assign _0467_ = _0466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58388" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[59];
  assign _0468_ = _0467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58388" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[60];
  assign _0469_ = _0468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58389" *) IntShiftRight_49U_6U_32U_mbits_fixed_1_sva[61];
  assign _0470_ = _0469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58389" *) _0306_;
  assign _0471_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58394" *) _0307_;
  assign _0472_ = IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58399" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[1];
  assign _0473_ = _0472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58399" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[2];
  assign _0474_ = _0473_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58400" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[3];
  assign _0475_ = _0474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58400" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[4];
  assign _0476_ = _0475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58401" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[5];
  assign _0477_ = _0476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58401" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[6];
  assign _0478_ = _0477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58402" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[7];
  assign _0479_ = _0478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58402" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[8];
  assign _0480_ = _0479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58403" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[9];
  assign _0481_ = _0480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58403" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[10];
  assign _0482_ = _0481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58404" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[11];
  assign _0483_ = _0482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58404" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[12];
  assign _0484_ = _0483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58405" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[13];
  assign _0485_ = _0484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58405" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[14];
  assign _0486_ = _0485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58406" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[15];
  assign _0487_ = _0486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58406" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[16];
  assign _0488_ = _0487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58407" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[17];
  assign _0489_ = _0488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58407" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[18];
  assign _0490_ = _0489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58408" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[19];
  assign _0491_ = _0490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58408" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[20];
  assign _0492_ = _0491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58409" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[21];
  assign _0493_ = _0492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58409" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[22];
  assign _0494_ = _0493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58410" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[23];
  assign _0495_ = _0494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58410" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[24];
  assign _0496_ = _0495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58411" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[25];
  assign _0497_ = _0496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58411" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[26];
  assign _0498_ = _0497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58412" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[27];
  assign _0499_ = _0498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58412" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[28];
  assign _0500_ = _0499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58413" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[29];
  assign _0501_ = _0500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58413" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[30];
  assign _0502_ = _0501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58414" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[31];
  assign _0503_ = _0502_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58414" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[32];
  assign _0504_ = _0503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58415" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[33];
  assign _0505_ = _0504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58415" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[34];
  assign _0506_ = _0505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58416" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[35];
  assign _0507_ = _0506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58416" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[36];
  assign _0508_ = _0507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58417" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[37];
  assign _0509_ = _0508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58417" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[38];
  assign _0510_ = _0509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58418" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[39];
  assign _0511_ = _0510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58418" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[40];
  assign _0512_ = _0511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58419" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[41];
  assign _0513_ = _0512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58419" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[42];
  assign _0514_ = _0513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58420" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[43];
  assign _0515_ = _0514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58420" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[44];
  assign _0516_ = _0515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58421" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[45];
  assign _0517_ = _0516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58421" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[46];
  assign _0518_ = _0517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58422" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[47];
  assign _0519_ = _0518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58422" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[48];
  assign _0520_ = _0519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58423" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[49];
  assign _0521_ = _0520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58423" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[50];
  assign _0522_ = _0521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58424" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[51];
  assign _0523_ = _0522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58424" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[52];
  assign _0524_ = _0523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58425" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[53];
  assign _0525_ = _0524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58425" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[54];
  assign _0526_ = _0525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58426" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[55];
  assign _0527_ = _0526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58426" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[56];
  assign _0528_ = _0527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58427" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[57];
  assign _0529_ = _0528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58427" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[58];
  assign _0530_ = _0529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58428" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[59];
  assign _0531_ = _0530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58428" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[60];
  assign _0532_ = _0531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58429" *) IntShiftRight_49U_6U_32U_mbits_fixed_2_sva[61];
  assign _0533_ = _0532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58429" *) _0309_;
  assign _0534_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58434" *) _0310_;
  assign _0535_ = IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58439" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[1];
  assign _0536_ = _0535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58439" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[2];
  assign _0537_ = _0536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58440" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[3];
  assign _0538_ = _0537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58440" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[4];
  assign _0539_ = _0538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58441" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[5];
  assign _0540_ = _0539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58441" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[6];
  assign _0541_ = _0540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58442" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[7];
  assign _0542_ = _0541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58442" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[8];
  assign _0543_ = _0542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58443" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[9];
  assign _0544_ = _0543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58443" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[10];
  assign _0545_ = _0544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58444" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[11];
  assign _0546_ = _0545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58444" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[12];
  assign _0547_ = _0546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58445" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[13];
  assign _0548_ = _0547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58445" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[14];
  assign _0549_ = _0548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58446" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[15];
  assign _0550_ = _0549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58446" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[16];
  assign _0551_ = _0550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58447" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[17];
  assign _0552_ = _0551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58447" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[18];
  assign _0553_ = _0552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58448" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[19];
  assign _0554_ = _0553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58448" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[20];
  assign _0555_ = _0554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58449" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[21];
  assign _0556_ = _0555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58449" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[22];
  assign _0557_ = _0556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58450" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[23];
  assign _0558_ = _0557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58450" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[24];
  assign _0559_ = _0558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58451" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[25];
  assign _0560_ = _0559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58451" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[26];
  assign _0561_ = _0560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58452" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[27];
  assign _0562_ = _0561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58452" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[28];
  assign _0563_ = _0562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58453" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[29];
  assign _0564_ = _0563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58453" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[30];
  assign _0565_ = _0564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58454" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[31];
  assign _0566_ = _0565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58454" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[32];
  assign _0567_ = _0566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58455" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[33];
  assign _0568_ = _0567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58455" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[34];
  assign _0569_ = _0568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58456" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[35];
  assign _0570_ = _0569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58456" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[36];
  assign _0571_ = _0570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58457" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[37];
  assign _0572_ = _0571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58457" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[38];
  assign _0573_ = _0572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58458" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[39];
  assign _0574_ = _0573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58458" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[40];
  assign _0575_ = _0574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58459" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[41];
  assign _0576_ = _0575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58459" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[42];
  assign _0577_ = _0576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58460" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[43];
  assign _0578_ = _0577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58460" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[44];
  assign _0579_ = _0578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58461" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[45];
  assign _0580_ = _0579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58461" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[46];
  assign _0581_ = _0580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58462" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[47];
  assign _0582_ = _0581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58462" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[48];
  assign _0583_ = _0582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58463" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[49];
  assign _0584_ = _0583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58463" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[50];
  assign _0585_ = _0584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58464" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[51];
  assign _0586_ = _0585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58464" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[52];
  assign _0587_ = _0586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58465" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[53];
  assign _0588_ = _0587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58465" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[54];
  assign _0589_ = _0588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58466" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[55];
  assign _0590_ = _0589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58466" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[56];
  assign _0591_ = _0590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58467" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[57];
  assign _0592_ = _0591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58467" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[58];
  assign _0593_ = _0592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58468" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[59];
  assign _0594_ = _0593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58468" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[60];
  assign _0595_ = _0594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58469" *) IntShiftRight_49U_6U_32U_mbits_fixed_3_sva[61];
  assign _0596_ = _0595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58469" *) _0312_;
  assign _0597_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58474" *) _0313_;
  assign _0598_ = IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58479" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[1];
  assign _0599_ = _0598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58479" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[2];
  assign _0600_ = _0599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58480" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[3];
  assign _0601_ = _0600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58480" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[4];
  assign _0602_ = _0601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58481" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[5];
  assign _0603_ = _0602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58481" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[6];
  assign _0604_ = _0603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58482" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[7];
  assign _0605_ = _0604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58482" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[8];
  assign _0606_ = _0605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58483" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[9];
  assign _0607_ = _0606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58483" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[10];
  assign _0608_ = _0607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58484" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[11];
  assign _0609_ = _0608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58484" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[12];
  assign _0610_ = _0609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58485" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[13];
  assign _0611_ = _0610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58485" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[14];
  assign _0612_ = _0611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58486" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[15];
  assign _0613_ = _0612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58486" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[16];
  assign _0614_ = _0613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58487" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[17];
  assign _0615_ = _0614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58487" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[18];
  assign _0616_ = _0615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58488" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[19];
  assign _0617_ = _0616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58488" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[20];
  assign _0618_ = _0617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58489" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[21];
  assign _0619_ = _0618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58489" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[22];
  assign _0620_ = _0619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58490" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[23];
  assign _0621_ = _0620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58490" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[24];
  assign _0622_ = _0621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58491" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[25];
  assign _0623_ = _0622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58491" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[26];
  assign _0624_ = _0623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58492" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[27];
  assign _0625_ = _0624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58492" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[28];
  assign _0626_ = _0625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58493" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[29];
  assign _0627_ = _0626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58493" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[30];
  assign _0628_ = _0627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58494" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[31];
  assign _0629_ = _0628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58494" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[32];
  assign _0630_ = _0629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58495" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[33];
  assign _0631_ = _0630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58495" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[34];
  assign _0632_ = _0631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58496" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[35];
  assign _0633_ = _0632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58496" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[36];
  assign _0634_ = _0633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58497" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[37];
  assign _0635_ = _0634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58497" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[38];
  assign _0636_ = _0635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58498" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[39];
  assign _0637_ = _0636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58498" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[40];
  assign _0638_ = _0637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58499" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[41];
  assign _0639_ = _0638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58499" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[42];
  assign _0640_ = _0639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58500" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[43];
  assign _0641_ = _0640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58500" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[44];
  assign _0642_ = _0641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58501" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[45];
  assign _0643_ = _0642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58501" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[46];
  assign _0644_ = _0643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58502" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[47];
  assign _0645_ = _0644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58502" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[48];
  assign _0646_ = _0645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58503" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[49];
  assign _0647_ = _0646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58503" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[50];
  assign _0648_ = _0647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58504" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[51];
  assign _0649_ = _0648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58504" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[52];
  assign _0650_ = _0649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58505" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[53];
  assign _0651_ = _0650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58505" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[54];
  assign _0652_ = _0651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58506" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[55];
  assign _0653_ = _0652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58506" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[56];
  assign _0654_ = _0653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58507" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[57];
  assign _0655_ = _0654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58507" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[58];
  assign _0656_ = _0655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58508" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[59];
  assign _0657_ = _0656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58508" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[60];
  assign _0658_ = _0657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58509" *) IntShiftRight_49U_6U_32U_mbits_fixed_4_sva[61];
  assign _0659_ = _0658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58509" *) _0315_;
  assign _0660_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58514" *) _0316_;
  assign _0661_ = IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58519" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[1];
  assign _0662_ = _0661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58519" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[2];
  assign _0663_ = _0662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58520" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[3];
  assign _0664_ = _0663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58520" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[4];
  assign _0665_ = _0664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58521" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[5];
  assign _0666_ = _0665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58521" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[6];
  assign _0667_ = _0666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58522" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[7];
  assign _0668_ = _0667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58522" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[8];
  assign _0669_ = _0668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58523" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[9];
  assign _0670_ = _0669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58523" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[10];
  assign _0671_ = _0670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58524" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[11];
  assign _0672_ = _0671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58524" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[12];
  assign _0673_ = _0672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58525" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[13];
  assign _0674_ = _0673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58525" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[14];
  assign _0675_ = _0674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58526" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[15];
  assign _0676_ = _0675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58526" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[16];
  assign _0677_ = _0676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58527" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[17];
  assign _0678_ = _0677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58527" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[18];
  assign _0679_ = _0678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58528" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[19];
  assign _0680_ = _0679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58528" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[20];
  assign _0681_ = _0680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58529" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[21];
  assign _0682_ = _0681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58529" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[22];
  assign _0683_ = _0682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58530" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[23];
  assign _0684_ = _0683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58530" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[24];
  assign _0685_ = _0684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58531" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[25];
  assign _0686_ = _0685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58531" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[26];
  assign _0687_ = _0686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58532" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[27];
  assign _0688_ = _0687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58532" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[28];
  assign _0689_ = _0688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58533" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[29];
  assign _0690_ = _0689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58533" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[30];
  assign _0691_ = _0690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58534" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[31];
  assign _0692_ = _0691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58534" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[32];
  assign _0693_ = _0692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58535" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[33];
  assign _0694_ = _0693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58535" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[34];
  assign _0695_ = _0694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58536" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[35];
  assign _0696_ = _0695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58536" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[36];
  assign _0697_ = _0696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58537" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[37];
  assign _0698_ = _0697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58537" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[38];
  assign _0699_ = _0698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58538" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[39];
  assign _0700_ = _0699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58538" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[40];
  assign _0701_ = _0700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58539" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[41];
  assign _0702_ = _0701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58539" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[42];
  assign _0703_ = _0702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58540" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[43];
  assign _0704_ = _0703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58540" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[44];
  assign _0705_ = _0704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58541" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[45];
  assign _0706_ = _0705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58541" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[46];
  assign _0707_ = _0706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58542" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[47];
  assign _0708_ = _0707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58542" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[48];
  assign _0709_ = _0708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58543" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[49];
  assign _0710_ = _0709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58543" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[50];
  assign _0711_ = _0710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58544" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[51];
  assign _0712_ = _0711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58544" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[52];
  assign _0713_ = _0712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58545" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[53];
  assign _0714_ = _0713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58545" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[54];
  assign _0715_ = _0714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58546" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[55];
  assign _0716_ = _0715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58546" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[56];
  assign _0717_ = _0716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58547" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[57];
  assign _0718_ = _0717_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58547" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[58];
  assign _0719_ = _0718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58548" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[59];
  assign _0720_ = _0719_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58548" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[60];
  assign _0721_ = _0720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58549" *) IntShiftRight_49U_6U_32U_mbits_fixed_5_sva[61];
  assign _0722_ = _0721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58549" *) _0318_;
  assign _0723_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58554" *) _0319_;
  assign _0724_ = IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58559" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[1];
  assign _0725_ = _0724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58559" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[2];
  assign _0726_ = _0725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58560" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[3];
  assign _0727_ = _0726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58560" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[4];
  assign _0728_ = _0727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58561" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[5];
  assign _0729_ = _0728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58561" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[6];
  assign _0730_ = _0729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58562" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[7];
  assign _0731_ = _0730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58562" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[8];
  assign _0732_ = _0731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58563" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[9];
  assign _0733_ = _0732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58563" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[10];
  assign _0734_ = _0733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58564" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[11];
  assign _0735_ = _0734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58564" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[12];
  assign _0736_ = _0735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58565" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[13];
  assign _0737_ = _0736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58565" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[14];
  assign _0738_ = _0737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58566" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[15];
  assign _0739_ = _0738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58566" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[16];
  assign _0740_ = _0739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58567" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[17];
  assign _0741_ = _0740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58567" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[18];
  assign _0742_ = _0741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58568" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[19];
  assign _0743_ = _0742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58568" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[20];
  assign _0744_ = _0743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58569" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[21];
  assign _0745_ = _0744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58569" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[22];
  assign _0746_ = _0745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58570" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[23];
  assign _0747_ = _0746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58570" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[24];
  assign _0748_ = _0747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58571" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[25];
  assign _0749_ = _0748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58571" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[26];
  assign _0750_ = _0749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58572" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[27];
  assign _0751_ = _0750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58572" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[28];
  assign _0752_ = _0751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58573" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[29];
  assign _0753_ = _0752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58573" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[30];
  assign _0754_ = _0753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58574" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[31];
  assign _0755_ = _0754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58574" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[32];
  assign _0756_ = _0755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58575" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[33];
  assign _0757_ = _0756_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58575" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[34];
  assign _0758_ = _0757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58576" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[35];
  assign _0759_ = _0758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58576" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[36];
  assign _0760_ = _0759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58577" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[37];
  assign _0761_ = _0760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58577" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[38];
  assign _0762_ = _0761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58578" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[39];
  assign _0763_ = _0762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58578" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[40];
  assign _0764_ = _0763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58579" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[41];
  assign _0765_ = _0764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58579" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[42];
  assign _0766_ = _0765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58580" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[43];
  assign _0767_ = _0766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58580" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[44];
  assign _0768_ = _0767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58581" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[45];
  assign _0769_ = _0768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58581" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[46];
  assign _0770_ = _0769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58582" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[47];
  assign _0771_ = _0770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58582" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[48];
  assign _0772_ = _0771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58583" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[49];
  assign _0773_ = _0772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58583" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[50];
  assign _0774_ = _0773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58584" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[51];
  assign _0775_ = _0774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58584" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[52];
  assign _0776_ = _0775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58585" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[53];
  assign _0777_ = _0776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58585" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[54];
  assign _0778_ = _0777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58586" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[55];
  assign _0779_ = _0778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58586" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[56];
  assign _0780_ = _0779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58587" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[57];
  assign _0781_ = _0780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58587" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[58];
  assign _0782_ = _0781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58588" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[59];
  assign _0783_ = _0782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58588" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[60];
  assign _0784_ = _0783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58589" *) IntShiftRight_49U_6U_32U_mbits_fixed_6_sva[61];
  assign _0785_ = _0784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58589" *) _0321_;
  assign _0786_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58594" *) _0322_;
  assign _0787_ = IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58599" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[1];
  assign _0788_ = _0787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58599" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[2];
  assign _0789_ = _0788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58600" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[3];
  assign _0790_ = _0789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58600" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[4];
  assign _0791_ = _0790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58601" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[5];
  assign _0792_ = _0791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58601" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[6];
  assign _0793_ = _0792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58602" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[7];
  assign _0794_ = _0793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58602" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[8];
  assign _0795_ = _0794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58603" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[9];
  assign _0796_ = _0795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58603" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[10];
  assign _0797_ = _0796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58604" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[11];
  assign _0798_ = _0797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58604" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[12];
  assign _0799_ = _0798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58605" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[13];
  assign _0800_ = _0799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58605" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[14];
  assign _0801_ = _0800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58606" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[15];
  assign _0802_ = _0801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58606" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[16];
  assign _0803_ = _0802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58607" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[17];
  assign _0804_ = _0803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58607" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[18];
  assign _0805_ = _0804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58608" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[19];
  assign _0806_ = _0805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58608" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[20];
  assign _0807_ = _0806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58609" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[21];
  assign _0808_ = _0807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58609" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[22];
  assign _0809_ = _0808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58610" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[23];
  assign _0810_ = _0809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58610" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[24];
  assign _0811_ = _0810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58611" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[25];
  assign _0812_ = _0811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58611" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[26];
  assign _0813_ = _0812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58612" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[27];
  assign _0814_ = _0813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58612" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[28];
  assign _0815_ = _0814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58613" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[29];
  assign _0816_ = _0815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58613" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[30];
  assign _0817_ = _0816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58614" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[31];
  assign _0818_ = _0817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58614" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[32];
  assign _0819_ = _0818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58615" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[33];
  assign _0820_ = _0819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58615" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[34];
  assign _0821_ = _0820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58616" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[35];
  assign _0822_ = _0821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58616" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[36];
  assign _0823_ = _0822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58617" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[37];
  assign _0824_ = _0823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58617" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[38];
  assign _0825_ = _0824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58618" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[39];
  assign _0826_ = _0825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58618" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[40];
  assign _0827_ = _0826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58619" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[41];
  assign _0828_ = _0827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58619" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[42];
  assign _0829_ = _0828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58620" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[43];
  assign _0830_ = _0829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58620" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[44];
  assign _0831_ = _0830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58621" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[45];
  assign _0832_ = _0831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58621" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[46];
  assign _0833_ = _0832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58622" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[47];
  assign _0834_ = _0833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58622" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[48];
  assign _0835_ = _0834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58623" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[49];
  assign _0836_ = _0835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58623" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[50];
  assign _0837_ = _0836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58624" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[51];
  assign _0838_ = _0837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58624" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[52];
  assign _0839_ = _0838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58625" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[53];
  assign _0840_ = _0839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58625" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[54];
  assign _0841_ = _0840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58626" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[55];
  assign _0842_ = _0841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58626" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[56];
  assign _0843_ = _0842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58627" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[57];
  assign _0844_ = _0843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58627" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[58];
  assign _0845_ = _0844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58628" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[59];
  assign _0846_ = _0845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58628" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[60];
  assign _0847_ = _0846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58629" *) IntShiftRight_49U_6U_32U_mbits_fixed_7_sva[61];
  assign _0848_ = _0847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58629" *) _0324_;
  assign _0849_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58634" *) _0325_;
  assign _0850_ = IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58639" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[1];
  assign _0851_ = _0850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58639" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[2];
  assign _0852_ = _0851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58640" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[3];
  assign _0853_ = _0852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58640" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[4];
  assign _0854_ = _0853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58641" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[5];
  assign _0855_ = _0854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58641" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[6];
  assign _0856_ = _0855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58642" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[7];
  assign _0857_ = _0856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58642" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[8];
  assign _0858_ = _0857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58643" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[9];
  assign _0859_ = _0858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58643" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[10];
  assign _0860_ = _0859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58644" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[11];
  assign _0861_ = _0860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58644" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[12];
  assign _0862_ = _0861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58645" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[13];
  assign _0863_ = _0862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58645" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[14];
  assign _0864_ = _0863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58646" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[15];
  assign _0865_ = _0864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58646" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[16];
  assign _0866_ = _0865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58647" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[17];
  assign _0867_ = _0866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58647" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[18];
  assign _0868_ = _0867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58648" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[19];
  assign _0869_ = _0868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58648" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[20];
  assign _0870_ = _0869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58649" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[21];
  assign _0871_ = _0870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58649" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[22];
  assign _0872_ = _0871_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58650" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[23];
  assign _0873_ = _0872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58650" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[24];
  assign _0874_ = _0873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58651" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[25];
  assign _0875_ = _0874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58651" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[26];
  assign _0876_ = _0875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58652" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[27];
  assign _0877_ = _0876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58652" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[28];
  assign _0878_ = _0877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58653" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[29];
  assign _0879_ = _0878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58653" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[30];
  assign _0880_ = _0879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58654" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[31];
  assign _0881_ = _0880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58654" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[32];
  assign _0882_ = _0881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58655" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[33];
  assign _0883_ = _0882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58655" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[34];
  assign _0884_ = _0883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58656" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[35];
  assign _0885_ = _0884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58656" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[36];
  assign _0886_ = _0885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58657" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[37];
  assign _0887_ = _0886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58657" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[38];
  assign _0888_ = _0887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58658" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[39];
  assign _0889_ = _0888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58658" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[40];
  assign _0890_ = _0889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58659" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[41];
  assign _0891_ = _0890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58659" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[42];
  assign _0892_ = _0891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58660" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[43];
  assign _0893_ = _0892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58660" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[44];
  assign _0894_ = _0893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58661" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[45];
  assign _0895_ = _0894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58661" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[46];
  assign _0896_ = _0895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58662" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[47];
  assign _0897_ = _0896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58662" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[48];
  assign _0898_ = _0897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58663" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[49];
  assign _0899_ = _0898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58663" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[50];
  assign _0900_ = _0899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58664" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[51];
  assign _0901_ = _0900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58664" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[52];
  assign _0902_ = _0901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58665" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[53];
  assign _0903_ = _0902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58665" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[54];
  assign _0904_ = _0903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58666" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[55];
  assign _0905_ = _0904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58666" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[56];
  assign _0906_ = _0905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58667" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[57];
  assign _0907_ = _0906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58667" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[58];
  assign _0908_ = _0907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58668" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[59];
  assign _0909_ = _0908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58668" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[60];
  assign _0910_ = _0909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58669" *) IntShiftRight_49U_6U_32U_mbits_fixed_8_sva[61];
  assign _0911_ = _0910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58669" *) _0327_;
  assign _0912_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58674" *) _0328_;
  assign _0913_ = IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58679" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[1];
  assign _0914_ = _0913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58679" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[2];
  assign _0915_ = _0914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58680" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[3];
  assign _0916_ = _0915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58680" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[4];
  assign _0917_ = _0916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58681" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[5];
  assign _0918_ = _0917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58681" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[6];
  assign _0919_ = _0918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58682" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[7];
  assign _0920_ = _0919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58682" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[8];
  assign _0921_ = _0920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58683" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[9];
  assign _0922_ = _0921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58683" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[10];
  assign _0923_ = _0922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58684" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[11];
  assign _0924_ = _0923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58684" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[12];
  assign _0925_ = _0924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58685" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[13];
  assign _0926_ = _0925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58685" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[14];
  assign _0927_ = _0926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58686" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[15];
  assign _0928_ = _0927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58686" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[16];
  assign _0929_ = _0928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58687" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[17];
  assign _0930_ = _0929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58687" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[18];
  assign _0931_ = _0930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58688" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[19];
  assign _0932_ = _0931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58688" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[20];
  assign _0933_ = _0932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58689" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[21];
  assign _0934_ = _0933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58689" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[22];
  assign _0935_ = _0934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58690" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[23];
  assign _0936_ = _0935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58690" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[24];
  assign _0937_ = _0936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58691" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[25];
  assign _0938_ = _0937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58691" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[26];
  assign _0939_ = _0938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58692" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[27];
  assign _0940_ = _0939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58692" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[28];
  assign _0941_ = _0940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58693" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[29];
  assign _0942_ = _0941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58693" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[30];
  assign _0943_ = _0942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58694" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[31];
  assign _0944_ = _0943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58694" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[32];
  assign _0945_ = _0944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58695" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[33];
  assign _0946_ = _0945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58695" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[34];
  assign _0947_ = _0946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58696" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[35];
  assign _0948_ = _0947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58696" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[36];
  assign _0949_ = _0948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58697" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[37];
  assign _0950_ = _0949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58697" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[38];
  assign _0951_ = _0950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58698" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[39];
  assign _0952_ = _0951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58698" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[40];
  assign _0953_ = _0952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58699" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[41];
  assign _0954_ = _0953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58699" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[42];
  assign _0955_ = _0954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58700" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[43];
  assign _0956_ = _0955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58700" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[44];
  assign _0957_ = _0956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58701" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[45];
  assign _0958_ = _0957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58701" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[46];
  assign _0959_ = _0958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58702" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[47];
  assign _0960_ = _0959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58702" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[48];
  assign _0961_ = _0960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58703" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[49];
  assign _0962_ = _0961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58703" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[50];
  assign _0963_ = _0962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58704" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[51];
  assign _0964_ = _0963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58704" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[52];
  assign _0965_ = _0964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58705" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[53];
  assign _0966_ = _0965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58705" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[54];
  assign _0967_ = _0966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58706" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[55];
  assign _0968_ = _0967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58706" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[56];
  assign _0969_ = _0968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58707" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[57];
  assign _0970_ = _0969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58707" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[58];
  assign _0971_ = _0970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58708" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[59];
  assign _0972_ = _0971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58708" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[60];
  assign _0973_ = _0972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58709" *) IntShiftRight_49U_6U_32U_mbits_fixed_9_sva[61];
  assign _0974_ = _0973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58709" *) _0330_;
  assign _0975_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58714" *) _0331_;
  assign _0976_ = IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58719" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[1];
  assign _0977_ = _0976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58719" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[2];
  assign _0978_ = _0977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58720" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[3];
  assign _0979_ = _0978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58720" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[4];
  assign _0980_ = _0979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58721" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[5];
  assign _0981_ = _0980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58721" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[6];
  assign _0982_ = _0981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58722" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[7];
  assign _0983_ = _0982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58722" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[8];
  assign _0984_ = _0983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58723" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[9];
  assign _0985_ = _0984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58723" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[10];
  assign _0986_ = _0985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58724" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[11];
  assign _0987_ = _0986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58724" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[12];
  assign _0988_ = _0987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58725" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[13];
  assign _0989_ = _0988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58725" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[14];
  assign _0990_ = _0989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58726" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[15];
  assign _0991_ = _0990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58726" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[16];
  assign _0992_ = _0991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58727" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[17];
  assign _0993_ = _0992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58727" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[18];
  assign _0994_ = _0993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58728" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[19];
  assign _0995_ = _0994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58728" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[20];
  assign _0996_ = _0995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58729" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[21];
  assign _0997_ = _0996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58729" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[22];
  assign _0998_ = _0997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58730" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[23];
  assign _0999_ = _0998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58730" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[24];
  assign _1000_ = _0999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58731" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[25];
  assign _1001_ = _1000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58731" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[26];
  assign _1002_ = _1001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58732" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[27];
  assign _1003_ = _1002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58732" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[28];
  assign _1004_ = _1003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58733" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[29];
  assign _1005_ = _1004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58733" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[30];
  assign _1006_ = _1005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58734" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[31];
  assign _1007_ = _1006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58734" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[32];
  assign _1008_ = _1007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58735" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[33];
  assign _1009_ = _1008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58735" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[34];
  assign _1010_ = _1009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58736" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[35];
  assign _1011_ = _1010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58736" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[36];
  assign _1012_ = _1011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58737" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[37];
  assign _1013_ = _1012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58737" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[38];
  assign _1014_ = _1013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58738" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[39];
  assign _1015_ = _1014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58738" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[40];
  assign _1016_ = _1015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58739" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[41];
  assign _1017_ = _1016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58739" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[42];
  assign _1018_ = _1017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58740" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[43];
  assign _1019_ = _1018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58740" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[44];
  assign _1020_ = _1019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58741" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[45];
  assign _1021_ = _1020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58741" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[46];
  assign _1022_ = _1021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58742" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[47];
  assign _1023_ = _1022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58742" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[48];
  assign _1024_ = _1023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58743" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[49];
  assign _1025_ = _1024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58743" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[50];
  assign _1026_ = _1025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58744" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[51];
  assign _1027_ = _1026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58744" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[52];
  assign _1028_ = _1027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58745" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[53];
  assign _1029_ = _1028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58745" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[54];
  assign _1030_ = _1029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58746" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[55];
  assign _1031_ = _1030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58746" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[56];
  assign _1032_ = _1031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58747" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[57];
  assign _1033_ = _1032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58747" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[58];
  assign _1034_ = _1033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58748" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[59];
  assign _1035_ = _1034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58748" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[60];
  assign _1036_ = _1035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58749" *) IntShiftRight_49U_6U_32U_mbits_fixed_10_sva[61];
  assign _1037_ = _1036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58749" *) _0333_;
  assign _1038_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58754" *) _0334_;
  assign _1039_ = IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58759" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[1];
  assign _1040_ = _1039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58759" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[2];
  assign _1041_ = _1040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58760" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[3];
  assign _1042_ = _1041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58760" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[4];
  assign _1043_ = _1042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58761" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[5];
  assign _1044_ = _1043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58761" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[6];
  assign _1045_ = _1044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58762" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[7];
  assign _1046_ = _1045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58762" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[8];
  assign _1047_ = _1046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58763" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[9];
  assign _1048_ = _1047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58763" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[10];
  assign _1049_ = _1048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58764" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[11];
  assign _1050_ = _1049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58764" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[12];
  assign _1051_ = _1050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58765" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[13];
  assign _1052_ = _1051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58765" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[14];
  assign _1053_ = _1052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58766" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[15];
  assign _1054_ = _1053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58766" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[16];
  assign _1055_ = _1054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58767" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[17];
  assign _1056_ = _1055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58767" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[18];
  assign _1057_ = _1056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58768" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[19];
  assign _1058_ = _1057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58768" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[20];
  assign _1059_ = _1058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58769" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[21];
  assign _1060_ = _1059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58769" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[22];
  assign _1061_ = _1060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58770" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[23];
  assign _1062_ = _1061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58770" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[24];
  assign _1063_ = _1062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58771" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[25];
  assign _1064_ = _1063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58771" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[26];
  assign _1065_ = _1064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58772" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[27];
  assign _1066_ = _1065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58772" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[28];
  assign _1067_ = _1066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58773" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[29];
  assign _1068_ = _1067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58773" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[30];
  assign _1069_ = _1068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58774" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[31];
  assign _1070_ = _1069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58774" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[32];
  assign _1071_ = _1070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58775" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[33];
  assign _1072_ = _1071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58775" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[34];
  assign _1073_ = _1072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58776" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[35];
  assign _1074_ = _1073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58776" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[36];
  assign _1075_ = _1074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58777" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[37];
  assign _1076_ = _1075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58777" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[38];
  assign _1077_ = _1076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58778" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[39];
  assign _1078_ = _1077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58778" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[40];
  assign _1079_ = _1078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58779" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[41];
  assign _1080_ = _1079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58779" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[42];
  assign _1081_ = _1080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58780" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[43];
  assign _1082_ = _1081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58780" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[44];
  assign _1083_ = _1082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58781" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[45];
  assign _1084_ = _1083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58781" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[46];
  assign _1085_ = _1084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58782" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[47];
  assign _1086_ = _1085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58782" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[48];
  assign _1087_ = _1086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58783" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[49];
  assign _1088_ = _1087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58783" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[50];
  assign _1089_ = _1088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58784" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[51];
  assign _1090_ = _1089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58784" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[52];
  assign _1091_ = _1090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58785" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[53];
  assign _1092_ = _1091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58785" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[54];
  assign _1093_ = _1092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58786" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[55];
  assign _1094_ = _1093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58786" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[56];
  assign _1095_ = _1094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58787" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[57];
  assign _1096_ = _1095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58787" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[58];
  assign _1097_ = _1096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58788" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[59];
  assign _1098_ = _1097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58788" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[60];
  assign _1099_ = _1098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58789" *) IntShiftRight_49U_6U_32U_mbits_fixed_11_sva[61];
  assign _1100_ = _1099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58789" *) _0336_;
  assign _1101_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58794" *) _0337_;
  assign _1102_ = IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58799" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[1];
  assign _1103_ = _1102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58799" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[2];
  assign _1104_ = _1103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58800" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[3];
  assign _1105_ = _1104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58800" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[4];
  assign _1106_ = _1105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58801" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[5];
  assign _1107_ = _1106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58801" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[6];
  assign _1108_ = _1107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58802" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[7];
  assign _1109_ = _1108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58802" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[8];
  assign _1110_ = _1109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58803" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[9];
  assign _1111_ = _1110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58803" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[10];
  assign _1112_ = _1111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58804" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[11];
  assign _1113_ = _1112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58804" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[12];
  assign _1114_ = _1113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58805" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[13];
  assign _1115_ = _1114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58805" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[14];
  assign _1116_ = _1115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58806" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[15];
  assign _1117_ = _1116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58806" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[16];
  assign _1118_ = _1117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58807" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[17];
  assign _1119_ = _1118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58807" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[18];
  assign _1120_ = _1119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58808" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[19];
  assign _1121_ = _1120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58808" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[20];
  assign _1122_ = _1121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58809" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[21];
  assign _1123_ = _1122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58809" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[22];
  assign _1124_ = _1123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58810" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[23];
  assign _1125_ = _1124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58810" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[24];
  assign _1126_ = _1125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58811" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[25];
  assign _1127_ = _1126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58811" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[26];
  assign _1128_ = _1127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58812" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[27];
  assign _1129_ = _1128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58812" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[28];
  assign _1130_ = _1129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58813" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[29];
  assign _1131_ = _1130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58813" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[30];
  assign _1132_ = _1131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58814" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[31];
  assign _1133_ = _1132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58814" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[32];
  assign _1134_ = _1133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58815" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[33];
  assign _1135_ = _1134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58815" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[34];
  assign _1136_ = _1135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58816" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[35];
  assign _1137_ = _1136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58816" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[36];
  assign _1138_ = _1137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58817" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[37];
  assign _1139_ = _1138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58817" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[38];
  assign _1140_ = _1139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58818" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[39];
  assign _1141_ = _1140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58818" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[40];
  assign _1142_ = _1141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58819" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[41];
  assign _1143_ = _1142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58819" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[42];
  assign _1144_ = _1143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58820" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[43];
  assign _1145_ = _1144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58820" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[44];
  assign _1146_ = _1145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58821" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[45];
  assign _1147_ = _1146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58821" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[46];
  assign _1148_ = _1147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58822" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[47];
  assign _1149_ = _1148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58822" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[48];
  assign _1150_ = _1149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58823" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[49];
  assign _1151_ = _1150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58823" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[50];
  assign _1152_ = _1151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58824" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[51];
  assign _1153_ = _1152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58824" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[52];
  assign _1154_ = _1153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58825" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[53];
  assign _1155_ = _1154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58825" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[54];
  assign _1156_ = _1155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58826" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[55];
  assign _1157_ = _1156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58826" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[56];
  assign _1158_ = _1157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58827" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[57];
  assign _1159_ = _1158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58827" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[58];
  assign _1160_ = _1159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58828" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[59];
  assign _1161_ = _1160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58828" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[60];
  assign _1162_ = _1161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58829" *) IntShiftRight_49U_6U_32U_mbits_fixed_12_sva[61];
  assign _1163_ = _1162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58829" *) _0339_;
  assign _1164_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58834" *) _0340_;
  assign _1165_ = IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58839" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[1];
  assign _1166_ = _1165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58839" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[2];
  assign _1167_ = _1166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58840" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[3];
  assign _1168_ = _1167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58840" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[4];
  assign _1169_ = _1168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58841" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[5];
  assign _1170_ = _1169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58841" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[6];
  assign _1171_ = _1170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58842" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[7];
  assign _1172_ = _1171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58842" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[8];
  assign _1173_ = _1172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58843" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[9];
  assign _1174_ = _1173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58843" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[10];
  assign _1175_ = _1174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58844" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[11];
  assign _1176_ = _1175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58844" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[12];
  assign _1177_ = _1176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58845" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[13];
  assign _1178_ = _1177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58845" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[14];
  assign _1179_ = _1178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58846" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[15];
  assign _1180_ = _1179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58846" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[16];
  assign _1181_ = _1180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58847" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[17];
  assign _1182_ = _1181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58847" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[18];
  assign _1183_ = _1182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58848" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[19];
  assign _1184_ = _1183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58848" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[20];
  assign _1185_ = _1184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58849" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[21];
  assign _1186_ = _1185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58849" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[22];
  assign _1187_ = _1186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58850" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[23];
  assign _1188_ = _1187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58850" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[24];
  assign _1189_ = _1188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58851" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[25];
  assign _1190_ = _1189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58851" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[26];
  assign _1191_ = _1190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58852" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[27];
  assign _1192_ = _1191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58852" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[28];
  assign _1193_ = _1192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58853" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[29];
  assign _1194_ = _1193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58853" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[30];
  assign _1195_ = _1194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58854" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[31];
  assign _1196_ = _1195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58854" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[32];
  assign _1197_ = _1196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58855" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[33];
  assign _1198_ = _1197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58855" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[34];
  assign _1199_ = _1198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58856" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[35];
  assign _1200_ = _1199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58856" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[36];
  assign _1201_ = _1200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58857" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[37];
  assign _1202_ = _1201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58857" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[38];
  assign _1203_ = _1202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58858" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[39];
  assign _1204_ = _1203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58858" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[40];
  assign _1205_ = _1204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58859" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[41];
  assign _1206_ = _1205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58859" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[42];
  assign _1207_ = _1206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58860" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[43];
  assign _1208_ = _1207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58860" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[44];
  assign _1209_ = _1208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58861" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[45];
  assign _1210_ = _1209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58861" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[46];
  assign _1211_ = _1210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58862" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[47];
  assign _1212_ = _1211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58862" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[48];
  assign _1213_ = _1212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58863" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[49];
  assign _1214_ = _1213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58863" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[50];
  assign _1215_ = _1214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58864" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[51];
  assign _1216_ = _1215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58864" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[52];
  assign _1217_ = _1216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58865" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[53];
  assign _1218_ = _1217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58865" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[54];
  assign _1219_ = _1218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58866" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[55];
  assign _1220_ = _1219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58866" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[56];
  assign _1221_ = _1220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58867" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[57];
  assign _1222_ = _1221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58867" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[58];
  assign _1223_ = _1222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58868" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[59];
  assign _1224_ = _1223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58868" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[60];
  assign _1225_ = _1224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58869" *) IntShiftRight_49U_6U_32U_mbits_fixed_13_sva[61];
  assign _1226_ = _1225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58869" *) _0342_;
  assign _1227_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58874" *) _0343_;
  assign _1228_ = IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58879" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[1];
  assign _1229_ = _1228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58879" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[2];
  assign _1230_ = _1229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58880" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[3];
  assign _1231_ = _1230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58880" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[4];
  assign _1232_ = _1231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58881" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[5];
  assign _1233_ = _1232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58881" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[6];
  assign _1234_ = _1233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58882" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[7];
  assign _1235_ = _1234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58882" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[8];
  assign _1236_ = _1235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58883" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[9];
  assign _1237_ = _1236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58883" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[10];
  assign _1238_ = _1237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58884" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[11];
  assign _1239_ = _1238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58884" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[12];
  assign _1240_ = _1239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58885" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[13];
  assign _1241_ = _1240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58885" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[14];
  assign _1242_ = _1241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58886" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[15];
  assign _1243_ = _1242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58886" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[16];
  assign _1244_ = _1243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58887" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[17];
  assign _1245_ = _1244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58887" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[18];
  assign _1246_ = _1245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58888" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[19];
  assign _1247_ = _1246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58888" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[20];
  assign _1248_ = _1247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58889" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[21];
  assign _1249_ = _1248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58889" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[22];
  assign _1250_ = _1249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58890" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[23];
  assign _1251_ = _1250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58890" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[24];
  assign _1252_ = _1251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58891" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[25];
  assign _1253_ = _1252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58891" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[26];
  assign _1254_ = _1253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58892" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[27];
  assign _1255_ = _1254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58892" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[28];
  assign _1256_ = _1255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58893" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[29];
  assign _1257_ = _1256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58893" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[30];
  assign _1258_ = _1257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58894" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[31];
  assign _1259_ = _1258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58894" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[32];
  assign _1260_ = _1259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58895" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[33];
  assign _1261_ = _1260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58895" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[34];
  assign _1262_ = _1261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58896" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[35];
  assign _1263_ = _1262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58896" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[36];
  assign _1264_ = _1263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58897" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[37];
  assign _1265_ = _1264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58897" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[38];
  assign _1266_ = _1265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58898" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[39];
  assign _1267_ = _1266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58898" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[40];
  assign _1268_ = _1267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58899" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[41];
  assign _1269_ = _1268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58899" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[42];
  assign _1270_ = _1269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58900" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[43];
  assign _1271_ = _1270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58900" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[44];
  assign _1272_ = _1271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58901" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[45];
  assign _1273_ = _1272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58901" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[46];
  assign _1274_ = _1273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58902" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[47];
  assign _1275_ = _1274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58902" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[48];
  assign _1276_ = _1275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58903" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[49];
  assign _1277_ = _1276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58903" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[50];
  assign _1278_ = _1277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58904" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[51];
  assign _1279_ = _1278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58904" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[52];
  assign _1280_ = _1279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58905" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[53];
  assign _1281_ = _1280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58905" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[54];
  assign _1282_ = _1281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58906" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[55];
  assign _1283_ = _1282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58906" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[56];
  assign _1284_ = _1283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58907" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[57];
  assign _1285_ = _1284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58907" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[58];
  assign _1286_ = _1285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58908" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[59];
  assign _1287_ = _1286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58908" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[60];
  assign _1288_ = _1287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58909" *) IntShiftRight_49U_6U_32U_mbits_fixed_14_sva[61];
  assign _1289_ = _1288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58909" *) _0345_;
  assign _1290_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58914" *) _0346_;
  assign _1291_ = IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58919" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[1];
  assign _1292_ = _1291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58919" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[2];
  assign _1293_ = _1292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58920" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[3];
  assign _1294_ = _1293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58920" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[4];
  assign _1295_ = _1294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58921" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[5];
  assign _1296_ = _1295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58921" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[6];
  assign _1297_ = _1296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58922" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[7];
  assign _1298_ = _1297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58922" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[8];
  assign _1299_ = _1298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58923" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[9];
  assign _1300_ = _1299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58923" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[10];
  assign _1301_ = _1300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58924" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[11];
  assign _1302_ = _1301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58924" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[12];
  assign _1303_ = _1302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58925" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[13];
  assign _1304_ = _1303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58925" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[14];
  assign _1305_ = _1304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58926" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[15];
  assign _1306_ = _1305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58926" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[16];
  assign _1307_ = _1306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58927" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[17];
  assign _1308_ = _1307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58927" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[18];
  assign _1309_ = _1308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58928" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[19];
  assign _1310_ = _1309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58928" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[20];
  assign _1311_ = _1310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58929" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[21];
  assign _1312_ = _1311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58929" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[22];
  assign _1313_ = _1312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58930" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[23];
  assign _1314_ = _1313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58930" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[24];
  assign _1315_ = _1314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58931" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[25];
  assign _1316_ = _1315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58931" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[26];
  assign _1317_ = _1316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58932" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[27];
  assign _1318_ = _1317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58932" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[28];
  assign _1319_ = _1318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58933" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[29];
  assign _1320_ = _1319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58933" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[30];
  assign _1321_ = _1320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58934" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[31];
  assign _1322_ = _1321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58934" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[32];
  assign _1323_ = _1322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58935" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[33];
  assign _1324_ = _1323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58935" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[34];
  assign _1325_ = _1324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58936" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[35];
  assign _1326_ = _1325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58936" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[36];
  assign _1327_ = _1326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58937" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[37];
  assign _1328_ = _1327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58937" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[38];
  assign _1329_ = _1328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58938" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[39];
  assign _1330_ = _1329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58938" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[40];
  assign _1331_ = _1330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58939" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[41];
  assign _1332_ = _1331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58939" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[42];
  assign _1333_ = _1332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58940" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[43];
  assign _1334_ = _1333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58940" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[44];
  assign _1335_ = _1334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58941" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[45];
  assign _1336_ = _1335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58941" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[46];
  assign _1337_ = _1336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58942" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[47];
  assign _1338_ = _1337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58942" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[48];
  assign _1339_ = _1338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58943" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[49];
  assign _1340_ = _1339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58943" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[50];
  assign _1341_ = _1340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58944" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[51];
  assign _1342_ = _1341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58944" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[52];
  assign _1343_ = _1342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58945" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[53];
  assign _1344_ = _1343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58945" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[54];
  assign _1345_ = _1344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58946" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[55];
  assign _1346_ = _1345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58946" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[56];
  assign _1347_ = _1346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58947" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[57];
  assign _1348_ = _1347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58947" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[58];
  assign _1349_ = _1348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58948" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[59];
  assign _1350_ = _1349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58948" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[60];
  assign _1351_ = _1350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58949" *) IntShiftRight_49U_6U_32U_mbits_fixed_15_sva[61];
  assign _1352_ = _1351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58949" *) _0348_;
  assign _1353_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58954" *) _0349_;
  assign _1354_ = IntShiftRight_49U_6U_32U_mbits_fixed_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58959" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[1];
  assign _1355_ = _1354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58959" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[2];
  assign _1356_ = _1355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58960" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[3];
  assign _1357_ = _1356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58960" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[4];
  assign _1358_ = _1357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58961" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[5];
  assign _1359_ = _1358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58961" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[6];
  assign _1360_ = _1359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58962" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[7];
  assign _1361_ = _1360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58962" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[8];
  assign _1362_ = _1361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58963" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[9];
  assign _1363_ = _1362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58963" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[10];
  assign _1364_ = _1363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58964" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[11];
  assign _1365_ = _1364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58964" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[12];
  assign _1366_ = _1365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58965" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[13];
  assign _1367_ = _1366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58965" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[14];
  assign _1368_ = _1367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58966" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[15];
  assign _1369_ = _1368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58966" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[16];
  assign _1370_ = _1369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58967" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[17];
  assign _1371_ = _1370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58967" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[18];
  assign _1372_ = _1371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58968" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[19];
  assign _1373_ = _1372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58968" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[20];
  assign _1374_ = _1373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58969" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[21];
  assign _1375_ = _1374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58969" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[22];
  assign _1376_ = _1375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58970" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[23];
  assign _1377_ = _1376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58970" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[24];
  assign _1378_ = _1377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58971" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[25];
  assign _1379_ = _1378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58971" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[26];
  assign _1380_ = _1379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58972" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[27];
  assign _1381_ = _1380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58972" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[28];
  assign _1382_ = _1381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58973" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[29];
  assign _1383_ = _1382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58973" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[30];
  assign _1384_ = _1383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58974" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[31];
  assign _1385_ = _1384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58974" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[32];
  assign _1386_ = _1385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58975" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[33];
  assign _1387_ = _1386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58975" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[34];
  assign _1388_ = _1387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58976" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[35];
  assign _1389_ = _1388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58976" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[36];
  assign _1390_ = _1389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58977" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[37];
  assign _1391_ = _1390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58977" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[38];
  assign _1392_ = _1391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58978" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[39];
  assign _1393_ = _1392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58978" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[40];
  assign _1394_ = _1393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58979" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[41];
  assign _1395_ = _1394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58979" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[42];
  assign _1396_ = _1395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58980" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[43];
  assign _1397_ = _1396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58980" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[44];
  assign _1398_ = _1397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58981" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[45];
  assign _1399_ = _1398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58981" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[46];
  assign _1400_ = _1399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58982" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[47];
  assign _1401_ = _1400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58982" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[48];
  assign _1402_ = _1401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58983" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[49];
  assign _1403_ = _1402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58983" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[50];
  assign _1404_ = _1403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58984" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[51];
  assign _1405_ = _1404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58984" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[52];
  assign _1406_ = _1405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58985" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[53];
  assign _1407_ = _1406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58985" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[54];
  assign _1408_ = _1407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58986" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[55];
  assign _1409_ = _1408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58986" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[56];
  assign _1410_ = _1409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58987" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[57];
  assign _1411_ = _1410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58987" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[58];
  assign _1412_ = _1411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58988" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[59];
  assign _1413_ = _1412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58988" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[60];
  assign _1414_ = _1413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58989" *) IntShiftRight_49U_6U_32U_mbits_fixed_sva[61];
  assign _1415_ = _1414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58989" *) _0351_;
  assign _1416_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58994" *) _0352_;
  assign _1417_ = chn_trt_out_rsci_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58997" *) _0354_;
  assign _1418_ = cfg_mul_shift_value_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58998" *) _0354_;
  assign or_dcpl = and_dcpl_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59000" *) _0354_;
  assign _1419_ = cfg_precision[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59008" *) _0355_;
  assign chn_trt_in_rsci_ld_core_psct_mx0c0 = and_4_mdf | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59016" *) fsm_output[0];
  assign chn_trt_out_rsci_d_0_mx0c1 = and_150_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59017" *) _0138_;
  assign _1420_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59020" *) chn_trt_in_rsci_d_mxwt[784];
  assign chn_trt_out_rsci_d_30_1_mx0c1 = _0140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59021" *) _0142_;
  assign _1421_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59024" *) chn_trt_in_rsci_d_mxwt[785];
  assign chn_trt_out_rsci_d_62_33_mx0c1 = _0144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59025" *) _0146_;
  assign _1422_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59028" *) chn_trt_in_rsci_d_mxwt[786];
  assign chn_trt_out_rsci_d_94_65_mx0c1 = _0148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59029" *) _0150_;
  assign _1423_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59032" *) chn_trt_in_rsci_d_mxwt[787];
  assign chn_trt_out_rsci_d_126_97_mx0c1 = _0152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59033" *) _0154_;
  assign _1424_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59036" *) chn_trt_in_rsci_d_mxwt[788];
  assign chn_trt_out_rsci_d_158_129_mx0c1 = _0156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59037" *) _0158_;
  assign _1425_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59040" *) chn_trt_in_rsci_d_mxwt[789];
  assign chn_trt_out_rsci_d_190_161_mx0c1 = _0160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59041" *) _0162_;
  assign _1426_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59044" *) chn_trt_in_rsci_d_mxwt[790];
  assign chn_trt_out_rsci_d_222_193_mx0c1 = _0164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59045" *) _0166_;
  assign _1427_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59048" *) chn_trt_in_rsci_d_mxwt[791];
  assign chn_trt_out_rsci_d_254_225_mx0c1 = _0168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59049" *) _0170_;
  assign _1428_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59052" *) chn_trt_in_rsci_d_mxwt[792];
  assign chn_trt_out_rsci_d_286_257_mx0c1 = _0172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59053" *) _0174_;
  assign _1429_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59056" *) chn_trt_in_rsci_d_mxwt[793];
  assign chn_trt_out_rsci_d_318_289_mx0c1 = _0176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59057" *) _0178_;
  assign _1430_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59060" *) chn_trt_in_rsci_d_mxwt[794];
  assign chn_trt_out_rsci_d_350_321_mx0c1 = _0180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59061" *) _0182_;
  assign _1431_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59064" *) chn_trt_in_rsci_d_mxwt[795];
  assign chn_trt_out_rsci_d_382_353_mx0c1 = _0184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59065" *) _0186_;
  assign _1432_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59068" *) chn_trt_in_rsci_d_mxwt[796];
  assign chn_trt_out_rsci_d_414_385_mx0c1 = _0188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59069" *) _0190_;
  assign _1433_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59072" *) chn_trt_in_rsci_d_mxwt[797];
  assign chn_trt_out_rsci_d_446_417_mx0c1 = _0192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59073" *) _0194_;
  assign _1434_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59076" *) chn_trt_in_rsci_d_mxwt[798];
  assign chn_trt_out_rsci_d_478_449_mx0c1 = _0196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59077" *) _0198_;
  assign _1435_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59080" *) chn_trt_in_rsci_d_mxwt[799];
  assign chn_trt_out_rsci_d_510_481_mx0c1 = _0200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59081" *) _0202_;
  assign _1436_ = and_148_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59106" *) _0205_;
  assign _1437_ = _1436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59106" *) chn_trt_out_rsci_d_0_mx0c1;
  assign _1438_ = _0209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59118" *) _0211_;
  assign _1439_ = _1438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59118" *) chn_trt_out_rsci_d_30_1_mx0c1;
  assign _1440_ = _0214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59228" *) _0215_;
  assign _1441_ = _1440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59228" *) chn_trt_out_rsci_d_62_33_mx0c1;
  assign _1442_ = _0218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59239" *) _0219_;
  assign _1443_ = _1442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59239" *) chn_trt_out_rsci_d_94_65_mx0c1;
  assign _1444_ = _0222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59250" *) _0223_;
  assign _1445_ = _1444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59250" *) chn_trt_out_rsci_d_126_97_mx0c1;
  assign _1446_ = _0226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59261" *) _0227_;
  assign _1447_ = _1446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59261" *) chn_trt_out_rsci_d_158_129_mx0c1;
  assign _1448_ = _0230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59272" *) _0231_;
  assign _1449_ = _1448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59272" *) chn_trt_out_rsci_d_190_161_mx0c1;
  assign _1450_ = _0234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59283" *) _0235_;
  assign _1451_ = _1450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59283" *) chn_trt_out_rsci_d_222_193_mx0c1;
  assign _1452_ = _0238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59294" *) _0239_;
  assign _1453_ = _1452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59294" *) chn_trt_out_rsci_d_254_225_mx0c1;
  assign _1454_ = _0242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59305" *) _0243_;
  assign _1455_ = _1454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59305" *) chn_trt_out_rsci_d_286_257_mx0c1;
  assign _1456_ = _0246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59316" *) _0247_;
  assign _1457_ = _1456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59316" *) chn_trt_out_rsci_d_318_289_mx0c1;
  assign _1458_ = _0250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59327" *) _0251_;
  assign _1459_ = _1458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59327" *) chn_trt_out_rsci_d_350_321_mx0c1;
  assign _1460_ = _0254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59338" *) _0255_;
  assign _1461_ = _1460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59338" *) chn_trt_out_rsci_d_382_353_mx0c1;
  assign _1462_ = _0258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59349" *) _0259_;
  assign _1463_ = _1462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59349" *) chn_trt_out_rsci_d_414_385_mx0c1;
  assign _1464_ = _0262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59360" *) _0263_;
  assign _1465_ = _1464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59360" *) chn_trt_out_rsci_d_446_417_mx0c1;
  assign _1466_ = _0266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59371" *) _0267_;
  assign _1467_ = _1466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59371" *) chn_trt_out_rsci_d_478_449_mx0c1;
  assign _1468_ = _0270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59382" *) _0271_;
  assign _1469_ = _1468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59382" *) chn_trt_out_rsci_d_510_481_mx0c1;
  assign _1470_ = or_tmp_150 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59391" *) and_dcpl_134;
  assign _1471_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59396" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva;
  assign _1472_ = _0376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59397" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva;
  assign _1473_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59406" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva;
  assign _1474_ = _0377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59407" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_1_sva;
  assign _1475_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59411" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva;
  assign _1476_ = _0378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59412" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva;
  assign _1477_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59416" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva;
  assign _1478_ = _0379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59417" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_2_sva;
  assign _1479_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59421" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva;
  assign _1480_ = _0380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59422" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva;
  assign _1481_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59426" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva;
  assign _1482_ = _0381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59427" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_3_sva;
  assign _1483_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59431" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva;
  assign _1484_ = _0382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59432" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva;
  assign _1485_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59436" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva;
  assign _1486_ = _0383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59437" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_4_sva;
  assign _1487_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59441" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva;
  assign _1488_ = _0384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59442" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva;
  assign _1489_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59446" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva;
  assign _1490_ = _0385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59447" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_5_sva;
  assign _1491_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59451" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva;
  assign _1492_ = _0386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59452" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva;
  assign _1493_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59456" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva;
  assign _1494_ = _0387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59457" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_6_sva;
  assign _1495_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59461" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva;
  assign _1496_ = _0388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59462" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva;
  assign _1497_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59466" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva;
  assign _1498_ = _0389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59467" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_7_sva;
  assign _1499_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59471" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva;
  assign _1500_ = _0390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59472" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva;
  assign _1501_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59476" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva;
  assign _1502_ = _0391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59477" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_8_sva;
  assign _1503_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59481" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva;
  assign _1504_ = _0392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59482" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva;
  assign _1505_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59486" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva;
  assign _1506_ = _0393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59487" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_9_sva;
  assign _1507_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59491" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva;
  assign _1508_ = _0394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59492" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva;
  assign _1509_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59496" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva;
  assign _1510_ = _0395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59497" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_10_sva;
  assign _1511_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59501" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva;
  assign _1512_ = _0396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59502" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva;
  assign _1513_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59506" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva;
  assign _1514_ = _0397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59507" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_11_sva;
  assign _1515_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59511" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva;
  assign _1516_ = _0398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59512" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva;
  assign _1517_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59516" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva;
  assign _1518_ = _0399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59517" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_12_sva;
  assign _1519_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59521" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva;
  assign _1520_ = _0400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59522" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva;
  assign _1521_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59526" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva;
  assign _1522_ = _0401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59527" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_13_sva;
  assign _1523_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59531" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva;
  assign _1524_ = _0402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59532" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva;
  assign _1525_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59536" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva;
  assign _1526_ = _0403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59537" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_14_sva;
  assign _1527_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59541" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva;
  assign _1528_ = _0404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59542" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva;
  assign _1529_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59546" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva;
  assign _1530_ = _0405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59547" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_15_sva;
  assign _1531_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59551" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva;
  assign _1532_ = _0406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59552" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva;
  assign _1533_ = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59556" *) IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva;
  assign _1534_ = _0407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59557" *) IntShiftRight_49U_6U_32U_obits_fixed_nor_ovfl_sva;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_trt_out_rsci_ld_core_psct_cse <= 1'b0;
    else
      reg_chn_trt_out_rsci_ld_core_psct_cse <= _0083_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_510_481 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_510_481 <= _0074_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_478_449 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_478_449 <= _0071_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_446_417 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_446_417 <= _0068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_414_385 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_414_385 <= _0065_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_382_353 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_382_353 <= _0062_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_350_321 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_350_321 <= _0059_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_318_289 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_318_289 <= _0054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_286_257 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_286_257 <= _0050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_254_225 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_254_225 <= _0047_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_222_193 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_222_193 <= _0044_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_190_161 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_190_161 <= _0041_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_158_129 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_158_129 <= _0038_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_126_97 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_126_97 <= _0035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_94_65 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_94_65 <= _0079_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_62_33 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_62_33 <= _0076_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_511 <= 1'b0;
    else
      chn_trt_out_rsci_d_511 <= _0075_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_480 <= 1'b0;
    else
      chn_trt_out_rsci_d_480 <= _0073_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_479 <= 1'b0;
    else
      chn_trt_out_rsci_d_479 <= _0072_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_448 <= 1'b0;
    else
      chn_trt_out_rsci_d_448 <= _0070_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_447 <= 1'b0;
    else
      chn_trt_out_rsci_d_447 <= _0069_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_416 <= 1'b0;
    else
      chn_trt_out_rsci_d_416 <= _0067_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_415 <= 1'b0;
    else
      chn_trt_out_rsci_d_415 <= _0066_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_384 <= 1'b0;
    else
      chn_trt_out_rsci_d_384 <= _0064_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_383 <= 1'b0;
    else
      chn_trt_out_rsci_d_383 <= _0063_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_352 <= 1'b0;
    else
      chn_trt_out_rsci_d_352 <= _0061_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_351 <= 1'b0;
    else
      chn_trt_out_rsci_d_351 <= _0060_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_320 <= 1'b0;
    else
      chn_trt_out_rsci_d_320 <= _0057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_319 <= 1'b0;
    else
      chn_trt_out_rsci_d_319 <= _0055_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_288 <= 1'b0;
    else
      chn_trt_out_rsci_d_288 <= _0052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_287 <= 1'b0;
    else
      chn_trt_out_rsci_d_287 <= _0051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_256 <= 1'b0;
    else
      chn_trt_out_rsci_d_256 <= _0049_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_255 <= 1'b0;
    else
      chn_trt_out_rsci_d_255 <= _0048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_224 <= 1'b0;
    else
      chn_trt_out_rsci_d_224 <= _0046_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_223 <= 1'b0;
    else
      chn_trt_out_rsci_d_223 <= _0045_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_192 <= 1'b0;
    else
      chn_trt_out_rsci_d_192 <= _0043_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_191 <= 1'b0;
    else
      chn_trt_out_rsci_d_191 <= _0042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_160 <= 1'b0;
    else
      chn_trt_out_rsci_d_160 <= _0040_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_159 <= 1'b0;
    else
      chn_trt_out_rsci_d_159 <= _0039_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_128 <= 1'b0;
    else
      chn_trt_out_rsci_d_128 <= _0037_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_127 <= 1'b0;
    else
      chn_trt_out_rsci_d_127 <= _0036_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_96 <= 1'b0;
    else
      chn_trt_out_rsci_d_96 <= _0081_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_95 <= 1'b0;
    else
      chn_trt_out_rsci_d_95 <= _0080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_64 <= 1'b0;
    else
      chn_trt_out_rsci_d_64 <= _0078_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_63 <= 1'b0;
    else
      chn_trt_out_rsci_d_63 <= _0077_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_32 <= 1'b0;
    else
      chn_trt_out_rsci_d_32 <= _0058_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_31 <= 1'b0;
    else
      chn_trt_out_rsci_d_31 <= _0056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_30_1 <= 30'b000000000000000000000000000000;
    else
      chn_trt_out_rsci_d_30_1 <= _0053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_out_rsci_d_0 <= 1'b0;
    else
      chn_trt_out_rsci_d_0 <= _0034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_in_rsci_ld_core_psct <= 1'b0;
    else
      chn_trt_in_rsci_ld_core_psct <= _0033_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_trt_in_rsci_iswt0 <= 1'b0;
    else
      chn_trt_in_rsci_iswt0 <= _0032_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
    else
      reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse <= _0082_;
  assign _0031_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0030_ = _1416_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0029_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_15_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0028_ = _1353_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0027_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_14_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0026_ = _1290_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0025_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_13_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0024_ = _1227_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0023_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_12_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0022_ = _1164_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0021_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_11_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0020_ = _1101_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0019_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_10_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0018_ = _1038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0017_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_9_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0016_ = _0975_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0015_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_8_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0014_ = _0912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0013_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_7_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0012_ = _0849_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0011_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_6_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0010_ = _0786_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0009_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_5_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0008_ = _0723_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0007_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_4_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0006_ = _0660_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0005_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_3_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0004_ = _0597_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[30:1] : 30'b111111111111111111111111111111;
  assign _0003_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_2_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0002_ = _0534_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[30:1] : 30'b111111111111111111111111111111;
  assign trt_loop_else_mux_143_nl = chn_trt_in_rsci_d_mxwt[799] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[766] : trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_142_nl = chn_trt_in_rsci_d_mxwt[799] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[735] : trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_141_nl = chn_trt_in_rsci_d_mxwt[798] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[717] : trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_140_nl = chn_trt_in_rsci_d_mxwt[798] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[686] : trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_139_nl = chn_trt_in_rsci_d_mxwt[797] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[668] : trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_138_nl = chn_trt_in_rsci_d_mxwt[797] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[637] : trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_137_nl = chn_trt_in_rsci_d_mxwt[796] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[619] : trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_136_nl = chn_trt_in_rsci_d_mxwt[796] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[588] : trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_135_nl = chn_trt_in_rsci_d_mxwt[795] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[570] : trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_134_nl = chn_trt_in_rsci_d_mxwt[795] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[539] : trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_133_nl = chn_trt_in_rsci_d_mxwt[794] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[521] : trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_132_nl = chn_trt_in_rsci_d_mxwt[794] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[490] : trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_131_nl = chn_trt_in_rsci_d_mxwt[793] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[472] : trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_130_nl = chn_trt_in_rsci_d_mxwt[793] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[441] : trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_129_nl = chn_trt_in_rsci_d_mxwt[792] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[423] : trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_128_nl = chn_trt_in_rsci_d_mxwt[792] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[392] : trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_127_nl = chn_trt_in_rsci_d_mxwt[791] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[374] : trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_126_nl = chn_trt_in_rsci_d_mxwt[791] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[343] : trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_125_nl = chn_trt_in_rsci_d_mxwt[790] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[325] : trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_124_nl = chn_trt_in_rsci_d_mxwt[790] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[294] : trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_123_nl = chn_trt_in_rsci_d_mxwt[789] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[276] : trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_122_nl = chn_trt_in_rsci_d_mxwt[789] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[245] : trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_121_nl = chn_trt_in_rsci_d_mxwt[788] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[227] : trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_120_nl = chn_trt_in_rsci_d_mxwt[788] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[196] : trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_119_nl = chn_trt_in_rsci_d_mxwt[787] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[178] : trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_118_nl = chn_trt_in_rsci_d_mxwt[787] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[147] : trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_117_nl = chn_trt_in_rsci_d_mxwt[786] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[129] : trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_116_nl = chn_trt_in_rsci_d_mxwt[786] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[98] : trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_115_nl = chn_trt_in_rsci_d_mxwt[785] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[80] : trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign trt_loop_else_mux_114_nl = chn_trt_in_rsci_d_mxwt[785] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[49] : trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign trt_loop_else_mux_113_nl = chn_trt_in_rsci_d_mxwt[784] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[31] : trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0001_ = IntShiftRight_49U_6U_32U_obits_fixed_and_unfl_1_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) 30'b111111111111111111111111111111 : trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_nor_2_nl;
  assign _0000_ = _0471_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[30:1] : 30'b111111111111111111111111111111;
  assign trt_loop_else_mux_112_nl = chn_trt_in_rsci_d_mxwt[784] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[0] : trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_1_nl;
  assign mux_19_nl = chn_trt_in_rsci_d_mxwt[799] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_18_nl = chn_trt_in_rsci_d_mxwt[798] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_17_nl = chn_trt_in_rsci_d_mxwt[797] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_16_nl = chn_trt_in_rsci_d_mxwt[796] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_15_nl = chn_trt_in_rsci_d_mxwt[795] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_14_nl = chn_trt_in_rsci_d_mxwt[794] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_13_nl = chn_trt_in_rsci_d_mxwt[793] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_12_nl = chn_trt_in_rsci_d_mxwt[792] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_11_nl = chn_trt_in_rsci_d_mxwt[791] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_10_nl = chn_trt_in_rsci_d_mxwt[790] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_9_nl = chn_trt_in_rsci_d_mxwt[789] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_8_nl = chn_trt_in_rsci_d_mxwt[788] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_7_nl = chn_trt_in_rsci_d_mxwt[787] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_6_nl = chn_trt_in_rsci_d_mxwt[786] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_5_nl = chn_trt_in_rsci_d_mxwt[785] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign mux_4_nl = chn_trt_in_rsci_d_mxwt[784] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) or_dcpl : not_tmp_9;
  assign _0083_ = _0273_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59391" *) _0375_ : reg_chn_trt_out_rsci_ld_core_psct_cse;
  assign _0131_ = chn_trt_out_rsci_d_510_481_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[765:736] : trt_loop_16_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0074_ = _0272_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59382" *) _0131_ : chn_trt_out_rsci_d_510_481;
  assign _0130_ = chn_trt_out_rsci_d_478_449_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[716:687] : trt_loop_15_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0071_ = _0268_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59371" *) _0130_ : chn_trt_out_rsci_d_478_449;
  assign _0129_ = chn_trt_out_rsci_d_446_417_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[667:638] : trt_loop_14_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0068_ = _0264_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59360" *) _0129_ : chn_trt_out_rsci_d_446_417;
  assign _0128_ = chn_trt_out_rsci_d_414_385_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[618:589] : trt_loop_13_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0065_ = _0260_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59349" *) _0128_ : chn_trt_out_rsci_d_414_385;
  assign _0127_ = chn_trt_out_rsci_d_382_353_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[569:540] : trt_loop_12_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0062_ = _0256_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59338" *) _0127_ : chn_trt_out_rsci_d_382_353;
  assign _0126_ = chn_trt_out_rsci_d_350_321_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[520:491] : trt_loop_11_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0059_ = _0252_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59327" *) _0126_ : chn_trt_out_rsci_d_350_321;
  assign _0125_ = chn_trt_out_rsci_d_318_289_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[471:442] : trt_loop_10_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0054_ = _0248_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59316" *) _0125_ : chn_trt_out_rsci_d_318_289;
  assign _0124_ = chn_trt_out_rsci_d_286_257_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[422:393] : trt_loop_9_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0050_ = _0244_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59305" *) _0124_ : chn_trt_out_rsci_d_286_257;
  assign _0123_ = chn_trt_out_rsci_d_254_225_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[373:344] : trt_loop_8_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0047_ = _0240_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59294" *) _0123_ : chn_trt_out_rsci_d_254_225;
  assign _0122_ = chn_trt_out_rsci_d_222_193_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[324:295] : trt_loop_7_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0044_ = _0236_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59283" *) _0122_ : chn_trt_out_rsci_d_222_193;
  assign _0121_ = chn_trt_out_rsci_d_190_161_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[275:246] : trt_loop_6_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0041_ = _0232_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59272" *) _0121_ : chn_trt_out_rsci_d_190_161;
  assign _0120_ = chn_trt_out_rsci_d_158_129_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[226:197] : trt_loop_5_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0038_ = _0228_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59261" *) _0120_ : chn_trt_out_rsci_d_158_129;
  assign _0119_ = chn_trt_out_rsci_d_126_97_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[177:148] : trt_loop_4_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0035_ = _0224_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59250" *) _0119_ : chn_trt_out_rsci_d_126_97;
  assign _0118_ = chn_trt_out_rsci_d_94_65_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[128:99] : trt_loop_3_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0079_ = _0220_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59239" *) _0118_ : chn_trt_out_rsci_d_94_65;
  assign _0117_ = chn_trt_out_rsci_d_62_33_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[79:50] : trt_loop_2_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0076_ = _0216_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59228" *) _0117_ : chn_trt_out_rsci_d_62_33;
  assign _0115_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[766] : trt_loop_else_mux_143_nl;
  assign _0114_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[735] : trt_loop_else_mux_142_nl;
  assign _0113_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[717] : trt_loop_else_mux_141_nl;
  assign _0112_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[686] : trt_loop_else_mux_140_nl;
  assign _0111_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[668] : trt_loop_else_mux_139_nl;
  assign _0110_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[637] : trt_loop_else_mux_138_nl;
  assign _0109_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[619] : trt_loop_else_mux_137_nl;
  assign _0108_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[588] : trt_loop_else_mux_136_nl;
  assign _0107_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[570] : trt_loop_else_mux_135_nl;
  assign _0106_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[539] : trt_loop_else_mux_134_nl;
  assign _0105_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[521] : trt_loop_else_mux_133_nl;
  assign _0104_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[490] : trt_loop_else_mux_132_nl;
  assign _0103_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[472] : trt_loop_else_mux_131_nl;
  assign _0102_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[441] : trt_loop_else_mux_130_nl;
  assign _0101_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[423] : trt_loop_else_mux_129_nl;
  assign _0100_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[392] : trt_loop_else_mux_128_nl;
  assign _0099_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[374] : trt_loop_else_mux_127_nl;
  assign _0098_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[343] : trt_loop_else_mux_126_nl;
  assign _0097_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[325] : trt_loop_else_mux_125_nl;
  assign _0096_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[294] : trt_loop_else_mux_124_nl;
  assign _0095_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[276] : trt_loop_else_mux_123_nl;
  assign _0094_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[245] : trt_loop_else_mux_122_nl;
  assign _0093_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[227] : trt_loop_else_mux_121_nl;
  assign _0092_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[196] : trt_loop_else_mux_120_nl;
  assign _0091_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[178] : trt_loop_else_mux_119_nl;
  assign _0090_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[147] : trt_loop_else_mux_118_nl;
  assign _0089_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[129] : trt_loop_else_mux_117_nl;
  assign _0088_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[98] : trt_loop_else_mux_116_nl;
  assign _0087_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[80] : trt_loop_else_mux_115_nl;
  assign _0086_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[49] : trt_loop_else_mux_114_nl;
  assign _0085_ = and_150_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[31] : trt_loop_else_mux_113_nl;
  assign _0056_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0085_ : chn_trt_out_rsci_d_31;
  assign _0058_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0086_ : chn_trt_out_rsci_d_32;
  assign _0077_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0087_ : chn_trt_out_rsci_d_63;
  assign _0078_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0088_ : chn_trt_out_rsci_d_64;
  assign _0080_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0089_ : chn_trt_out_rsci_d_95;
  assign _0081_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0090_ : chn_trt_out_rsci_d_96;
  assign _0036_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0091_ : chn_trt_out_rsci_d_127;
  assign _0037_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0092_ : chn_trt_out_rsci_d_128;
  assign _0039_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0093_ : chn_trt_out_rsci_d_159;
  assign _0040_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0094_ : chn_trt_out_rsci_d_160;
  assign _0042_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0095_ : chn_trt_out_rsci_d_191;
  assign _0043_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0096_ : chn_trt_out_rsci_d_192;
  assign _0045_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0097_ : chn_trt_out_rsci_d_223;
  assign _0046_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0098_ : chn_trt_out_rsci_d_224;
  assign _0048_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0099_ : chn_trt_out_rsci_d_255;
  assign _0049_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0100_ : chn_trt_out_rsci_d_256;
  assign _0051_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0101_ : chn_trt_out_rsci_d_287;
  assign _0052_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0102_ : chn_trt_out_rsci_d_288;
  assign _0055_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0103_ : chn_trt_out_rsci_d_319;
  assign _0057_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0104_ : chn_trt_out_rsci_d_320;
  assign _0060_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0105_ : chn_trt_out_rsci_d_351;
  assign _0061_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0106_ : chn_trt_out_rsci_d_352;
  assign _0063_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0107_ : chn_trt_out_rsci_d_383;
  assign _0064_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0108_ : chn_trt_out_rsci_d_384;
  assign _0066_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0109_ : chn_trt_out_rsci_d_415;
  assign _0067_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0110_ : chn_trt_out_rsci_d_416;
  assign _0069_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0111_ : chn_trt_out_rsci_d_447;
  assign _0070_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0112_ : chn_trt_out_rsci_d_448;
  assign _0072_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0113_ : chn_trt_out_rsci_d_479;
  assign _0073_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0114_ : chn_trt_out_rsci_d_480;
  assign _0075_ = chn_trt_out_and_2_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59157" *) _0115_ : chn_trt_out_rsci_d_511;
  assign _0116_ = chn_trt_out_rsci_d_30_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59659|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59658" *) chn_trt_in_rsci_d_mxwt[30:1] : trt_loop_1_IntShiftRight_49U_6U_32U_obits_fixed_IntShiftRight_49U_6U_32U_obits_fixed_nor_nl;
  assign _0053_ = _0212_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59118" *) _0116_ : chn_trt_out_rsci_d_30_1;
  assign _0084_ = chn_trt_out_rsci_d_0_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59642|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59641" *) chn_trt_in_rsci_d_mxwt[0] : trt_loop_else_mux_112_nl;
  assign _0034_ = _0206_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59107" *) _0084_ : chn_trt_out_rsci_d_0;
  assign _0033_ = _0204_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59098" *) chn_trt_in_rsci_ld_core_psct_mx0c0 : chn_trt_in_rsci_ld_core_psct;
  assign _0082_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59089" *) or_tmp_150 : reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse;
  assign _0032_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:59089" *) _0358_ : chn_trt_in_rsci_iswt0;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58331" *)
  SDP_X_X_trt_core_cfg_mul_shift_value_rsc_triosy_obj X_trt_core_cfg_mul_shift_value_rsc_triosy_obj_inst (
    .cfg_mul_shift_value_rsc_triosy_lz(cfg_mul_shift_value_rsc_triosy_lz),
    .cfg_mul_shift_value_rsc_triosy_obj_bawt(cfg_mul_shift_value_rsc_triosy_obj_bawt),
    .cfg_mul_shift_value_rsc_triosy_obj_iswt0(reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_mul_shift_value_rsc_triosy_obj_oswt(cfg_mul_shift_value_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58299" *)
  SDP_X_X_trt_core_chn_trt_in_rsci X_trt_core_chn_trt_in_rsci_inst (
    .chn_trt_in_rsc_lz(chn_trt_in_rsc_lz),
    .chn_trt_in_rsc_slz(chn_trt_in_rsc_slz),
    .chn_trt_in_rsc_sz(chn_trt_in_rsc_sz),
    .chn_trt_in_rsc_vz(chn_trt_in_rsc_vz),
    .chn_trt_in_rsc_z(chn_trt_in_rsc_z),
    .chn_trt_in_rsci_bawt(chn_trt_in_rsci_bawt),
    .chn_trt_in_rsci_d_mxwt(chn_trt_in_rsci_d_mxwt),
    .chn_trt_in_rsci_iswt0(chn_trt_in_rsci_iswt0),
    .chn_trt_in_rsci_ld_core_psct(chn_trt_in_rsci_ld_core_psct),
    .chn_trt_in_rsci_oswt(chn_trt_in_rsci_oswt),
    .chn_trt_in_rsci_wen_comp(chn_trt_in_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58316" *)
  SDP_X_X_trt_core_chn_trt_out_rsci X_trt_core_chn_trt_out_rsci_inst (
    .chn_trt_out_rsc_lz(chn_trt_out_rsc_lz),
    .chn_trt_out_rsc_vz(chn_trt_out_rsc_vz),
    .chn_trt_out_rsc_z(chn_trt_out_rsc_z),
    .chn_trt_out_rsci_bawt(chn_trt_out_rsci_bawt),
    .chn_trt_out_rsci_d({ chn_trt_out_rsci_d_511, chn_trt_out_rsci_d_510_481, chn_trt_out_rsci_d_480, chn_trt_out_rsci_d_479, chn_trt_out_rsci_d_478_449, chn_trt_out_rsci_d_448, chn_trt_out_rsci_d_447, chn_trt_out_rsci_d_446_417, chn_trt_out_rsci_d_416, chn_trt_out_rsci_d_415, chn_trt_out_rsci_d_414_385, chn_trt_out_rsci_d_384, chn_trt_out_rsci_d_383, chn_trt_out_rsci_d_382_353, chn_trt_out_rsci_d_352, chn_trt_out_rsci_d_351, chn_trt_out_rsci_d_350_321, chn_trt_out_rsci_d_320, chn_trt_out_rsci_d_319, chn_trt_out_rsci_d_318_289, chn_trt_out_rsci_d_288, chn_trt_out_rsci_d_287, chn_trt_out_rsci_d_286_257, chn_trt_out_rsci_d_256, chn_trt_out_rsci_d_255, chn_trt_out_rsci_d_254_225, chn_trt_out_rsci_d_224, chn_trt_out_rsci_d_223, chn_trt_out_rsci_d_222_193, chn_trt_out_rsci_d_192, chn_trt_out_rsci_d_191, chn_trt_out_rsci_d_190_161, chn_trt_out_rsci_d_160, chn_trt_out_rsci_d_159, chn_trt_out_rsci_d_158_129, chn_trt_out_rsci_d_128, chn_trt_out_rsci_d_127, chn_trt_out_rsci_d_126_97, chn_trt_out_rsci_d_96, chn_trt_out_rsci_d_95, chn_trt_out_rsci_d_94_65, chn_trt_out_rsci_d_64, chn_trt_out_rsci_d_63, chn_trt_out_rsci_d_62_33, chn_trt_out_rsci_d_32, chn_trt_out_rsci_d_31, chn_trt_out_rsci_d_30_1, chn_trt_out_rsci_d_0 }),
    .chn_trt_out_rsci_iswt0(reg_cfg_mul_shift_value_rsc_triosy_obj_ld_core_psct_cse),
    .chn_trt_out_rsci_ld_core_psct(reg_chn_trt_out_rsci_ld_core_psct_cse),
    .chn_trt_out_rsci_oswt(chn_trt_out_rsci_oswt),
    .chn_trt_out_rsci_wen_comp(chn_trt_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58350" *)
  SDP_X_X_trt_core_core_fsm X_trt_core_core_fsm_inst (
    .core_wen(core_wen),
    .fsm_output(fsm_output),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58342" *)
  SDP_X_X_trt_core_staller X_trt_core_staller_inst (
    .chn_trt_in_rsci_wen_comp(chn_trt_in_rsci_wen_comp),
    .chn_trt_out_rsci_wen_comp(chn_trt_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58236" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_10_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[489:441], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_10_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58245" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_11_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[538:490], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_11_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58254" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_12_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[587:539], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_12_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58263" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_13_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[636:588], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_13_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58272" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_14_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[685:637], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_14_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58281" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_15_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[734:686], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_15_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58290" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_16_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[783:735], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58164" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_1_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[48:0], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58172" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_2_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[97:49], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58180" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_3_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[146:98], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58188" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_4_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[195:147], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_4_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58196" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_5_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[244:196], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_5_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58204" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_6_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[293:245], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_6_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58212" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_7_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[342:294], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_7_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58220" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_8_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[391:343], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_8_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:58228" *)
  \$paramod\SDP_X_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  trt_loop_9_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg (
    .a({ chn_trt_in_rsci_d_mxwt[440:392], 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_mul_shift_value_rsci_d),
    .z(IntShiftRight_49U_6U_32U_mbits_fixed_9_sva)
  );
  assign chn_trt_in_rsci_oswt_unreg = or_tmp_150;
  assign chn_trt_out_rsci_oswt_unreg_pff = and_dcpl_3;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_10_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_11_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_12_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_13_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_14_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_15_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_1_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_2_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_3_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_4_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_5_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_6_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_7_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_8_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_9_sva;
  assign nl_IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva[49:0] = IntShiftRight_49U_6U_32U_obits_fixed_acc_sat_sva;
  assign nl_X_trt_core_chn_trt_out_rsci_inst_chn_trt_out_rsci_d = { chn_trt_out_rsci_d_511, chn_trt_out_rsci_d_510_481, chn_trt_out_rsci_d_480, chn_trt_out_rsci_d_479, chn_trt_out_rsci_d_478_449, chn_trt_out_rsci_d_448, chn_trt_out_rsci_d_447, chn_trt_out_rsci_d_446_417, chn_trt_out_rsci_d_416, chn_trt_out_rsci_d_415, chn_trt_out_rsci_d_414_385, chn_trt_out_rsci_d_384, chn_trt_out_rsci_d_383, chn_trt_out_rsci_d_382_353, chn_trt_out_rsci_d_352, chn_trt_out_rsci_d_351, chn_trt_out_rsci_d_350_321, chn_trt_out_rsci_d_320, chn_trt_out_rsci_d_319, chn_trt_out_rsci_d_318_289, chn_trt_out_rsci_d_288, chn_trt_out_rsci_d_287, chn_trt_out_rsci_d_286_257, chn_trt_out_rsci_d_256, chn_trt_out_rsci_d_255, chn_trt_out_rsci_d_254_225, chn_trt_out_rsci_d_224, chn_trt_out_rsci_d_223, chn_trt_out_rsci_d_222_193, chn_trt_out_rsci_d_192, chn_trt_out_rsci_d_191, chn_trt_out_rsci_d_190_161, chn_trt_out_rsci_d_160, chn_trt_out_rsci_d_159, chn_trt_out_rsci_d_158_129, chn_trt_out_rsci_d_128, chn_trt_out_rsci_d_127, chn_trt_out_rsci_d_126_97, chn_trt_out_rsci_d_96, chn_trt_out_rsci_d_95, chn_trt_out_rsci_d_94_65, chn_trt_out_rsci_d_64, chn_trt_out_rsci_d_63, chn_trt_out_rsci_d_62_33, chn_trt_out_rsci_d_32, chn_trt_out_rsci_d_31, chn_trt_out_rsci_d_30_1, chn_trt_out_rsci_d_0 };
  assign nl_trt_loop_10_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[489:441], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_11_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[538:490], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_12_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[587:539], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_13_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[636:588], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_14_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[685:637], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_15_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[734:686], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_16_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[783:735], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_1_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[48:0], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_2_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[97:49], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_3_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[146:98], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_4_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[195:147], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_5_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[244:196], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_6_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[293:245], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_7_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[342:294], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_8_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[391:343], 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_trt_loop_9_IntShiftRight_49U_6U_32U_mbits_fixed_rshift_rg_a = { chn_trt_in_rsci_d_mxwt[440:392], 63'b000000000000000000000000000000000000000000000000000000000000000 };
endmodule
