module \$paramod\SDP_Y_CORE_mgc_in_wire_v1\rscid=7\width=10 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:376" *)
  output [9:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:377" *)
  input [9:0] z;
  assign d = z;
endmodule
