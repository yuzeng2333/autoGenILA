module SDP_Y_CORE_leading_sign_49_0(mantissa, rtn);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:244" *)
  wire _000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:258" *)
  wire _001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:258" *)
  wire _002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:271" *)
  wire _003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:277" *)
  wire _004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *)
  wire _005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *)
  wire _006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:280" *)
  wire _007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *)
  wire _008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *)
  wire _009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *)
  wire _010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *)
  wire _011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:283" *)
  wire _012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:286" *)
  wire _013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *)
  wire _014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *)
  wire _015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:288" *)
  wire _016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:289" *)
  wire _017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:290" *)
  wire _018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *)
  wire _019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *)
  wire _020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *)
  wire _021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *)
  wire _022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:293" *)
  wire _023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *)
  wire _024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *)
  wire _025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *)
  wire _026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:295" *)
  wire _027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *)
  wire _033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *)
  wire _040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *)
  wire _041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *)
  wire _042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *)
  wire _043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:307" *)
  wire _050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:307" *)
  wire _051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:236" *)
  wire _052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:243" *)
  wire _053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:249" *)
  wire _054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:257" *)
  wire _055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:263" *)
  wire _056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:270" *)
  wire _057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:232" *)
  wire _058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:233" *)
  wire _059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:234" *)
  wire _060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:238" *)
  wire _061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:239" *)
  wire _062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:240" *)
  wire _063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:245" *)
  wire _064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:246" *)
  wire _065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:247" *)
  wire _066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:251" *)
  wire _067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:252" *)
  wire _068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:253" *)
  wire _069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:259" *)
  wire _070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:260" *)
  wire _071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:261" *)
  wire _072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:265" *)
  wire _073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:266" *)
  wire _074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:267" *)
  wire _075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *)
  wire _076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *)
  wire _080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *)
  wire _084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *)
  wire _085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *)
  wire _086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *)
  wire _087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:275" *)
  wire _088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:277" *)
  wire _089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *)
  wire _090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *)
  wire _091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *)
  wire _092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:280" *)
  wire _093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *)
  wire _094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *)
  wire _095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *)
  wire _096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *)
  wire _097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *)
  wire _098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:283" *)
  wire _099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *)
  wire _100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *)
  wire _101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:290" *)
  wire _102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *)
  wire _103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *)
  wire _104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *)
  wire _105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *)
  wire _106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *)
  wire _107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *)
  wire _108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:295" *)
  wire _109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *)
  wire _110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *)
  wire _111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *)
  wire _120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *)
  wire _121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *)
  wire _131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *)
  wire _132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *)
  wire _133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *)
  wire _134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *)
  wire _135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *)
  wire _136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *)
  wire _137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *)
  wire _138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:275" *)
  wire _145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:277" *)
  wire _146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:280" *)
  wire _147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *)
  wire _148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *)
  wire _149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:283" *)
  wire _150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:285" *)
  wire _151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *)
  wire _152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:289" *)
  wire _153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:290" *)
  wire _154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:292" *)
  wire _155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *)
  wire _156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:295" *)
  wire _157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *)
  wire _158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *)
  wire _160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *)
  wire _161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *)
  wire _162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *)
  wire _164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *)
  wire _165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *)
  wire _166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *)
  wire _167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *)
  wire _168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *)
  wire _169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *)
  wire _170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:230" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:227" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:226" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:228" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:229" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:211" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:199" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:212" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:200" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:213" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:201" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:203" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:191" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:204" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:192" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:205" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:193" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:206" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:194" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:207" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:195" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:202" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:190" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:208" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:196" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:209" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:197" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:210" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:198" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:218" *)
  wire c_h_1_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:219" *)
  wire c_h_1_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:220" *)
  wire c_h_1_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:221" *)
  wire c_h_1_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:214" *)
  wire c_h_1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:222" *)
  wire c_h_1_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:223" *)
  wire c_h_1_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:224" *)
  wire c_h_1_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:225" *)
  wire c_h_1_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:215" *)
  wire c_h_1_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:216" *)
  wire c_h_1_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:217" *)
  wire c_h_1_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:187" *)
  input [48:0] mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:188" *)
  output [5:0] rtn;
  assign c_h_1_2 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:235" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3 = _052_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:237" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:241" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:242" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _053_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:244" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:244" *) c_h_1_5;
  assign c_h_1_9 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:248" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3 = _054_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:250" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  assign c_h_1_12 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:254" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:255" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:256" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign _001_ = _055_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:258" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  assign _002_ = _001_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:258" *) c_h_1_12;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5 = _002_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:258" *) c_h_1_13;
  assign c_h_1_17 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:262" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3 = _056_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:264" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  assign c_h_1_20 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:268" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:269" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign _003_ = _057_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:271" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4 = _003_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:271" *) c_h_1_20;
  assign c_h_1_22 = c_h_1_21 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:272" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_23 = c_h_1_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:273" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl = c_h_1_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:275" *) _145_;
  assign _004_ = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:277" *) _146_;
  assign _005_ = c_h_1_21 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *) _090_;
  assign _006_ = _091_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl = _004_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *) _092_;
  assign _007_ = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:280" *) _147_;
  assign _008_ = c_h_1_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *) _148_;
  assign _009_ = _095_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *) c_h_1_14;
  assign _010_ = _007_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *) _096_;
  assign _011_ = c_h_1_17 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *) _149_;
  assign _012_ = _150_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:283" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl = _010_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:283" *) _099_;
  assign _013_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:286" *) _151_;
  assign _014_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *) _152_;
  assign _015_ = _100_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *) c_h_1_6;
  assign _016_ = _013_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:288" *) _101_;
  assign _017_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:289" *) _153_;
  assign _018_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:290" *) _154_;
  assign _019_ = _102_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *) c_h_1_13;
  assign _020_ = _017_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *) _103_;
  assign _021_ = _104_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *) c_h_1_14;
  assign _022_ = _016_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *) _105_;
  assign _023_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:293" *) _155_;
  assign _024_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *) _156_;
  assign _025_ = _106_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *) c_h_1_21;
  assign _026_ = _023_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *) _107_;
  assign _027_ = _157_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:295" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl = _022_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:295" *) _109_;
  assign _028_ = _159_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) c_h_1_2;
  assign _029_ = _111_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) _113_;
  assign _030_ = _161_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) c_h_1_5;
  assign _031_ = _115_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) _117_;
  assign _032_ = _118_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) c_h_1_6;
  assign _033_ = _029_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *) _119_;
  assign _034_ = _163_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) c_h_1_9;
  assign _035_ = _121_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) _123_;
  assign _036_ = _165_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) c_h_1_12;
  assign _037_ = _125_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _127_;
  assign _038_ = _128_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) c_h_1_13;
  assign _039_ = _035_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _129_;
  assign _040_ = _130_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *) c_h_1_14;
  assign _041_ = _033_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *) _131_;
  assign _042_ = _167_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *) c_h_1_17;
  assign _043_ = _133_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *) _135_;
  assign _044_ = _169_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) c_h_1_20;
  assign _045_ = _137_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _139_;
  assign _046_ = _140_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) c_h_1_21;
  assign _047_ = _043_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _141_;
  assign _048_ = _170_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) c_h_1_23;
  assign _049_ = _041_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _143_;
  assign _050_ = _144_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:307" *) c_h_1_22;
  assign _051_ = _050_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:307" *) c_h_1_23;
  assign _052_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:236" *) mantissa[42:41];
  assign _053_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:243" *) mantissa[34:33];
  assign _054_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:249" *) mantissa[26:25];
  assign _055_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:257" *) mantissa[18:17];
  assign _056_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:263" *) mantissa[10:9];
  assign _057_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:270" *) mantissa[2:1];
  assign _058_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:232" *) mantissa[46:45];
  assign _059_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:233" *) mantissa[48:47];
  assign _060_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:234" *) mantissa[44:43];
  assign _061_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:238" *) mantissa[38:37];
  assign _062_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:239" *) mantissa[40:39];
  assign _063_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:240" *) mantissa[36:35];
  assign _064_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:245" *) mantissa[30:29];
  assign _065_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:246" *) mantissa[32:31];
  assign _066_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:247" *) mantissa[28:27];
  assign _067_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:251" *) mantissa[22:21];
  assign _068_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:252" *) mantissa[24:23];
  assign _069_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:253" *) mantissa[20:19];
  assign _070_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:259" *) mantissa[14:13];
  assign _071_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:260" *) mantissa[16:15];
  assign _072_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:261" *) mantissa[12:11];
  assign _073_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:265" *) mantissa[6:5];
  assign _074_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:266" *) mantissa[8:7];
  assign _075_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:267" *) mantissa[4:3];
  assign _076_ = mantissa[47:46] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *) 1'b1;
  assign _077_ = mantissa[43:42] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) 1'b1;
  assign _078_ = mantissa[39:38] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) 1'b1;
  assign _079_ = mantissa[35:34] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) 1'b1;
  assign _080_ = mantissa[31:30] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *) 1'b1;
  assign _081_ = mantissa[27:26] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) 1'b1;
  assign _082_ = mantissa[23:22] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) 1'b1;
  assign _083_ = mantissa[19:18] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) 1'b1;
  assign _084_ = mantissa[15:14] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *) 1'b1;
  assign _085_ = mantissa[11:10] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *) 1'b1;
  assign _086_ = mantissa[7:6] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *) 1'b1;
  assign _087_ = mantissa[3:2] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *) 1'b1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:232" *) _058_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:233" *) _059_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:234" *) _060_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:238" *) _061_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:239" *) _062_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:240" *) _063_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:245" *) _064_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:246" *) _065_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:247" *) _066_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:251" *) _067_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:252" *) _068_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:253" *) _069_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:259" *) _070_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:260" *) _071_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:261" *) _072_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:265" *) _073_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:266" *) _074_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:267" *) _075_;
  assign _088_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:275" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign _089_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:277" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign _090_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign _091_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *) _005_;
  assign _092_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:278" *) _006_;
  assign _093_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:280" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign _094_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign _095_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *) _008_;
  assign _096_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *) _009_;
  assign _097_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign _098_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *) _011_;
  assign _099_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:283" *) _012_;
  assign _100_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *) _014_;
  assign _101_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *) _015_;
  assign _102_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:290" *) _018_;
  assign _103_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *) _019_;
  assign _104_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *) _020_;
  assign _105_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:291" *) _021_;
  assign _106_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *) _024_;
  assign _107_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *) _025_;
  assign _108_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *) _026_;
  assign _109_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:295" *) _027_;
  assign _110_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *) _076_;
  assign _111_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *) _158_;
  assign _112_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) _077_;
  assign _113_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) _028_;
  assign _114_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) _078_;
  assign _115_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) _160_;
  assign _116_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) _079_;
  assign _117_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) _030_;
  assign _118_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) _031_;
  assign _119_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) _032_;
  assign _120_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *) _080_;
  assign _121_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *) _162_;
  assign _122_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) _081_;
  assign _123_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) _034_;
  assign _124_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) _082_;
  assign _125_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) _164_;
  assign _126_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _083_;
  assign _127_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _036_;
  assign _128_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _037_;
  assign _129_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _038_;
  assign _130_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _039_;
  assign _131_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *) _040_;
  assign _132_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *) _084_;
  assign _133_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *) _166_;
  assign _134_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *) _085_;
  assign _135_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *) _042_;
  assign _136_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *) _086_;
  assign _137_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *) _168_;
  assign _138_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *) _087_;
  assign _139_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _044_;
  assign _140_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _045_;
  assign _141_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _046_;
  assign _142_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _047_;
  assign _143_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) _048_;
  assign _144_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) mantissa[0];
  assign _145_ = c_h_1_22 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:275" *) _088_;
  assign _146_ = c_h_1_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:277" *) _089_;
  assign _147_ = c_h_1_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:280" *) _093_;
  assign _148_ = c_h_1_12 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:281" *) _094_;
  assign _149_ = c_h_1_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:282" *) _097_;
  assign _150_ = _098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:283" *) c_h_1_22;
  assign _151_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:285" *) _058_;
  assign _152_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:287" *) _061_;
  assign _153_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:289" *) _064_;
  assign _154_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:290" *) _067_;
  assign _155_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:292" *) _070_;
  assign _156_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:294" *) _073_;
  assign _157_ = _108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:295" *) c_h_1_22;
  assign _158_ = mantissa[48] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:297" *) _110_;
  assign _159_ = mantissa[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) _112_;
  assign _160_ = mantissa[40] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:298" *) _114_;
  assign _161_ = mantissa[36] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:299" *) _116_;
  assign _162_ = mantissa[32] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:300" *) _120_;
  assign _163_ = mantissa[28] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) _122_;
  assign _164_ = mantissa[24] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:301" *) _124_;
  assign _165_ = mantissa[20] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:302" *) _126_;
  assign _166_ = mantissa[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:303" *) _132_;
  assign _167_ = mantissa[12] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:304" *) _134_;
  assign _168_ = mantissa[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *) _136_;
  assign _169_ = mantissa[4] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:305" *) _138_;
  assign _170_ = _142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:306" *) c_h_1_22;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl = _049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:307" *) _051_;
  assign rtn = { c_h_1_23, IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl, IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl };
endmodule
