module bar__DOT__i1(
__START__,
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
in,
rcon,
out_1,
out_2,
__COUNTER_start__n0
);
input            __START__;
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg    [127:0] in;
output reg      [7:0] rcon;
output reg    [127:0] out_1;
output reg    [127:0] out_2;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire            __START__;
wire    [127:0] bv_128_0_n1;
wire      [7:0] bv_8_0_n583;
wire      [7:0] bv_8_100_n417;
wire      [7:0] bv_8_101_n261;
wire      [7:0] bv_8_102_n176;
wire      [7:0] bv_8_103_n525;
wire      [7:0] bv_8_104_n39;
wire      [7:0] bv_8_105_n113;
wire      [7:0] bv_8_106_n516;
wire      [7:0] bv_8_107_n513;
wire      [7:0] bv_8_108_n272;
wire      [7:0] bv_8_109_n289;
wire      [7:0] bv_8_10_n343;
wire      [7:0] bv_8_110_n504;
wire      [7:0] bv_8_111_n501;
wire      [7:0] bv_8_112_n188;
wire      [7:0] bv_8_113_n495;
wire      [7:0] bv_8_114_n491;
wire      [7:0] bv_8_115_n408;
wire      [7:0] bv_8_116_n211;
wire      [7:0] bv_8_117_n484;
wire      [7:0] bv_8_118_n480;
wire      [7:0] bv_8_119_n477;
wire      [7:0] bv_8_11_n359;
wire      [7:0] bv_8_120_n243;
wire      [7:0] bv_8_121_n302;
wire      [7:0] bv_8_122_n257;
wire      [7:0] bv_8_123_n467;
wire      [7:0] bv_8_124_n463;
wire      [7:0] bv_8_125_n460;
wire      [7:0] bv_8_126_n423;
wire      [7:0] bv_8_127_n455;
wire      [7:0] bv_8_128_n452;
wire      [7:0] bv_8_129_n401;
wire      [7:0] bv_8_12_n450;
wire      [7:0] bv_8_130_n445;
wire      [7:0] bv_8_131_n442;
wire      [7:0] bv_8_132_n438;
wire      [7:0] bv_8_133_n435;
wire      [7:0] bv_8_134_n142;
wire      [7:0] bv_8_135_n91;
wire      [7:0] bv_8_136_n381;
wire      [7:0] bv_8_137_n59;
wire      [7:0] bv_8_138_n192;
wire      [7:0] bv_8_139_n195;
wire      [7:0] bv_8_13_n55;
wire      [7:0] bv_8_140_n67;
wire      [7:0] bv_8_141_n285;
wire      [7:0] bv_8_142_n105;
wire      [7:0] bv_8_143_n406;
wire      [7:0] bv_8_144_n385;
wire      [7:0] bv_8_145_n312;
wire      [7:0] bv_8_146_n396;
wire      [7:0] bv_8_147_n393;
wire      [7:0] bv_8_148_n102;
wire      [7:0] bv_8_149_n308;
wire      [7:0] bv_8_14_n161;
wire      [7:0] bv_8_150_n383;
wire      [7:0] bv_8_151_n379;
wire      [7:0] bv_8_152_n121;
wire      [7:0] bv_8_153_n31;
wire      [7:0] bv_8_154_n371;
wire      [7:0] bv_8_155_n98;
wire      [7:0] bv_8_156_n365;
wire      [7:0] bv_8_157_n361;
wire      [7:0] bv_8_158_n130;
wire      [7:0] bv_8_159_n355;
wire      [7:0] bv_8_15_n23;
wire      [7:0] bv_8_160_n352;
wire      [7:0] bv_8_161_n63;
wire      [7:0] bv_8_162_n345;
wire      [7:0] bv_8_163_n341;
wire      [7:0] bv_8_164_n337;
wire      [7:0] bv_8_165_n333;
wire      [7:0] bv_8_166_n228;
wire      [7:0] bv_8_167_n326;
wire      [7:0] bv_8_168_n323;
wire      [7:0] bv_8_169_n276;
wire      [7:0] bv_8_16_n465;
wire      [7:0] bv_8_170_n318;
wire      [7:0] bv_8_171_n314;
wire      [7:0] bv_8_172_n310;
wire      [7:0] bv_8_173_n306;
wire      [7:0] bv_8_174_n254;
wire      [7:0] bv_8_175_n300;
wire      [7:0] bv_8_176_n19;
wire      [7:0] bv_8_177_n295;
wire      [7:0] bv_8_178_n291;
wire      [7:0] bv_8_179_n287;
wire      [7:0] bv_8_17_n117;
wire      [7:0] bv_8_180_n224;
wire      [7:0] bv_8_181_n180;
wire      [7:0] bv_8_182_n278;
wire      [7:0] bv_8_183_n274;
wire      [7:0] bv_8_184_n270;
wire      [7:0] bv_8_185_n146;
wire      [7:0] bv_8_186_n247;
wire      [7:0] bv_8_187_n11;
wire      [7:0] bv_8_188_n259;
wire      [7:0] bv_8_189_n199;
wire      [7:0] bv_8_18_n644;
wire      [7:0] bv_8_190_n252;
wire      [7:0] bv_8_191_n51;
wire      [7:0] bv_8_192_n245;
wire      [7:0] bv_8_193_n138;
wire      [7:0] bv_8_194_n238;
wire      [7:0] bv_8_195_n234;
wire      [7:0] bv_8_196_n230;
wire      [7:0] bv_8_197_n226;
wire      [7:0] bv_8_198_n221;
wire      [7:0] bv_8_199_n219;
wire      [7:0] bv_8_19_n447;
wire      [7:0] bv_8_1_n753;
wire      [7:0] bv_8_200_n216;
wire      [7:0] bv_8_201_n213;
wire      [7:0] bv_8_202_n209;
wire      [7:0] bv_8_203_n205;
wire      [7:0] bv_8_204_n201;
wire      [7:0] bv_8_205_n197;
wire      [7:0] bv_8_206_n83;
wire      [7:0] bv_8_207_n190;
wire      [7:0] bv_8_208_n186;
wire      [7:0] bv_8_209_n182;
wire      [7:0] bv_8_20_n369;
wire      [7:0] bv_8_210_n178;
wire      [7:0] bv_8_211_n174;
wire      [7:0] bv_8_212_n170;
wire      [7:0] bv_8_213_n166;
wire      [7:0] bv_8_214_n163;
wire      [7:0] bv_8_215_n159;
wire      [7:0] bv_8_216_n155;
wire      [7:0] bv_8_217_n109;
wire      [7:0] bv_8_218_n148;
wire      [7:0] bv_8_219_n144;
wire      [7:0] bv_8_21_n674;
wire      [7:0] bv_8_220_n140;
wire      [7:0] bv_8_221_n136;
wire      [7:0] bv_8_222_n132;
wire      [7:0] bv_8_223_n71;
wire      [7:0] bv_8_224_n126;
wire      [7:0] bv_8_225_n123;
wire      [7:0] bv_8_226_n119;
wire      [7:0] bv_8_227_n115;
wire      [7:0] bv_8_228_n111;
wire      [7:0] bv_8_229_n107;
wire      [7:0] bv_8_22_n7;
wire      [7:0] bv_8_230_n47;
wire      [7:0] bv_8_231_n100;
wire      [7:0] bv_8_232_n96;
wire      [7:0] bv_8_233_n87;
wire      [7:0] bv_8_234_n89;
wire      [7:0] bv_8_235_n85;
wire      [7:0] bv_8_236_n81;
wire      [7:0] bv_8_237_n77;
wire      [7:0] bv_8_238_n73;
wire      [7:0] bv_8_239_n69;
wire      [7:0] bv_8_23_n430;
wire      [7:0] bv_8_240_n65;
wire      [7:0] bv_8_241_n61;
wire      [7:0] bv_8_242_n57;
wire      [7:0] bv_8_243_n53;
wire      [7:0] bv_8_244_n49;
wire      [7:0] bv_8_245_n45;
wire      [7:0] bv_8_246_n41;
wire      [7:0] bv_8_247_n37;
wire      [7:0] bv_8_248_n33;
wire      [7:0] bv_8_249_n29;
wire      [7:0] bv_8_24_n659;
wire      [7:0] bv_8_250_n25;
wire      [7:0] bv_8_251_n21;
wire      [7:0] bv_8_252_n17;
wire      [7:0] bv_8_253_n13;
wire      [7:0] bv_8_254_n9;
wire      [7:0] bv_8_255_n5;
wire      [7:0] bv_8_25_n411;
wire      [7:0] bv_8_26_n619;
wire      [7:0] bv_8_27_n616;
wire      [7:0] bv_8_28_n232;
wire      [7:0] bv_8_29_n134;
wire      [7:0] bv_8_2_n518;
wire      [7:0] bv_8_30_n94;
wire      [7:0] bv_8_31_n207;
wire      [7:0] bv_8_32_n576;
wire      [7:0] bv_8_33_n469;
wire      [7:0] bv_8_34_n391;
wire      [7:0] bv_8_35_n664;
wire      [7:0] bv_8_36_n331;
wire      [7:0] bv_8_37_n240;
wire      [7:0] bv_8_38_n693;
wire      [7:0] bv_8_39_n635;
wire      [7:0] bv_8_3_n168;
wire      [7:0] bv_8_40_n75;
wire      [7:0] bv_8_41_n597;
wire      [7:0] bv_8_42_n388;
wire      [7:0] bv_8_43_n682;
wire      [7:0] bv_8_44_n622;
wire      [7:0] bv_8_45_n27;
wire      [7:0] bv_8_46_n236;
wire      [7:0] bv_8_47_n592;
wire      [7:0] bv_8_48_n669;
wire      [7:0] bv_8_49_n666;
wire      [7:0] bv_8_4_n671;
wire      [7:0] bv_8_50_n350;
wire      [7:0] bv_8_51_n529;
wire      [7:0] bv_8_52_n657;
wire      [7:0] bv_8_53_n153;
wire      [7:0] bv_8_54_n651;
wire      [7:0] bv_8_55_n293;
wire      [7:0] bv_8_56_n482;
wire      [7:0] bv_8_57_n559;
wire      [7:0] bv_8_58_n347;
wire      [7:0] bv_8_59_n604;
wire      [7:0] bv_8_5_n653;
wire      [7:0] bv_8_60_n508;
wire      [7:0] bv_8_61_n420;
wire      [7:0] bv_8_62_n184;
wire      [7:0] bv_8_63_n629;
wire      [7:0] bv_8_64_n493;
wire      [7:0] bv_8_65_n35;
wire      [7:0] bv_8_66_n43;
wire      [7:0] bv_8_67_n535;
wire      [7:0] bv_8_68_n433;
wire      [7:0] bv_8_69_n523;
wire      [7:0] bv_8_6_n335;
wire      [7:0] bv_8_70_n377;
wire      [7:0] bv_8_71_n608;
wire      [7:0] bv_8_72_n172;
wire      [7:0] bv_8_73_n339;
wire      [7:0] bv_8_74_n555;
wire      [7:0] bv_8_75_n203;
wire      [7:0] bv_8_76_n552;
wire      [7:0] bv_8_77_n532;
wire      [7:0] bv_8_78_n280;
wire      [7:0] bv_8_79_n398;
wire      [7:0] bv_8_7_n647;
wire      [7:0] bv_8_80_n511;
wire      [7:0] bv_8_81_n499;
wire      [7:0] bv_8_82_n581;
wire      [7:0] bv_8_83_n578;
wire      [7:0] bv_8_84_n15;
wire      [7:0] bv_8_85_n79;
wire      [7:0] bv_8_86_n268;
wire      [7:0] bv_8_87_n150;
wire      [7:0] bv_8_88_n549;
wire      [7:0] bv_8_89_n564;
wire      [7:0] bv_8_8_n250;
wire      [7:0] bv_8_90_n561;
wire      [7:0] bv_8_91_n557;
wire      [7:0] bv_8_92_n328;
wire      [7:0] bv_8_93_n414;
wire      [7:0] bv_8_94_n363;
wire      [7:0] bv_8_95_n440;
wire      [7:0] bv_8_96_n404;
wire      [7:0] bv_8_97_n157;
wire      [7:0] bv_8_98_n316;
wire      [7:0] bv_8_99_n537;
wire      [7:0] bv_8_9_n627;
wire            clk;
(* keep *) wire    [127:0] in_randinit;
wire            n10;
wire      [7:0] n1000;
wire      [7:0] n1001;
wire      [7:0] n1002;
wire      [7:0] n1003;
wire      [7:0] n1004;
wire      [7:0] n1005;
wire      [7:0] n1006;
wire      [7:0] n1007;
wire      [7:0] n1008;
wire      [7:0] n1009;
wire            n101;
wire      [7:0] n1010;
wire      [7:0] n1011;
wire      [7:0] n1012;
wire      [7:0] n1013;
wire      [7:0] n1014;
wire      [7:0] n1015;
wire      [7:0] n1016;
wire      [7:0] n1017;
wire      [7:0] n1018;
wire      [7:0] n1019;
wire      [7:0] n1020;
wire      [7:0] n1021;
wire      [7:0] n1022;
wire      [7:0] n1023;
wire      [7:0] n1024;
wire      [7:0] n1025;
wire      [7:0] n1026;
wire      [7:0] n1027;
wire      [7:0] n1028;
wire      [7:0] n1029;
wire      [7:0] n103;
wire      [7:0] n1030;
wire            n1031;
wire      [7:0] n1032;
wire            n1033;
wire      [7:0] n1034;
wire            n1035;
wire      [7:0] n1036;
wire            n1037;
wire      [7:0] n1038;
wire            n1039;
wire            n104;
wire      [7:0] n1040;
wire            n1041;
wire      [7:0] n1042;
wire            n1043;
wire      [7:0] n1044;
wire            n1045;
wire      [7:0] n1046;
wire            n1047;
wire      [7:0] n1048;
wire            n1049;
wire      [7:0] n1050;
wire            n1051;
wire      [7:0] n1052;
wire            n1053;
wire      [7:0] n1054;
wire            n1055;
wire      [7:0] n1056;
wire            n1057;
wire      [7:0] n1058;
wire            n1059;
wire      [7:0] n106;
wire      [7:0] n1060;
wire            n1061;
wire      [7:0] n1062;
wire            n1063;
wire      [7:0] n1064;
wire            n1065;
wire      [7:0] n1066;
wire            n1067;
wire      [7:0] n1068;
wire            n1069;
wire      [7:0] n1070;
wire            n1071;
wire      [7:0] n1072;
wire            n1073;
wire      [7:0] n1074;
wire            n1075;
wire      [7:0] n1076;
wire            n1077;
wire      [7:0] n1078;
wire            n1079;
wire            n108;
wire      [7:0] n1080;
wire            n1081;
wire      [7:0] n1082;
wire            n1083;
wire      [7:0] n1084;
wire            n1085;
wire      [7:0] n1086;
wire            n1087;
wire      [7:0] n1088;
wire            n1089;
wire      [7:0] n1090;
wire            n1091;
wire      [7:0] n1092;
wire            n1093;
wire      [7:0] n1094;
wire            n1095;
wire      [7:0] n1096;
wire            n1097;
wire      [7:0] n1098;
wire            n1099;
wire      [7:0] n110;
wire      [7:0] n1100;
wire            n1101;
wire      [7:0] n1102;
wire            n1103;
wire      [7:0] n1104;
wire            n1105;
wire      [7:0] n1106;
wire            n1107;
wire      [7:0] n1108;
wire            n1109;
wire      [7:0] n1110;
wire            n1111;
wire      [7:0] n1112;
wire            n1113;
wire      [7:0] n1114;
wire            n1115;
wire      [7:0] n1116;
wire            n1117;
wire      [7:0] n1118;
wire            n1119;
wire            n112;
wire      [7:0] n1120;
wire            n1121;
wire      [7:0] n1122;
wire            n1123;
wire      [7:0] n1124;
wire            n1125;
wire      [7:0] n1126;
wire            n1127;
wire      [7:0] n1128;
wire            n1129;
wire      [7:0] n1130;
wire            n1131;
wire      [7:0] n1132;
wire            n1133;
wire      [7:0] n1134;
wire            n1135;
wire      [7:0] n1136;
wire            n1137;
wire      [7:0] n1138;
wire            n1139;
wire      [7:0] n114;
wire      [7:0] n1140;
wire            n1141;
wire      [7:0] n1142;
wire            n1143;
wire      [7:0] n1144;
wire            n1145;
wire      [7:0] n1146;
wire            n1147;
wire      [7:0] n1148;
wire            n1149;
wire      [7:0] n1150;
wire            n1151;
wire      [7:0] n1152;
wire            n1153;
wire      [7:0] n1154;
wire            n1155;
wire      [7:0] n1156;
wire            n1157;
wire      [7:0] n1158;
wire            n1159;
wire            n116;
wire      [7:0] n1160;
wire            n1161;
wire      [7:0] n1162;
wire            n1163;
wire      [7:0] n1164;
wire            n1165;
wire      [7:0] n1166;
wire            n1167;
wire      [7:0] n1168;
wire            n1169;
wire      [7:0] n1170;
wire            n1171;
wire      [7:0] n1172;
wire            n1173;
wire      [7:0] n1174;
wire            n1175;
wire      [7:0] n1176;
wire            n1177;
wire      [7:0] n1178;
wire            n1179;
wire      [7:0] n118;
wire      [7:0] n1180;
wire            n1181;
wire      [7:0] n1182;
wire            n1183;
wire      [7:0] n1184;
wire            n1185;
wire      [7:0] n1186;
wire            n1187;
wire      [7:0] n1188;
wire            n1189;
wire      [7:0] n1190;
wire            n1191;
wire      [7:0] n1192;
wire            n1193;
wire      [7:0] n1194;
wire            n1195;
wire      [7:0] n1196;
wire            n1197;
wire      [7:0] n1198;
wire            n1199;
wire      [7:0] n12;
wire            n120;
wire      [7:0] n1200;
wire            n1201;
wire      [7:0] n1202;
wire            n1203;
wire      [7:0] n1204;
wire            n1205;
wire      [7:0] n1206;
wire            n1207;
wire      [7:0] n1208;
wire            n1209;
wire      [7:0] n1210;
wire            n1211;
wire      [7:0] n1212;
wire            n1213;
wire      [7:0] n1214;
wire            n1215;
wire      [7:0] n1216;
wire            n1217;
wire      [7:0] n1218;
wire            n1219;
wire      [7:0] n122;
wire      [7:0] n1220;
wire            n1221;
wire      [7:0] n1222;
wire            n1223;
wire      [7:0] n1224;
wire            n1225;
wire      [7:0] n1226;
wire            n1227;
wire      [7:0] n1228;
wire            n1229;
wire      [7:0] n1230;
wire            n1231;
wire      [7:0] n1232;
wire            n1233;
wire      [7:0] n1234;
wire            n1235;
wire      [7:0] n1236;
wire            n1237;
wire      [7:0] n1238;
wire            n1239;
wire            n124;
wire      [7:0] n1240;
wire            n1241;
wire      [7:0] n1242;
wire            n1243;
wire      [7:0] n1244;
wire            n1245;
wire      [7:0] n1246;
wire            n1247;
wire      [7:0] n1248;
wire            n1249;
wire      [7:0] n125;
wire      [7:0] n1250;
wire            n1251;
wire      [7:0] n1252;
wire            n1253;
wire      [7:0] n1254;
wire            n1255;
wire      [7:0] n1256;
wire            n1257;
wire      [7:0] n1258;
wire            n1259;
wire      [7:0] n1260;
wire            n1261;
wire      [7:0] n1262;
wire            n1263;
wire      [7:0] n1264;
wire            n1265;
wire      [7:0] n1266;
wire            n1267;
wire      [7:0] n1268;
wire            n1269;
wire            n127;
wire      [7:0] n1270;
wire            n1271;
wire      [7:0] n1272;
wire            n1273;
wire      [7:0] n1274;
wire            n1275;
wire      [7:0] n1276;
wire            n1277;
wire      [7:0] n1278;
wire            n1279;
wire      [7:0] n128;
wire      [7:0] n1280;
wire            n1281;
wire      [7:0] n1282;
wire            n1283;
wire      [7:0] n1284;
wire            n1285;
wire      [7:0] n1286;
wire            n1287;
wire      [7:0] n1288;
wire            n1289;
wire            n129;
wire      [7:0] n1290;
wire            n1291;
wire      [7:0] n1292;
wire            n1293;
wire      [7:0] n1294;
wire            n1295;
wire      [7:0] n1296;
wire            n1297;
wire      [7:0] n1298;
wire            n1299;
wire      [7:0] n1300;
wire            n1301;
wire      [7:0] n1302;
wire            n1303;
wire      [7:0] n1304;
wire            n1305;
wire      [7:0] n1306;
wire            n1307;
wire      [7:0] n1308;
wire            n1309;
wire      [7:0] n131;
wire      [7:0] n1310;
wire            n1311;
wire      [7:0] n1312;
wire            n1313;
wire      [7:0] n1314;
wire            n1315;
wire      [7:0] n1316;
wire            n1317;
wire      [7:0] n1318;
wire            n1319;
wire      [7:0] n1320;
wire            n1321;
wire      [7:0] n1322;
wire            n1323;
wire      [7:0] n1324;
wire            n1325;
wire      [7:0] n1326;
wire            n1327;
wire      [7:0] n1328;
wire            n1329;
wire            n133;
wire      [7:0] n1330;
wire            n1331;
wire      [7:0] n1332;
wire            n1333;
wire      [7:0] n1334;
wire            n1335;
wire      [7:0] n1336;
wire            n1337;
wire      [7:0] n1338;
wire            n1339;
wire      [7:0] n1340;
wire            n1341;
wire      [7:0] n1342;
wire            n1343;
wire      [7:0] n1344;
wire            n1345;
wire      [7:0] n1346;
wire            n1347;
wire      [7:0] n1348;
wire            n1349;
wire      [7:0] n135;
wire      [7:0] n1350;
wire            n1351;
wire      [7:0] n1352;
wire            n1353;
wire      [7:0] n1354;
wire            n1355;
wire      [7:0] n1356;
wire            n1357;
wire      [7:0] n1358;
wire            n1359;
wire      [7:0] n1360;
wire            n1361;
wire      [7:0] n1362;
wire            n1363;
wire      [7:0] n1364;
wire            n1365;
wire      [7:0] n1366;
wire            n1367;
wire      [7:0] n1368;
wire            n1369;
wire            n137;
wire      [7:0] n1370;
wire            n1371;
wire      [7:0] n1372;
wire            n1373;
wire      [7:0] n1374;
wire            n1375;
wire      [7:0] n1376;
wire            n1377;
wire      [7:0] n1378;
wire            n1379;
wire      [7:0] n1380;
wire            n1381;
wire      [7:0] n1382;
wire            n1383;
wire      [7:0] n1384;
wire            n1385;
wire      [7:0] n1386;
wire            n1387;
wire      [7:0] n1388;
wire            n1389;
wire      [7:0] n139;
wire      [7:0] n1390;
wire            n1391;
wire      [7:0] n1392;
wire            n1393;
wire      [7:0] n1394;
wire            n1395;
wire      [7:0] n1396;
wire            n1397;
wire      [7:0] n1398;
wire            n1399;
wire            n14;
wire      [7:0] n1400;
wire            n1401;
wire      [7:0] n1402;
wire            n1403;
wire      [7:0] n1404;
wire            n1405;
wire      [7:0] n1406;
wire            n1407;
wire      [7:0] n1408;
wire            n1409;
wire            n141;
wire      [7:0] n1410;
wire            n1411;
wire      [7:0] n1412;
wire            n1413;
wire      [7:0] n1414;
wire            n1415;
wire      [7:0] n1416;
wire            n1417;
wire      [7:0] n1418;
wire            n1419;
wire      [7:0] n1420;
wire            n1421;
wire      [7:0] n1422;
wire            n1423;
wire      [7:0] n1424;
wire            n1425;
wire      [7:0] n1426;
wire            n1427;
wire      [7:0] n1428;
wire            n1429;
wire      [7:0] n143;
wire      [7:0] n1430;
wire            n1431;
wire      [7:0] n1432;
wire            n1433;
wire      [7:0] n1434;
wire            n1435;
wire      [7:0] n1436;
wire            n1437;
wire      [7:0] n1438;
wire            n1439;
wire      [7:0] n1440;
wire            n1441;
wire      [7:0] n1442;
wire            n1443;
wire      [7:0] n1444;
wire            n1445;
wire      [7:0] n1446;
wire            n1447;
wire      [7:0] n1448;
wire            n1449;
wire            n145;
wire      [7:0] n1450;
wire            n1451;
wire      [7:0] n1452;
wire            n1453;
wire      [7:0] n1454;
wire            n1455;
wire      [7:0] n1456;
wire            n1457;
wire      [7:0] n1458;
wire            n1459;
wire      [7:0] n1460;
wire            n1461;
wire      [7:0] n1462;
wire            n1463;
wire      [7:0] n1464;
wire            n1465;
wire      [7:0] n1466;
wire            n1467;
wire      [7:0] n1468;
wire            n1469;
wire      [7:0] n147;
wire      [7:0] n1470;
wire            n1471;
wire      [7:0] n1472;
wire            n1473;
wire      [7:0] n1474;
wire            n1475;
wire      [7:0] n1476;
wire            n1477;
wire      [7:0] n1478;
wire            n1479;
wire      [7:0] n1480;
wire            n1481;
wire      [7:0] n1482;
wire            n1483;
wire      [7:0] n1484;
wire            n1485;
wire      [7:0] n1486;
wire            n1487;
wire      [7:0] n1488;
wire            n1489;
wire            n149;
wire      [7:0] n1490;
wire            n1491;
wire      [7:0] n1492;
wire            n1493;
wire      [7:0] n1494;
wire            n1495;
wire      [7:0] n1496;
wire            n1497;
wire      [7:0] n1498;
wire            n1499;
wire      [7:0] n1500;
wire            n1501;
wire      [7:0] n1502;
wire            n1503;
wire      [7:0] n1504;
wire            n1505;
wire      [7:0] n1506;
wire            n1507;
wire      [7:0] n1508;
wire            n1509;
wire      [7:0] n151;
wire      [7:0] n1510;
wire            n1511;
wire      [7:0] n1512;
wire            n1513;
wire      [7:0] n1514;
wire            n1515;
wire      [7:0] n1516;
wire            n1517;
wire      [7:0] n1518;
wire            n1519;
wire            n152;
wire      [7:0] n1520;
wire            n1521;
wire      [7:0] n1522;
wire            n1523;
wire      [7:0] n1524;
wire            n1525;
wire      [7:0] n1526;
wire            n1527;
wire      [7:0] n1528;
wire            n1529;
wire      [7:0] n1530;
wire            n1531;
wire      [7:0] n1532;
wire            n1533;
wire      [7:0] n1534;
wire            n1535;
wire      [7:0] n1536;
wire            n1537;
wire      [7:0] n1538;
wire            n1539;
wire      [7:0] n154;
wire      [7:0] n1540;
wire            n1541;
wire      [7:0] n1542;
wire      [7:0] n1543;
wire      [7:0] n1544;
wire      [7:0] n1545;
wire      [7:0] n1546;
wire      [7:0] n1547;
wire      [7:0] n1548;
wire      [7:0] n1549;
wire      [7:0] n1550;
wire      [7:0] n1551;
wire      [7:0] n1552;
wire      [7:0] n1553;
wire      [7:0] n1554;
wire      [7:0] n1555;
wire      [7:0] n1556;
wire      [7:0] n1557;
wire      [7:0] n1558;
wire      [7:0] n1559;
wire            n156;
wire      [7:0] n1560;
wire      [7:0] n1561;
wire      [7:0] n1562;
wire      [7:0] n1563;
wire      [7:0] n1564;
wire      [7:0] n1565;
wire      [7:0] n1566;
wire      [7:0] n1567;
wire      [7:0] n1568;
wire      [7:0] n1569;
wire      [7:0] n1570;
wire      [7:0] n1571;
wire      [7:0] n1572;
wire      [7:0] n1573;
wire      [7:0] n1574;
wire      [7:0] n1575;
wire      [7:0] n1576;
wire      [7:0] n1577;
wire      [7:0] n1578;
wire      [7:0] n1579;
wire      [7:0] n158;
wire      [7:0] n1580;
wire      [7:0] n1581;
wire      [7:0] n1582;
wire      [7:0] n1583;
wire      [7:0] n1584;
wire      [7:0] n1585;
wire      [7:0] n1586;
wire      [7:0] n1587;
wire      [7:0] n1588;
wire      [7:0] n1589;
wire      [7:0] n1590;
wire      [7:0] n1591;
wire      [7:0] n1592;
wire      [7:0] n1593;
wire      [7:0] n1594;
wire      [7:0] n1595;
wire      [7:0] n1596;
wire      [7:0] n1597;
wire      [7:0] n1598;
wire      [7:0] n1599;
wire      [7:0] n16;
wire            n160;
wire      [7:0] n1600;
wire      [7:0] n1601;
wire      [7:0] n1602;
wire      [7:0] n1603;
wire      [7:0] n1604;
wire      [7:0] n1605;
wire      [7:0] n1606;
wire      [7:0] n1607;
wire      [7:0] n1608;
wire      [7:0] n1609;
wire      [7:0] n1610;
wire      [7:0] n1611;
wire      [7:0] n1612;
wire      [7:0] n1613;
wire      [7:0] n1614;
wire      [7:0] n1615;
wire      [7:0] n1616;
wire      [7:0] n1617;
wire      [7:0] n1618;
wire      [7:0] n1619;
wire      [7:0] n162;
wire      [7:0] n1620;
wire      [7:0] n1621;
wire      [7:0] n1622;
wire      [7:0] n1623;
wire      [7:0] n1624;
wire      [7:0] n1625;
wire      [7:0] n1626;
wire      [7:0] n1627;
wire      [7:0] n1628;
wire      [7:0] n1629;
wire      [7:0] n1630;
wire      [7:0] n1631;
wire      [7:0] n1632;
wire      [7:0] n1633;
wire      [7:0] n1634;
wire      [7:0] n1635;
wire      [7:0] n1636;
wire      [7:0] n1637;
wire      [7:0] n1638;
wire      [7:0] n1639;
wire            n164;
wire      [7:0] n1640;
wire      [7:0] n1641;
wire      [7:0] n1642;
wire      [7:0] n1643;
wire      [7:0] n1644;
wire      [7:0] n1645;
wire      [7:0] n1646;
wire      [7:0] n1647;
wire      [7:0] n1648;
wire      [7:0] n1649;
wire      [7:0] n165;
wire      [7:0] n1650;
wire      [7:0] n1651;
wire      [7:0] n1652;
wire      [7:0] n1653;
wire      [7:0] n1654;
wire      [7:0] n1655;
wire      [7:0] n1656;
wire      [7:0] n1657;
wire      [7:0] n1658;
wire      [7:0] n1659;
wire      [7:0] n1660;
wire      [7:0] n1661;
wire      [7:0] n1662;
wire      [7:0] n1663;
wire      [7:0] n1664;
wire      [7:0] n1665;
wire      [7:0] n1666;
wire      [7:0] n1667;
wire      [7:0] n1668;
wire      [7:0] n1669;
wire            n167;
wire      [7:0] n1670;
wire      [7:0] n1671;
wire      [7:0] n1672;
wire      [7:0] n1673;
wire      [7:0] n1674;
wire      [7:0] n1675;
wire      [7:0] n1676;
wire      [7:0] n1677;
wire      [7:0] n1678;
wire      [7:0] n1679;
wire      [7:0] n1680;
wire      [7:0] n1681;
wire      [7:0] n1682;
wire      [7:0] n1683;
wire      [7:0] n1684;
wire      [7:0] n1685;
wire      [7:0] n1686;
wire      [7:0] n1687;
wire      [7:0] n1688;
wire      [7:0] n1689;
wire      [7:0] n169;
wire      [7:0] n1690;
wire      [7:0] n1691;
wire      [7:0] n1692;
wire      [7:0] n1693;
wire      [7:0] n1694;
wire      [7:0] n1695;
wire      [7:0] n1696;
wire      [7:0] n1697;
wire      [7:0] n1698;
wire      [7:0] n1699;
wire      [7:0] n1700;
wire      [7:0] n1701;
wire      [7:0] n1702;
wire      [7:0] n1703;
wire      [7:0] n1704;
wire      [7:0] n1705;
wire      [7:0] n1706;
wire      [7:0] n1707;
wire      [7:0] n1708;
wire      [7:0] n1709;
wire            n171;
wire      [7:0] n1710;
wire      [7:0] n1711;
wire      [7:0] n1712;
wire      [7:0] n1713;
wire      [7:0] n1714;
wire      [7:0] n1715;
wire      [7:0] n1716;
wire      [7:0] n1717;
wire      [7:0] n1718;
wire      [7:0] n1719;
wire      [7:0] n1720;
wire      [7:0] n1721;
wire      [7:0] n1722;
wire      [7:0] n1723;
wire      [7:0] n1724;
wire      [7:0] n1725;
wire      [7:0] n1726;
wire      [7:0] n1727;
wire      [7:0] n1728;
wire      [7:0] n1729;
wire      [7:0] n173;
wire      [7:0] n1730;
wire      [7:0] n1731;
wire      [7:0] n1732;
wire      [7:0] n1733;
wire      [7:0] n1734;
wire      [7:0] n1735;
wire      [7:0] n1736;
wire      [7:0] n1737;
wire      [7:0] n1738;
wire      [7:0] n1739;
wire      [7:0] n1740;
wire      [7:0] n1741;
wire      [7:0] n1742;
wire      [7:0] n1743;
wire      [7:0] n1744;
wire      [7:0] n1745;
wire      [7:0] n1746;
wire      [7:0] n1747;
wire      [7:0] n1748;
wire      [7:0] n1749;
wire            n175;
wire      [7:0] n1750;
wire      [7:0] n1751;
wire      [7:0] n1752;
wire      [7:0] n1753;
wire      [7:0] n1754;
wire      [7:0] n1755;
wire      [7:0] n1756;
wire      [7:0] n1757;
wire      [7:0] n1758;
wire      [7:0] n1759;
wire      [7:0] n1760;
wire      [7:0] n1761;
wire      [7:0] n1762;
wire      [7:0] n1763;
wire      [7:0] n1764;
wire      [7:0] n1765;
wire      [7:0] n1766;
wire      [7:0] n1767;
wire      [7:0] n1768;
wire      [7:0] n1769;
wire      [7:0] n177;
wire      [7:0] n1770;
wire      [7:0] n1771;
wire      [7:0] n1772;
wire      [7:0] n1773;
wire      [7:0] n1774;
wire      [7:0] n1775;
wire      [7:0] n1776;
wire      [7:0] n1777;
wire      [7:0] n1778;
wire      [7:0] n1779;
wire      [7:0] n1780;
wire      [7:0] n1781;
wire      [7:0] n1782;
wire      [7:0] n1783;
wire      [7:0] n1784;
wire      [7:0] n1785;
wire      [7:0] n1786;
wire      [7:0] n1787;
wire      [7:0] n1788;
wire      [7:0] n1789;
wire            n179;
wire      [7:0] n1790;
wire      [7:0] n1791;
wire      [7:0] n1792;
wire      [7:0] n1793;
wire      [7:0] n1794;
wire      [7:0] n1795;
wire      [7:0] n1796;
wire      [7:0] n1797;
wire      [7:0] n1798;
wire     [15:0] n1799;
wire            n18;
wire      [7:0] n1800;
wire      [7:0] n1801;
wire            n1802;
wire      [7:0] n1803;
wire            n1804;
wire      [7:0] n1805;
wire            n1806;
wire      [7:0] n1807;
wire            n1808;
wire      [7:0] n1809;
wire      [7:0] n181;
wire            n1810;
wire      [7:0] n1811;
wire            n1812;
wire      [7:0] n1813;
wire            n1814;
wire      [7:0] n1815;
wire            n1816;
wire      [7:0] n1817;
wire            n1818;
wire      [7:0] n1819;
wire            n1820;
wire      [7:0] n1821;
wire            n1822;
wire      [7:0] n1823;
wire            n1824;
wire      [7:0] n1825;
wire            n1826;
wire      [7:0] n1827;
wire            n1828;
wire      [7:0] n1829;
wire            n183;
wire            n1830;
wire      [7:0] n1831;
wire            n1832;
wire      [7:0] n1833;
wire            n1834;
wire      [7:0] n1835;
wire            n1836;
wire      [7:0] n1837;
wire            n1838;
wire      [7:0] n1839;
wire            n1840;
wire      [7:0] n1841;
wire            n1842;
wire      [7:0] n1843;
wire            n1844;
wire      [7:0] n1845;
wire            n1846;
wire      [7:0] n1847;
wire            n1848;
wire      [7:0] n1849;
wire      [7:0] n185;
wire            n1850;
wire      [7:0] n1851;
wire            n1852;
wire      [7:0] n1853;
wire            n1854;
wire      [7:0] n1855;
wire            n1856;
wire      [7:0] n1857;
wire            n1858;
wire      [7:0] n1859;
wire            n1860;
wire      [7:0] n1861;
wire            n1862;
wire      [7:0] n1863;
wire            n1864;
wire      [7:0] n1865;
wire            n1866;
wire      [7:0] n1867;
wire            n1868;
wire      [7:0] n1869;
wire            n187;
wire            n1870;
wire      [7:0] n1871;
wire            n1872;
wire      [7:0] n1873;
wire            n1874;
wire      [7:0] n1875;
wire            n1876;
wire      [7:0] n1877;
wire            n1878;
wire      [7:0] n1879;
wire            n1880;
wire      [7:0] n1881;
wire            n1882;
wire      [7:0] n1883;
wire            n1884;
wire      [7:0] n1885;
wire            n1886;
wire      [7:0] n1887;
wire            n1888;
wire      [7:0] n1889;
wire      [7:0] n189;
wire            n1890;
wire      [7:0] n1891;
wire            n1892;
wire      [7:0] n1893;
wire            n1894;
wire      [7:0] n1895;
wire            n1896;
wire      [7:0] n1897;
wire            n1898;
wire      [7:0] n1899;
wire            n1900;
wire      [7:0] n1901;
wire            n1902;
wire      [7:0] n1903;
wire            n1904;
wire      [7:0] n1905;
wire            n1906;
wire      [7:0] n1907;
wire            n1908;
wire      [7:0] n1909;
wire            n191;
wire            n1910;
wire      [7:0] n1911;
wire            n1912;
wire      [7:0] n1913;
wire            n1914;
wire      [7:0] n1915;
wire            n1916;
wire      [7:0] n1917;
wire            n1918;
wire      [7:0] n1919;
wire            n1920;
wire      [7:0] n1921;
wire            n1922;
wire      [7:0] n1923;
wire            n1924;
wire      [7:0] n1925;
wire            n1926;
wire      [7:0] n1927;
wire            n1928;
wire      [7:0] n1929;
wire      [7:0] n193;
wire            n1930;
wire      [7:0] n1931;
wire            n1932;
wire      [7:0] n1933;
wire            n1934;
wire      [7:0] n1935;
wire            n1936;
wire      [7:0] n1937;
wire            n1938;
wire      [7:0] n1939;
wire            n194;
wire            n1940;
wire      [7:0] n1941;
wire            n1942;
wire      [7:0] n1943;
wire            n1944;
wire      [7:0] n1945;
wire            n1946;
wire      [7:0] n1947;
wire            n1948;
wire      [7:0] n1949;
wire            n1950;
wire      [7:0] n1951;
wire            n1952;
wire      [7:0] n1953;
wire            n1954;
wire      [7:0] n1955;
wire            n1956;
wire      [7:0] n1957;
wire            n1958;
wire      [7:0] n1959;
wire      [7:0] n196;
wire            n1960;
wire      [7:0] n1961;
wire            n1962;
wire      [7:0] n1963;
wire            n1964;
wire      [7:0] n1965;
wire            n1966;
wire      [7:0] n1967;
wire            n1968;
wire      [7:0] n1969;
wire            n1970;
wire      [7:0] n1971;
wire            n1972;
wire      [7:0] n1973;
wire            n1974;
wire      [7:0] n1975;
wire            n1976;
wire      [7:0] n1977;
wire            n1978;
wire      [7:0] n1979;
wire            n198;
wire            n1980;
wire      [7:0] n1981;
wire            n1982;
wire      [7:0] n1983;
wire            n1984;
wire      [7:0] n1985;
wire            n1986;
wire      [7:0] n1987;
wire            n1988;
wire      [7:0] n1989;
wire            n1990;
wire      [7:0] n1991;
wire            n1992;
wire      [7:0] n1993;
wire            n1994;
wire      [7:0] n1995;
wire            n1996;
wire      [7:0] n1997;
wire            n1998;
wire      [7:0] n1999;
wire      [7:0] n2;
wire      [7:0] n20;
wire      [7:0] n200;
wire            n2000;
wire      [7:0] n2001;
wire            n2002;
wire      [7:0] n2003;
wire            n2004;
wire      [7:0] n2005;
wire            n2006;
wire      [7:0] n2007;
wire            n2008;
wire      [7:0] n2009;
wire            n2010;
wire      [7:0] n2011;
wire            n2012;
wire      [7:0] n2013;
wire            n2014;
wire      [7:0] n2015;
wire            n2016;
wire      [7:0] n2017;
wire            n2018;
wire      [7:0] n2019;
wire            n202;
wire            n2020;
wire      [7:0] n2021;
wire            n2022;
wire      [7:0] n2023;
wire            n2024;
wire      [7:0] n2025;
wire            n2026;
wire      [7:0] n2027;
wire            n2028;
wire      [7:0] n2029;
wire            n2030;
wire      [7:0] n2031;
wire            n2032;
wire      [7:0] n2033;
wire            n2034;
wire      [7:0] n2035;
wire            n2036;
wire      [7:0] n2037;
wire            n2038;
wire      [7:0] n2039;
wire      [7:0] n204;
wire            n2040;
wire      [7:0] n2041;
wire            n2042;
wire      [7:0] n2043;
wire            n2044;
wire      [7:0] n2045;
wire            n2046;
wire      [7:0] n2047;
wire            n2048;
wire      [7:0] n2049;
wire            n2050;
wire      [7:0] n2051;
wire            n2052;
wire      [7:0] n2053;
wire            n2054;
wire      [7:0] n2055;
wire            n2056;
wire      [7:0] n2057;
wire            n2058;
wire      [7:0] n2059;
wire            n206;
wire            n2060;
wire      [7:0] n2061;
wire            n2062;
wire      [7:0] n2063;
wire            n2064;
wire      [7:0] n2065;
wire            n2066;
wire      [7:0] n2067;
wire            n2068;
wire      [7:0] n2069;
wire            n2070;
wire      [7:0] n2071;
wire            n2072;
wire      [7:0] n2073;
wire            n2074;
wire      [7:0] n2075;
wire            n2076;
wire      [7:0] n2077;
wire            n2078;
wire      [7:0] n2079;
wire      [7:0] n208;
wire            n2080;
wire      [7:0] n2081;
wire            n2082;
wire      [7:0] n2083;
wire            n2084;
wire      [7:0] n2085;
wire            n2086;
wire      [7:0] n2087;
wire            n2088;
wire      [7:0] n2089;
wire            n2090;
wire      [7:0] n2091;
wire            n2092;
wire      [7:0] n2093;
wire            n2094;
wire      [7:0] n2095;
wire            n2096;
wire      [7:0] n2097;
wire            n2098;
wire      [7:0] n2099;
wire            n210;
wire            n2100;
wire      [7:0] n2101;
wire            n2102;
wire      [7:0] n2103;
wire            n2104;
wire      [7:0] n2105;
wire            n2106;
wire      [7:0] n2107;
wire            n2108;
wire      [7:0] n2109;
wire            n2110;
wire      [7:0] n2111;
wire            n2112;
wire      [7:0] n2113;
wire            n2114;
wire      [7:0] n2115;
wire            n2116;
wire      [7:0] n2117;
wire            n2118;
wire      [7:0] n2119;
wire      [7:0] n212;
wire            n2120;
wire      [7:0] n2121;
wire            n2122;
wire      [7:0] n2123;
wire            n2124;
wire      [7:0] n2125;
wire            n2126;
wire      [7:0] n2127;
wire            n2128;
wire      [7:0] n2129;
wire            n2130;
wire      [7:0] n2131;
wire            n2132;
wire      [7:0] n2133;
wire            n2134;
wire      [7:0] n2135;
wire            n2136;
wire      [7:0] n2137;
wire            n2138;
wire      [7:0] n2139;
wire            n214;
wire            n2140;
wire      [7:0] n2141;
wire            n2142;
wire      [7:0] n2143;
wire            n2144;
wire      [7:0] n2145;
wire            n2146;
wire      [7:0] n2147;
wire            n2148;
wire      [7:0] n2149;
wire      [7:0] n215;
wire            n2150;
wire      [7:0] n2151;
wire            n2152;
wire      [7:0] n2153;
wire            n2154;
wire      [7:0] n2155;
wire            n2156;
wire      [7:0] n2157;
wire            n2158;
wire      [7:0] n2159;
wire            n2160;
wire      [7:0] n2161;
wire            n2162;
wire      [7:0] n2163;
wire            n2164;
wire      [7:0] n2165;
wire            n2166;
wire      [7:0] n2167;
wire            n2168;
wire      [7:0] n2169;
wire            n217;
wire            n2170;
wire      [7:0] n2171;
wire            n2172;
wire      [7:0] n2173;
wire            n2174;
wire      [7:0] n2175;
wire            n2176;
wire      [7:0] n2177;
wire            n2178;
wire      [7:0] n2179;
wire      [7:0] n218;
wire            n2180;
wire      [7:0] n2181;
wire            n2182;
wire      [7:0] n2183;
wire            n2184;
wire      [7:0] n2185;
wire            n2186;
wire      [7:0] n2187;
wire            n2188;
wire      [7:0] n2189;
wire            n2190;
wire      [7:0] n2191;
wire            n2192;
wire      [7:0] n2193;
wire            n2194;
wire      [7:0] n2195;
wire            n2196;
wire      [7:0] n2197;
wire            n2198;
wire      [7:0] n2199;
wire            n22;
wire            n220;
wire            n2200;
wire      [7:0] n2201;
wire            n2202;
wire      [7:0] n2203;
wire            n2204;
wire      [7:0] n2205;
wire            n2206;
wire      [7:0] n2207;
wire            n2208;
wire      [7:0] n2209;
wire            n2210;
wire      [7:0] n2211;
wire            n2212;
wire      [7:0] n2213;
wire            n2214;
wire      [7:0] n2215;
wire            n2216;
wire      [7:0] n2217;
wire            n2218;
wire      [7:0] n2219;
wire      [7:0] n222;
wire            n2220;
wire      [7:0] n2221;
wire            n2222;
wire      [7:0] n2223;
wire            n2224;
wire      [7:0] n2225;
wire            n2226;
wire      [7:0] n2227;
wire            n2228;
wire      [7:0] n2229;
wire            n223;
wire            n2230;
wire      [7:0] n2231;
wire            n2232;
wire      [7:0] n2233;
wire            n2234;
wire      [7:0] n2235;
wire            n2236;
wire      [7:0] n2237;
wire            n2238;
wire      [7:0] n2239;
wire            n2240;
wire      [7:0] n2241;
wire            n2242;
wire      [7:0] n2243;
wire            n2244;
wire      [7:0] n2245;
wire            n2246;
wire      [7:0] n2247;
wire            n2248;
wire      [7:0] n2249;
wire      [7:0] n225;
wire            n2250;
wire      [7:0] n2251;
wire            n2252;
wire      [7:0] n2253;
wire            n2254;
wire      [7:0] n2255;
wire            n2256;
wire      [7:0] n2257;
wire            n2258;
wire      [7:0] n2259;
wire            n2260;
wire      [7:0] n2261;
wire            n2262;
wire      [7:0] n2263;
wire            n2264;
wire      [7:0] n2265;
wire            n2266;
wire      [7:0] n2267;
wire            n2268;
wire      [7:0] n2269;
wire            n227;
wire            n2270;
wire      [7:0] n2271;
wire            n2272;
wire      [7:0] n2273;
wire            n2274;
wire      [7:0] n2275;
wire            n2276;
wire      [7:0] n2277;
wire            n2278;
wire      [7:0] n2279;
wire            n2280;
wire      [7:0] n2281;
wire            n2282;
wire      [7:0] n2283;
wire            n2284;
wire      [7:0] n2285;
wire            n2286;
wire      [7:0] n2287;
wire            n2288;
wire      [7:0] n2289;
wire      [7:0] n229;
wire            n2290;
wire      [7:0] n2291;
wire            n2292;
wire      [7:0] n2293;
wire            n2294;
wire      [7:0] n2295;
wire            n2296;
wire      [7:0] n2297;
wire            n2298;
wire      [7:0] n2299;
wire            n2300;
wire      [7:0] n2301;
wire            n2302;
wire      [7:0] n2303;
wire            n2304;
wire      [7:0] n2305;
wire            n2306;
wire      [7:0] n2307;
wire            n2308;
wire      [7:0] n2309;
wire            n231;
wire            n2310;
wire      [7:0] n2311;
wire            n2312;
wire      [7:0] n2313;
wire      [7:0] n2314;
wire      [7:0] n2315;
wire      [7:0] n2316;
wire      [7:0] n2317;
wire      [7:0] n2318;
wire      [7:0] n2319;
wire      [7:0] n2320;
wire      [7:0] n2321;
wire      [7:0] n2322;
wire      [7:0] n2323;
wire      [7:0] n2324;
wire      [7:0] n2325;
wire      [7:0] n2326;
wire      [7:0] n2327;
wire      [7:0] n2328;
wire      [7:0] n2329;
wire      [7:0] n233;
wire      [7:0] n2330;
wire      [7:0] n2331;
wire      [7:0] n2332;
wire      [7:0] n2333;
wire      [7:0] n2334;
wire      [7:0] n2335;
wire      [7:0] n2336;
wire      [7:0] n2337;
wire      [7:0] n2338;
wire      [7:0] n2339;
wire      [7:0] n2340;
wire      [7:0] n2341;
wire      [7:0] n2342;
wire      [7:0] n2343;
wire      [7:0] n2344;
wire      [7:0] n2345;
wire      [7:0] n2346;
wire      [7:0] n2347;
wire      [7:0] n2348;
wire      [7:0] n2349;
wire            n235;
wire      [7:0] n2350;
wire      [7:0] n2351;
wire      [7:0] n2352;
wire      [7:0] n2353;
wire      [7:0] n2354;
wire      [7:0] n2355;
wire      [7:0] n2356;
wire      [7:0] n2357;
wire      [7:0] n2358;
wire      [7:0] n2359;
wire      [7:0] n2360;
wire      [7:0] n2361;
wire      [7:0] n2362;
wire      [7:0] n2363;
wire      [7:0] n2364;
wire      [7:0] n2365;
wire      [7:0] n2366;
wire      [7:0] n2367;
wire      [7:0] n2368;
wire      [7:0] n2369;
wire      [7:0] n237;
wire      [7:0] n2370;
wire      [7:0] n2371;
wire      [7:0] n2372;
wire      [7:0] n2373;
wire      [7:0] n2374;
wire      [7:0] n2375;
wire      [7:0] n2376;
wire      [7:0] n2377;
wire      [7:0] n2378;
wire      [7:0] n2379;
wire      [7:0] n2380;
wire      [7:0] n2381;
wire      [7:0] n2382;
wire      [7:0] n2383;
wire      [7:0] n2384;
wire      [7:0] n2385;
wire      [7:0] n2386;
wire      [7:0] n2387;
wire      [7:0] n2388;
wire      [7:0] n2389;
wire            n239;
wire      [7:0] n2390;
wire      [7:0] n2391;
wire      [7:0] n2392;
wire      [7:0] n2393;
wire      [7:0] n2394;
wire      [7:0] n2395;
wire      [7:0] n2396;
wire      [7:0] n2397;
wire      [7:0] n2398;
wire      [7:0] n2399;
wire      [7:0] n24;
wire      [7:0] n2400;
wire      [7:0] n2401;
wire      [7:0] n2402;
wire      [7:0] n2403;
wire      [7:0] n2404;
wire      [7:0] n2405;
wire      [7:0] n2406;
wire      [7:0] n2407;
wire      [7:0] n2408;
wire      [7:0] n2409;
wire      [7:0] n241;
wire      [7:0] n2410;
wire      [7:0] n2411;
wire      [7:0] n2412;
wire      [7:0] n2413;
wire      [7:0] n2414;
wire      [7:0] n2415;
wire      [7:0] n2416;
wire      [7:0] n2417;
wire      [7:0] n2418;
wire      [7:0] n2419;
wire            n242;
wire      [7:0] n2420;
wire      [7:0] n2421;
wire      [7:0] n2422;
wire      [7:0] n2423;
wire      [7:0] n2424;
wire      [7:0] n2425;
wire      [7:0] n2426;
wire      [7:0] n2427;
wire      [7:0] n2428;
wire      [7:0] n2429;
wire      [7:0] n2430;
wire      [7:0] n2431;
wire      [7:0] n2432;
wire      [7:0] n2433;
wire      [7:0] n2434;
wire      [7:0] n2435;
wire      [7:0] n2436;
wire      [7:0] n2437;
wire      [7:0] n2438;
wire      [7:0] n2439;
wire      [7:0] n244;
wire      [7:0] n2440;
wire      [7:0] n2441;
wire      [7:0] n2442;
wire      [7:0] n2443;
wire      [7:0] n2444;
wire      [7:0] n2445;
wire      [7:0] n2446;
wire      [7:0] n2447;
wire      [7:0] n2448;
wire      [7:0] n2449;
wire      [7:0] n2450;
wire      [7:0] n2451;
wire      [7:0] n2452;
wire      [7:0] n2453;
wire      [7:0] n2454;
wire      [7:0] n2455;
wire      [7:0] n2456;
wire      [7:0] n2457;
wire      [7:0] n2458;
wire      [7:0] n2459;
wire            n246;
wire      [7:0] n2460;
wire      [7:0] n2461;
wire      [7:0] n2462;
wire      [7:0] n2463;
wire      [7:0] n2464;
wire      [7:0] n2465;
wire      [7:0] n2466;
wire      [7:0] n2467;
wire      [7:0] n2468;
wire      [7:0] n2469;
wire      [7:0] n2470;
wire      [7:0] n2471;
wire      [7:0] n2472;
wire      [7:0] n2473;
wire      [7:0] n2474;
wire      [7:0] n2475;
wire      [7:0] n2476;
wire      [7:0] n2477;
wire      [7:0] n2478;
wire      [7:0] n2479;
wire      [7:0] n248;
wire      [7:0] n2480;
wire      [7:0] n2481;
wire      [7:0] n2482;
wire      [7:0] n2483;
wire      [7:0] n2484;
wire      [7:0] n2485;
wire      [7:0] n2486;
wire      [7:0] n2487;
wire      [7:0] n2488;
wire      [7:0] n2489;
wire            n249;
wire      [7:0] n2490;
wire      [7:0] n2491;
wire      [7:0] n2492;
wire      [7:0] n2493;
wire      [7:0] n2494;
wire      [7:0] n2495;
wire      [7:0] n2496;
wire      [7:0] n2497;
wire      [7:0] n2498;
wire      [7:0] n2499;
wire      [7:0] n2500;
wire      [7:0] n2501;
wire      [7:0] n2502;
wire      [7:0] n2503;
wire      [7:0] n2504;
wire      [7:0] n2505;
wire      [7:0] n2506;
wire      [7:0] n2507;
wire      [7:0] n2508;
wire      [7:0] n2509;
wire      [7:0] n251;
wire      [7:0] n2510;
wire      [7:0] n2511;
wire      [7:0] n2512;
wire      [7:0] n2513;
wire      [7:0] n2514;
wire      [7:0] n2515;
wire      [7:0] n2516;
wire      [7:0] n2517;
wire      [7:0] n2518;
wire      [7:0] n2519;
wire      [7:0] n2520;
wire      [7:0] n2521;
wire      [7:0] n2522;
wire      [7:0] n2523;
wire      [7:0] n2524;
wire      [7:0] n2525;
wire      [7:0] n2526;
wire      [7:0] n2527;
wire      [7:0] n2528;
wire      [7:0] n2529;
wire            n253;
wire      [7:0] n2530;
wire      [7:0] n2531;
wire      [7:0] n2532;
wire      [7:0] n2533;
wire      [7:0] n2534;
wire      [7:0] n2535;
wire      [7:0] n2536;
wire      [7:0] n2537;
wire      [7:0] n2538;
wire      [7:0] n2539;
wire      [7:0] n2540;
wire      [7:0] n2541;
wire      [7:0] n2542;
wire      [7:0] n2543;
wire      [7:0] n2544;
wire      [7:0] n2545;
wire      [7:0] n2546;
wire      [7:0] n2547;
wire      [7:0] n2548;
wire      [7:0] n2549;
wire      [7:0] n255;
wire      [7:0] n2550;
wire      [7:0] n2551;
wire      [7:0] n2552;
wire      [7:0] n2553;
wire      [7:0] n2554;
wire      [7:0] n2555;
wire      [7:0] n2556;
wire      [7:0] n2557;
wire      [7:0] n2558;
wire      [7:0] n2559;
wire            n256;
wire      [7:0] n2560;
wire      [7:0] n2561;
wire      [7:0] n2562;
wire      [7:0] n2563;
wire      [7:0] n2564;
wire      [7:0] n2565;
wire      [7:0] n2566;
wire      [7:0] n2567;
wire      [7:0] n2568;
wire      [7:0] n2569;
wire     [23:0] n2570;
wire      [7:0] n2571;
wire      [7:0] n2572;
wire            n2573;
wire      [7:0] n2574;
wire            n2575;
wire      [7:0] n2576;
wire            n2577;
wire      [7:0] n2578;
wire            n2579;
wire      [7:0] n258;
wire      [7:0] n2580;
wire            n2581;
wire      [7:0] n2582;
wire            n2583;
wire      [7:0] n2584;
wire            n2585;
wire      [7:0] n2586;
wire            n2587;
wire      [7:0] n2588;
wire            n2589;
wire      [7:0] n2590;
wire            n2591;
wire      [7:0] n2592;
wire            n2593;
wire      [7:0] n2594;
wire            n2595;
wire      [7:0] n2596;
wire            n2597;
wire      [7:0] n2598;
wire            n2599;
wire            n26;
wire            n260;
wire      [7:0] n2600;
wire            n2601;
wire      [7:0] n2602;
wire            n2603;
wire      [7:0] n2604;
wire            n2605;
wire      [7:0] n2606;
wire            n2607;
wire      [7:0] n2608;
wire            n2609;
wire      [7:0] n2610;
wire            n2611;
wire      [7:0] n2612;
wire            n2613;
wire      [7:0] n2614;
wire            n2615;
wire      [7:0] n2616;
wire            n2617;
wire      [7:0] n2618;
wire            n2619;
wire      [7:0] n262;
wire      [7:0] n2620;
wire            n2621;
wire      [7:0] n2622;
wire            n2623;
wire      [7:0] n2624;
wire            n2625;
wire      [7:0] n2626;
wire            n2627;
wire      [7:0] n2628;
wire            n2629;
wire            n263;
wire      [7:0] n2630;
wire            n2631;
wire      [7:0] n2632;
wire            n2633;
wire      [7:0] n2634;
wire            n2635;
wire      [7:0] n2636;
wire            n2637;
wire      [7:0] n2638;
wire            n2639;
wire      [7:0] n264;
wire      [7:0] n2640;
wire            n2641;
wire      [7:0] n2642;
wire            n2643;
wire      [7:0] n2644;
wire            n2645;
wire      [7:0] n2646;
wire            n2647;
wire      [7:0] n2648;
wire            n2649;
wire            n265;
wire      [7:0] n2650;
wire            n2651;
wire      [7:0] n2652;
wire            n2653;
wire      [7:0] n2654;
wire            n2655;
wire      [7:0] n2656;
wire            n2657;
wire      [7:0] n2658;
wire            n2659;
wire      [7:0] n266;
wire      [7:0] n2660;
wire            n2661;
wire      [7:0] n2662;
wire            n2663;
wire      [7:0] n2664;
wire            n2665;
wire      [7:0] n2666;
wire            n2667;
wire      [7:0] n2668;
wire            n2669;
wire            n267;
wire      [7:0] n2670;
wire            n2671;
wire      [7:0] n2672;
wire            n2673;
wire      [7:0] n2674;
wire            n2675;
wire      [7:0] n2676;
wire            n2677;
wire      [7:0] n2678;
wire            n2679;
wire      [7:0] n2680;
wire            n2681;
wire      [7:0] n2682;
wire            n2683;
wire      [7:0] n2684;
wire            n2685;
wire      [7:0] n2686;
wire            n2687;
wire      [7:0] n2688;
wire            n2689;
wire      [7:0] n269;
wire      [7:0] n2690;
wire            n2691;
wire      [7:0] n2692;
wire            n2693;
wire      [7:0] n2694;
wire            n2695;
wire      [7:0] n2696;
wire            n2697;
wire      [7:0] n2698;
wire            n2699;
wire      [7:0] n2700;
wire            n2701;
wire      [7:0] n2702;
wire            n2703;
wire      [7:0] n2704;
wire            n2705;
wire      [7:0] n2706;
wire            n2707;
wire      [7:0] n2708;
wire            n2709;
wire            n271;
wire      [7:0] n2710;
wire            n2711;
wire      [7:0] n2712;
wire            n2713;
wire      [7:0] n2714;
wire            n2715;
wire      [7:0] n2716;
wire            n2717;
wire      [7:0] n2718;
wire            n2719;
wire      [7:0] n2720;
wire            n2721;
wire      [7:0] n2722;
wire            n2723;
wire      [7:0] n2724;
wire            n2725;
wire      [7:0] n2726;
wire            n2727;
wire      [7:0] n2728;
wire            n2729;
wire      [7:0] n273;
wire      [7:0] n2730;
wire            n2731;
wire      [7:0] n2732;
wire            n2733;
wire      [7:0] n2734;
wire            n2735;
wire      [7:0] n2736;
wire            n2737;
wire      [7:0] n2738;
wire            n2739;
wire      [7:0] n2740;
wire            n2741;
wire      [7:0] n2742;
wire            n2743;
wire      [7:0] n2744;
wire            n2745;
wire      [7:0] n2746;
wire            n2747;
wire      [7:0] n2748;
wire            n2749;
wire            n275;
wire      [7:0] n2750;
wire            n2751;
wire      [7:0] n2752;
wire            n2753;
wire      [7:0] n2754;
wire            n2755;
wire      [7:0] n2756;
wire            n2757;
wire      [7:0] n2758;
wire            n2759;
wire      [7:0] n2760;
wire            n2761;
wire      [7:0] n2762;
wire            n2763;
wire      [7:0] n2764;
wire            n2765;
wire      [7:0] n2766;
wire            n2767;
wire      [7:0] n2768;
wire            n2769;
wire      [7:0] n277;
wire      [7:0] n2770;
wire            n2771;
wire      [7:0] n2772;
wire            n2773;
wire      [7:0] n2774;
wire            n2775;
wire      [7:0] n2776;
wire            n2777;
wire      [7:0] n2778;
wire            n2779;
wire      [7:0] n2780;
wire            n2781;
wire      [7:0] n2782;
wire            n2783;
wire      [7:0] n2784;
wire            n2785;
wire      [7:0] n2786;
wire            n2787;
wire      [7:0] n2788;
wire            n2789;
wire            n279;
wire      [7:0] n2790;
wire            n2791;
wire      [7:0] n2792;
wire            n2793;
wire      [7:0] n2794;
wire            n2795;
wire      [7:0] n2796;
wire            n2797;
wire      [7:0] n2798;
wire            n2799;
wire      [7:0] n28;
wire      [7:0] n2800;
wire            n2801;
wire      [7:0] n2802;
wire            n2803;
wire      [7:0] n2804;
wire            n2805;
wire      [7:0] n2806;
wire            n2807;
wire      [7:0] n2808;
wire            n2809;
wire      [7:0] n281;
wire      [7:0] n2810;
wire            n2811;
wire      [7:0] n2812;
wire            n2813;
wire      [7:0] n2814;
wire            n2815;
wire      [7:0] n2816;
wire            n2817;
wire      [7:0] n2818;
wire            n2819;
wire            n282;
wire      [7:0] n2820;
wire            n2821;
wire      [7:0] n2822;
wire            n2823;
wire      [7:0] n2824;
wire            n2825;
wire      [7:0] n2826;
wire            n2827;
wire      [7:0] n2828;
wire            n2829;
wire      [7:0] n283;
wire      [7:0] n2830;
wire            n2831;
wire      [7:0] n2832;
wire            n2833;
wire      [7:0] n2834;
wire            n2835;
wire      [7:0] n2836;
wire            n2837;
wire      [7:0] n2838;
wire            n2839;
wire            n284;
wire      [7:0] n2840;
wire            n2841;
wire      [7:0] n2842;
wire            n2843;
wire      [7:0] n2844;
wire            n2845;
wire      [7:0] n2846;
wire            n2847;
wire      [7:0] n2848;
wire            n2849;
wire      [7:0] n2850;
wire            n2851;
wire      [7:0] n2852;
wire            n2853;
wire      [7:0] n2854;
wire            n2855;
wire      [7:0] n2856;
wire            n2857;
wire      [7:0] n2858;
wire            n2859;
wire      [7:0] n286;
wire      [7:0] n2860;
wire            n2861;
wire      [7:0] n2862;
wire            n2863;
wire      [7:0] n2864;
wire            n2865;
wire      [7:0] n2866;
wire            n2867;
wire      [7:0] n2868;
wire            n2869;
wire      [7:0] n2870;
wire            n2871;
wire      [7:0] n2872;
wire            n2873;
wire      [7:0] n2874;
wire            n2875;
wire      [7:0] n2876;
wire            n2877;
wire      [7:0] n2878;
wire            n2879;
wire            n288;
wire      [7:0] n2880;
wire            n2881;
wire      [7:0] n2882;
wire            n2883;
wire      [7:0] n2884;
wire            n2885;
wire      [7:0] n2886;
wire            n2887;
wire      [7:0] n2888;
wire            n2889;
wire      [7:0] n2890;
wire            n2891;
wire      [7:0] n2892;
wire            n2893;
wire      [7:0] n2894;
wire            n2895;
wire      [7:0] n2896;
wire            n2897;
wire      [7:0] n2898;
wire            n2899;
wire      [7:0] n290;
wire      [7:0] n2900;
wire            n2901;
wire      [7:0] n2902;
wire            n2903;
wire      [7:0] n2904;
wire            n2905;
wire      [7:0] n2906;
wire            n2907;
wire      [7:0] n2908;
wire            n2909;
wire      [7:0] n2910;
wire            n2911;
wire      [7:0] n2912;
wire            n2913;
wire      [7:0] n2914;
wire            n2915;
wire      [7:0] n2916;
wire            n2917;
wire      [7:0] n2918;
wire            n2919;
wire            n292;
wire      [7:0] n2920;
wire            n2921;
wire      [7:0] n2922;
wire            n2923;
wire      [7:0] n2924;
wire            n2925;
wire      [7:0] n2926;
wire            n2927;
wire      [7:0] n2928;
wire            n2929;
wire      [7:0] n2930;
wire            n2931;
wire      [7:0] n2932;
wire            n2933;
wire      [7:0] n2934;
wire            n2935;
wire      [7:0] n2936;
wire            n2937;
wire      [7:0] n2938;
wire            n2939;
wire      [7:0] n294;
wire      [7:0] n2940;
wire            n2941;
wire      [7:0] n2942;
wire            n2943;
wire      [7:0] n2944;
wire            n2945;
wire      [7:0] n2946;
wire            n2947;
wire      [7:0] n2948;
wire            n2949;
wire      [7:0] n2950;
wire            n2951;
wire      [7:0] n2952;
wire            n2953;
wire      [7:0] n2954;
wire            n2955;
wire      [7:0] n2956;
wire            n2957;
wire      [7:0] n2958;
wire            n2959;
wire            n296;
wire      [7:0] n2960;
wire            n2961;
wire      [7:0] n2962;
wire            n2963;
wire      [7:0] n2964;
wire            n2965;
wire      [7:0] n2966;
wire            n2967;
wire      [7:0] n2968;
wire            n2969;
wire      [7:0] n297;
wire      [7:0] n2970;
wire            n2971;
wire      [7:0] n2972;
wire            n2973;
wire      [7:0] n2974;
wire            n2975;
wire      [7:0] n2976;
wire            n2977;
wire      [7:0] n2978;
wire            n2979;
wire            n298;
wire      [7:0] n2980;
wire            n2981;
wire      [7:0] n2982;
wire            n2983;
wire      [7:0] n2984;
wire            n2985;
wire      [7:0] n2986;
wire            n2987;
wire      [7:0] n2988;
wire            n2989;
wire      [7:0] n299;
wire      [7:0] n2990;
wire            n2991;
wire      [7:0] n2992;
wire            n2993;
wire      [7:0] n2994;
wire            n2995;
wire      [7:0] n2996;
wire            n2997;
wire      [7:0] n2998;
wire            n2999;
wire      [7:0] n3;
wire            n30;
wire      [7:0] n3000;
wire            n3001;
wire      [7:0] n3002;
wire            n3003;
wire      [7:0] n3004;
wire            n3005;
wire      [7:0] n3006;
wire            n3007;
wire      [7:0] n3008;
wire            n3009;
wire            n301;
wire      [7:0] n3010;
wire            n3011;
wire      [7:0] n3012;
wire            n3013;
wire      [7:0] n3014;
wire            n3015;
wire      [7:0] n3016;
wire            n3017;
wire      [7:0] n3018;
wire            n3019;
wire      [7:0] n3020;
wire            n3021;
wire      [7:0] n3022;
wire            n3023;
wire      [7:0] n3024;
wire            n3025;
wire      [7:0] n3026;
wire            n3027;
wire      [7:0] n3028;
wire            n3029;
wire      [7:0] n303;
wire      [7:0] n3030;
wire            n3031;
wire      [7:0] n3032;
wire            n3033;
wire      [7:0] n3034;
wire            n3035;
wire      [7:0] n3036;
wire            n3037;
wire      [7:0] n3038;
wire            n3039;
wire            n304;
wire      [7:0] n3040;
wire            n3041;
wire      [7:0] n3042;
wire            n3043;
wire      [7:0] n3044;
wire            n3045;
wire      [7:0] n3046;
wire            n3047;
wire      [7:0] n3048;
wire            n3049;
wire      [7:0] n305;
wire      [7:0] n3050;
wire            n3051;
wire      [7:0] n3052;
wire            n3053;
wire      [7:0] n3054;
wire            n3055;
wire      [7:0] n3056;
wire            n3057;
wire      [7:0] n3058;
wire            n3059;
wire      [7:0] n3060;
wire            n3061;
wire      [7:0] n3062;
wire            n3063;
wire      [7:0] n3064;
wire            n3065;
wire      [7:0] n3066;
wire            n3067;
wire      [7:0] n3068;
wire            n3069;
wire            n307;
wire      [7:0] n3070;
wire            n3071;
wire      [7:0] n3072;
wire            n3073;
wire      [7:0] n3074;
wire            n3075;
wire      [7:0] n3076;
wire            n3077;
wire      [7:0] n3078;
wire            n3079;
wire      [7:0] n3080;
wire            n3081;
wire      [7:0] n3082;
wire            n3083;
wire      [7:0] n3084;
wire      [7:0] n3085;
wire      [7:0] n3086;
wire      [7:0] n3087;
wire      [7:0] n3088;
wire      [7:0] n3089;
wire      [7:0] n309;
wire      [7:0] n3090;
wire      [7:0] n3091;
wire      [7:0] n3092;
wire      [7:0] n3093;
wire      [7:0] n3094;
wire      [7:0] n3095;
wire      [7:0] n3096;
wire      [7:0] n3097;
wire      [7:0] n3098;
wire      [7:0] n3099;
wire      [7:0] n3100;
wire      [7:0] n3101;
wire      [7:0] n3102;
wire      [7:0] n3103;
wire      [7:0] n3104;
wire      [7:0] n3105;
wire      [7:0] n3106;
wire      [7:0] n3107;
wire      [7:0] n3108;
wire      [7:0] n3109;
wire            n311;
wire      [7:0] n3110;
wire      [7:0] n3111;
wire      [7:0] n3112;
wire      [7:0] n3113;
wire      [7:0] n3114;
wire      [7:0] n3115;
wire      [7:0] n3116;
wire      [7:0] n3117;
wire      [7:0] n3118;
wire      [7:0] n3119;
wire      [7:0] n3120;
wire      [7:0] n3121;
wire      [7:0] n3122;
wire      [7:0] n3123;
wire      [7:0] n3124;
wire      [7:0] n3125;
wire      [7:0] n3126;
wire      [7:0] n3127;
wire      [7:0] n3128;
wire      [7:0] n3129;
wire      [7:0] n313;
wire      [7:0] n3130;
wire      [7:0] n3131;
wire      [7:0] n3132;
wire      [7:0] n3133;
wire      [7:0] n3134;
wire      [7:0] n3135;
wire      [7:0] n3136;
wire      [7:0] n3137;
wire      [7:0] n3138;
wire      [7:0] n3139;
wire      [7:0] n3140;
wire      [7:0] n3141;
wire      [7:0] n3142;
wire      [7:0] n3143;
wire      [7:0] n3144;
wire      [7:0] n3145;
wire      [7:0] n3146;
wire      [7:0] n3147;
wire      [7:0] n3148;
wire      [7:0] n3149;
wire            n315;
wire      [7:0] n3150;
wire      [7:0] n3151;
wire      [7:0] n3152;
wire      [7:0] n3153;
wire      [7:0] n3154;
wire      [7:0] n3155;
wire      [7:0] n3156;
wire      [7:0] n3157;
wire      [7:0] n3158;
wire      [7:0] n3159;
wire      [7:0] n3160;
wire      [7:0] n3161;
wire      [7:0] n3162;
wire      [7:0] n3163;
wire      [7:0] n3164;
wire      [7:0] n3165;
wire      [7:0] n3166;
wire      [7:0] n3167;
wire      [7:0] n3168;
wire      [7:0] n3169;
wire      [7:0] n317;
wire      [7:0] n3170;
wire      [7:0] n3171;
wire      [7:0] n3172;
wire      [7:0] n3173;
wire      [7:0] n3174;
wire      [7:0] n3175;
wire      [7:0] n3176;
wire      [7:0] n3177;
wire      [7:0] n3178;
wire      [7:0] n3179;
wire      [7:0] n3180;
wire      [7:0] n3181;
wire      [7:0] n3182;
wire      [7:0] n3183;
wire      [7:0] n3184;
wire      [7:0] n3185;
wire      [7:0] n3186;
wire      [7:0] n3187;
wire      [7:0] n3188;
wire      [7:0] n3189;
wire            n319;
wire      [7:0] n3190;
wire      [7:0] n3191;
wire      [7:0] n3192;
wire      [7:0] n3193;
wire      [7:0] n3194;
wire      [7:0] n3195;
wire      [7:0] n3196;
wire      [7:0] n3197;
wire      [7:0] n3198;
wire      [7:0] n3199;
wire      [7:0] n32;
wire      [7:0] n320;
wire      [7:0] n3200;
wire      [7:0] n3201;
wire      [7:0] n3202;
wire      [7:0] n3203;
wire      [7:0] n3204;
wire      [7:0] n3205;
wire      [7:0] n3206;
wire      [7:0] n3207;
wire      [7:0] n3208;
wire      [7:0] n3209;
wire            n321;
wire      [7:0] n3210;
wire      [7:0] n3211;
wire      [7:0] n3212;
wire      [7:0] n3213;
wire      [7:0] n3214;
wire      [7:0] n3215;
wire      [7:0] n3216;
wire      [7:0] n3217;
wire      [7:0] n3218;
wire      [7:0] n3219;
wire      [7:0] n322;
wire      [7:0] n3220;
wire      [7:0] n3221;
wire      [7:0] n3222;
wire      [7:0] n3223;
wire      [7:0] n3224;
wire      [7:0] n3225;
wire      [7:0] n3226;
wire      [7:0] n3227;
wire      [7:0] n3228;
wire      [7:0] n3229;
wire      [7:0] n3230;
wire      [7:0] n3231;
wire      [7:0] n3232;
wire      [7:0] n3233;
wire      [7:0] n3234;
wire      [7:0] n3235;
wire      [7:0] n3236;
wire      [7:0] n3237;
wire      [7:0] n3238;
wire      [7:0] n3239;
wire            n324;
wire      [7:0] n3240;
wire      [7:0] n3241;
wire      [7:0] n3242;
wire      [7:0] n3243;
wire      [7:0] n3244;
wire      [7:0] n3245;
wire      [7:0] n3246;
wire      [7:0] n3247;
wire      [7:0] n3248;
wire      [7:0] n3249;
wire      [7:0] n325;
wire      [7:0] n3250;
wire      [7:0] n3251;
wire      [7:0] n3252;
wire      [7:0] n3253;
wire      [7:0] n3254;
wire      [7:0] n3255;
wire      [7:0] n3256;
wire      [7:0] n3257;
wire      [7:0] n3258;
wire      [7:0] n3259;
wire      [7:0] n3260;
wire      [7:0] n3261;
wire      [7:0] n3262;
wire      [7:0] n3263;
wire      [7:0] n3264;
wire      [7:0] n3265;
wire      [7:0] n3266;
wire      [7:0] n3267;
wire      [7:0] n3268;
wire      [7:0] n3269;
wire            n327;
wire      [7:0] n3270;
wire      [7:0] n3271;
wire      [7:0] n3272;
wire      [7:0] n3273;
wire      [7:0] n3274;
wire      [7:0] n3275;
wire      [7:0] n3276;
wire      [7:0] n3277;
wire      [7:0] n3278;
wire      [7:0] n3279;
wire      [7:0] n3280;
wire      [7:0] n3281;
wire      [7:0] n3282;
wire      [7:0] n3283;
wire      [7:0] n3284;
wire      [7:0] n3285;
wire      [7:0] n3286;
wire      [7:0] n3287;
wire      [7:0] n3288;
wire      [7:0] n3289;
wire      [7:0] n329;
wire      [7:0] n3290;
wire      [7:0] n3291;
wire      [7:0] n3292;
wire      [7:0] n3293;
wire      [7:0] n3294;
wire      [7:0] n3295;
wire      [7:0] n3296;
wire      [7:0] n3297;
wire      [7:0] n3298;
wire      [7:0] n3299;
wire            n330;
wire      [7:0] n3300;
wire      [7:0] n3301;
wire      [7:0] n3302;
wire      [7:0] n3303;
wire      [7:0] n3304;
wire      [7:0] n3305;
wire      [7:0] n3306;
wire      [7:0] n3307;
wire      [7:0] n3308;
wire      [7:0] n3309;
wire      [7:0] n3310;
wire      [7:0] n3311;
wire      [7:0] n3312;
wire      [7:0] n3313;
wire      [7:0] n3314;
wire      [7:0] n3315;
wire      [7:0] n3316;
wire      [7:0] n3317;
wire      [7:0] n3318;
wire      [7:0] n3319;
wire      [7:0] n332;
wire      [7:0] n3320;
wire      [7:0] n3321;
wire      [7:0] n3322;
wire      [7:0] n3323;
wire      [7:0] n3324;
wire      [7:0] n3325;
wire      [7:0] n3326;
wire      [7:0] n3327;
wire      [7:0] n3328;
wire      [7:0] n3329;
wire      [7:0] n3330;
wire      [7:0] n3331;
wire      [7:0] n3332;
wire      [7:0] n3333;
wire      [7:0] n3334;
wire      [7:0] n3335;
wire      [7:0] n3336;
wire      [7:0] n3337;
wire      [7:0] n3338;
wire      [7:0] n3339;
wire            n334;
wire      [7:0] n3340;
wire     [31:0] n3341;
wire      [7:0] n3342;
wire      [7:0] n3343;
wire      [7:0] n3344;
wire      [7:0] n3345;
wire      [7:0] n3346;
wire     [39:0] n3347;
wire      [7:0] n3348;
wire      [7:0] n3349;
wire      [7:0] n3350;
wire      [7:0] n3351;
wire     [47:0] n3352;
wire      [7:0] n3353;
wire      [7:0] n3354;
wire      [7:0] n3355;
wire      [7:0] n3356;
wire     [55:0] n3357;
wire      [7:0] n3358;
wire      [7:0] n3359;
wire      [7:0] n336;
wire      [7:0] n3360;
wire      [7:0] n3361;
wire     [63:0] n3362;
wire      [7:0] n3363;
wire      [7:0] n3364;
wire      [7:0] n3365;
wire      [7:0] n3366;
wire      [7:0] n3367;
wire      [7:0] n3368;
wire      [7:0] n3369;
wire     [71:0] n3370;
wire      [7:0] n3371;
wire      [7:0] n3372;
wire      [7:0] n3373;
wire      [7:0] n3374;
wire      [7:0] n3375;
wire      [7:0] n3376;
wire     [79:0] n3377;
wire      [7:0] n3378;
wire      [7:0] n3379;
wire            n338;
wire      [7:0] n3380;
wire      [7:0] n3381;
wire      [7:0] n3382;
wire      [7:0] n3383;
wire     [87:0] n3384;
wire      [7:0] n3385;
wire      [7:0] n3386;
wire      [7:0] n3387;
wire      [7:0] n3388;
wire      [7:0] n3389;
wire      [7:0] n3390;
wire     [95:0] n3391;
wire      [7:0] n3392;
wire      [7:0] n3393;
wire      [7:0] n3394;
wire      [7:0] n3395;
wire      [7:0] n3396;
wire      [7:0] n3397;
wire      [7:0] n3398;
wire      [7:0] n3399;
wire            n34;
wire      [7:0] n340;
wire      [7:0] n3400;
wire    [103:0] n3401;
wire      [7:0] n3402;
wire      [7:0] n3403;
wire      [7:0] n3404;
wire      [7:0] n3405;
wire      [7:0] n3406;
wire      [7:0] n3407;
wire      [7:0] n3408;
wire      [7:0] n3409;
wire    [111:0] n3410;
wire      [7:0] n3411;
wire      [7:0] n3412;
wire      [7:0] n3413;
wire      [7:0] n3414;
wire      [7:0] n3415;
wire      [7:0] n3416;
wire      [7:0] n3417;
wire      [7:0] n3418;
wire    [119:0] n3419;
wire            n342;
wire      [7:0] n3420;
wire      [7:0] n3421;
wire      [7:0] n3422;
wire      [7:0] n3423;
wire      [7:0] n3424;
wire      [7:0] n3425;
wire      [7:0] n3426;
wire      [7:0] n3427;
wire    [127:0] n3428;
wire    [127:0] n3429;
wire      [7:0] n3430;
wire      [7:0] n3431;
wire      [7:0] n3432;
wire            n3433;
wire      [7:0] n3434;
wire            n3435;
wire      [7:0] n3436;
wire            n3437;
wire      [7:0] n3438;
wire            n3439;
wire      [7:0] n344;
wire      [7:0] n3440;
wire            n3441;
wire      [7:0] n3442;
wire            n3443;
wire      [7:0] n3444;
wire            n3445;
wire      [7:0] n3446;
wire            n3447;
wire      [7:0] n3448;
wire            n3449;
wire      [7:0] n3450;
wire            n3451;
wire      [7:0] n3452;
wire            n3453;
wire      [7:0] n3454;
wire            n3455;
wire      [7:0] n3456;
wire            n3457;
wire      [7:0] n3458;
wire            n3459;
wire            n346;
wire      [7:0] n3460;
wire            n3461;
wire      [7:0] n3462;
wire            n3463;
wire      [7:0] n3464;
wire            n3465;
wire      [7:0] n3466;
wire            n3467;
wire      [7:0] n3468;
wire            n3469;
wire      [7:0] n3470;
wire            n3471;
wire      [7:0] n3472;
wire            n3473;
wire      [7:0] n3474;
wire            n3475;
wire      [7:0] n3476;
wire            n3477;
wire      [7:0] n3478;
wire            n3479;
wire      [7:0] n348;
wire      [7:0] n3480;
wire            n3481;
wire      [7:0] n3482;
wire            n3483;
wire      [7:0] n3484;
wire            n3485;
wire      [7:0] n3486;
wire            n3487;
wire      [7:0] n3488;
wire            n3489;
wire            n349;
wire      [7:0] n3490;
wire            n3491;
wire      [7:0] n3492;
wire            n3493;
wire      [7:0] n3494;
wire            n3495;
wire      [7:0] n3496;
wire            n3497;
wire      [7:0] n3498;
wire            n3499;
wire      [7:0] n3500;
wire            n3501;
wire      [7:0] n3502;
wire            n3503;
wire      [7:0] n3504;
wire            n3505;
wire      [7:0] n3506;
wire            n3507;
wire      [7:0] n3508;
wire            n3509;
wire      [7:0] n351;
wire      [7:0] n3510;
wire            n3511;
wire      [7:0] n3512;
wire            n3513;
wire      [7:0] n3514;
wire            n3515;
wire      [7:0] n3516;
wire            n3517;
wire      [7:0] n3518;
wire            n3519;
wire      [7:0] n3520;
wire            n3521;
wire      [7:0] n3522;
wire            n3523;
wire      [7:0] n3524;
wire            n3525;
wire      [7:0] n3526;
wire            n3527;
wire      [7:0] n3528;
wire            n3529;
wire            n353;
wire      [7:0] n3530;
wire            n3531;
wire      [7:0] n3532;
wire            n3533;
wire      [7:0] n3534;
wire            n3535;
wire      [7:0] n3536;
wire            n3537;
wire      [7:0] n3538;
wire            n3539;
wire      [7:0] n354;
wire      [7:0] n3540;
wire            n3541;
wire      [7:0] n3542;
wire            n3543;
wire      [7:0] n3544;
wire            n3545;
wire      [7:0] n3546;
wire            n3547;
wire      [7:0] n3548;
wire            n3549;
wire      [7:0] n3550;
wire            n3551;
wire      [7:0] n3552;
wire            n3553;
wire      [7:0] n3554;
wire            n3555;
wire      [7:0] n3556;
wire            n3557;
wire      [7:0] n3558;
wire            n3559;
wire            n356;
wire      [7:0] n3560;
wire            n3561;
wire      [7:0] n3562;
wire            n3563;
wire      [7:0] n3564;
wire            n3565;
wire      [7:0] n3566;
wire            n3567;
wire      [7:0] n3568;
wire            n3569;
wire      [7:0] n357;
wire      [7:0] n3570;
wire            n3571;
wire      [7:0] n3572;
wire            n3573;
wire      [7:0] n3574;
wire            n3575;
wire      [7:0] n3576;
wire            n3577;
wire      [7:0] n3578;
wire            n3579;
wire            n358;
wire      [7:0] n3580;
wire            n3581;
wire      [7:0] n3582;
wire            n3583;
wire      [7:0] n3584;
wire            n3585;
wire      [7:0] n3586;
wire            n3587;
wire      [7:0] n3588;
wire            n3589;
wire      [7:0] n3590;
wire            n3591;
wire      [7:0] n3592;
wire            n3593;
wire      [7:0] n3594;
wire            n3595;
wire      [7:0] n3596;
wire            n3597;
wire      [7:0] n3598;
wire            n3599;
wire      [7:0] n36;
wire      [7:0] n360;
wire      [7:0] n3600;
wire            n3601;
wire      [7:0] n3602;
wire            n3603;
wire      [7:0] n3604;
wire            n3605;
wire      [7:0] n3606;
wire            n3607;
wire      [7:0] n3608;
wire            n3609;
wire      [7:0] n3610;
wire            n3611;
wire      [7:0] n3612;
wire            n3613;
wire      [7:0] n3614;
wire            n3615;
wire      [7:0] n3616;
wire            n3617;
wire      [7:0] n3618;
wire            n3619;
wire            n362;
wire      [7:0] n3620;
wire            n3621;
wire      [7:0] n3622;
wire            n3623;
wire      [7:0] n3624;
wire            n3625;
wire      [7:0] n3626;
wire            n3627;
wire      [7:0] n3628;
wire            n3629;
wire      [7:0] n3630;
wire            n3631;
wire      [7:0] n3632;
wire            n3633;
wire      [7:0] n3634;
wire            n3635;
wire      [7:0] n3636;
wire            n3637;
wire      [7:0] n3638;
wire            n3639;
wire      [7:0] n364;
wire      [7:0] n3640;
wire            n3641;
wire      [7:0] n3642;
wire            n3643;
wire      [7:0] n3644;
wire            n3645;
wire      [7:0] n3646;
wire            n3647;
wire      [7:0] n3648;
wire            n3649;
wire      [7:0] n3650;
wire            n3651;
wire      [7:0] n3652;
wire            n3653;
wire      [7:0] n3654;
wire            n3655;
wire      [7:0] n3656;
wire            n3657;
wire      [7:0] n3658;
wire            n3659;
wire            n366;
wire      [7:0] n3660;
wire            n3661;
wire      [7:0] n3662;
wire            n3663;
wire      [7:0] n3664;
wire            n3665;
wire      [7:0] n3666;
wire            n3667;
wire      [7:0] n3668;
wire            n3669;
wire      [7:0] n367;
wire      [7:0] n3670;
wire            n3671;
wire      [7:0] n3672;
wire            n3673;
wire      [7:0] n3674;
wire            n3675;
wire      [7:0] n3676;
wire            n3677;
wire      [7:0] n3678;
wire            n3679;
wire            n368;
wire      [7:0] n3680;
wire            n3681;
wire      [7:0] n3682;
wire            n3683;
wire      [7:0] n3684;
wire            n3685;
wire      [7:0] n3686;
wire            n3687;
wire      [7:0] n3688;
wire            n3689;
wire      [7:0] n3690;
wire            n3691;
wire      [7:0] n3692;
wire            n3693;
wire      [7:0] n3694;
wire            n3695;
wire      [7:0] n3696;
wire            n3697;
wire      [7:0] n3698;
wire            n3699;
wire      [7:0] n370;
wire      [7:0] n3700;
wire            n3701;
wire      [7:0] n3702;
wire            n3703;
wire      [7:0] n3704;
wire            n3705;
wire      [7:0] n3706;
wire            n3707;
wire      [7:0] n3708;
wire            n3709;
wire      [7:0] n3710;
wire            n3711;
wire      [7:0] n3712;
wire            n3713;
wire      [7:0] n3714;
wire            n3715;
wire      [7:0] n3716;
wire            n3717;
wire      [7:0] n3718;
wire            n3719;
wire            n372;
wire      [7:0] n3720;
wire            n3721;
wire      [7:0] n3722;
wire            n3723;
wire      [7:0] n3724;
wire            n3725;
wire      [7:0] n3726;
wire            n3727;
wire      [7:0] n3728;
wire            n3729;
wire      [7:0] n373;
wire      [7:0] n3730;
wire            n3731;
wire      [7:0] n3732;
wire            n3733;
wire      [7:0] n3734;
wire            n3735;
wire      [7:0] n3736;
wire            n3737;
wire      [7:0] n3738;
wire            n3739;
wire            n374;
wire      [7:0] n3740;
wire            n3741;
wire      [7:0] n3742;
wire            n3743;
wire      [7:0] n3744;
wire            n3745;
wire      [7:0] n3746;
wire            n3747;
wire      [7:0] n3748;
wire            n3749;
wire      [7:0] n375;
wire      [7:0] n3750;
wire            n3751;
wire      [7:0] n3752;
wire            n3753;
wire      [7:0] n3754;
wire            n3755;
wire      [7:0] n3756;
wire            n3757;
wire      [7:0] n3758;
wire            n3759;
wire            n376;
wire      [7:0] n3760;
wire            n3761;
wire      [7:0] n3762;
wire            n3763;
wire      [7:0] n3764;
wire            n3765;
wire      [7:0] n3766;
wire            n3767;
wire      [7:0] n3768;
wire            n3769;
wire      [7:0] n3770;
wire            n3771;
wire      [7:0] n3772;
wire            n3773;
wire      [7:0] n3774;
wire            n3775;
wire      [7:0] n3776;
wire            n3777;
wire      [7:0] n3778;
wire            n3779;
wire      [7:0] n378;
wire      [7:0] n3780;
wire            n3781;
wire      [7:0] n3782;
wire            n3783;
wire      [7:0] n3784;
wire            n3785;
wire      [7:0] n3786;
wire            n3787;
wire      [7:0] n3788;
wire            n3789;
wire      [7:0] n3790;
wire            n3791;
wire      [7:0] n3792;
wire            n3793;
wire      [7:0] n3794;
wire            n3795;
wire      [7:0] n3796;
wire            n3797;
wire      [7:0] n3798;
wire            n3799;
wire            n38;
wire            n380;
wire      [7:0] n3800;
wire            n3801;
wire      [7:0] n3802;
wire            n3803;
wire      [7:0] n3804;
wire            n3805;
wire      [7:0] n3806;
wire            n3807;
wire      [7:0] n3808;
wire            n3809;
wire      [7:0] n3810;
wire            n3811;
wire      [7:0] n3812;
wire            n3813;
wire      [7:0] n3814;
wire            n3815;
wire      [7:0] n3816;
wire            n3817;
wire      [7:0] n3818;
wire            n3819;
wire      [7:0] n382;
wire      [7:0] n3820;
wire            n3821;
wire      [7:0] n3822;
wire            n3823;
wire      [7:0] n3824;
wire            n3825;
wire      [7:0] n3826;
wire            n3827;
wire      [7:0] n3828;
wire            n3829;
wire      [7:0] n3830;
wire            n3831;
wire      [7:0] n3832;
wire            n3833;
wire      [7:0] n3834;
wire            n3835;
wire      [7:0] n3836;
wire            n3837;
wire      [7:0] n3838;
wire            n3839;
wire            n384;
wire      [7:0] n3840;
wire            n3841;
wire      [7:0] n3842;
wire            n3843;
wire      [7:0] n3844;
wire            n3845;
wire      [7:0] n3846;
wire            n3847;
wire      [7:0] n3848;
wire            n3849;
wire      [7:0] n3850;
wire            n3851;
wire      [7:0] n3852;
wire            n3853;
wire      [7:0] n3854;
wire            n3855;
wire      [7:0] n3856;
wire            n3857;
wire      [7:0] n3858;
wire            n3859;
wire      [7:0] n386;
wire      [7:0] n3860;
wire            n3861;
wire      [7:0] n3862;
wire            n3863;
wire      [7:0] n3864;
wire            n3865;
wire      [7:0] n3866;
wire            n3867;
wire      [7:0] n3868;
wire            n3869;
wire            n387;
wire      [7:0] n3870;
wire            n3871;
wire      [7:0] n3872;
wire            n3873;
wire      [7:0] n3874;
wire            n3875;
wire      [7:0] n3876;
wire            n3877;
wire      [7:0] n3878;
wire            n3879;
wire      [7:0] n3880;
wire            n3881;
wire      [7:0] n3882;
wire            n3883;
wire      [7:0] n3884;
wire            n3885;
wire      [7:0] n3886;
wire            n3887;
wire      [7:0] n3888;
wire            n3889;
wire      [7:0] n389;
wire      [7:0] n3890;
wire            n3891;
wire      [7:0] n3892;
wire            n3893;
wire      [7:0] n3894;
wire            n3895;
wire      [7:0] n3896;
wire            n3897;
wire      [7:0] n3898;
wire            n3899;
wire            n390;
wire      [7:0] n3900;
wire            n3901;
wire      [7:0] n3902;
wire            n3903;
wire      [7:0] n3904;
wire            n3905;
wire      [7:0] n3906;
wire            n3907;
wire      [7:0] n3908;
wire            n3909;
wire      [7:0] n3910;
wire            n3911;
wire      [7:0] n3912;
wire            n3913;
wire      [7:0] n3914;
wire            n3915;
wire      [7:0] n3916;
wire            n3917;
wire      [7:0] n3918;
wire            n3919;
wire      [7:0] n392;
wire      [7:0] n3920;
wire            n3921;
wire      [7:0] n3922;
wire            n3923;
wire      [7:0] n3924;
wire            n3925;
wire      [7:0] n3926;
wire            n3927;
wire      [7:0] n3928;
wire            n3929;
wire      [7:0] n3930;
wire            n3931;
wire      [7:0] n3932;
wire            n3933;
wire      [7:0] n3934;
wire            n3935;
wire      [7:0] n3936;
wire            n3937;
wire      [7:0] n3938;
wire            n3939;
wire            n394;
wire      [7:0] n3940;
wire            n3941;
wire      [7:0] n3942;
wire            n3943;
wire      [7:0] n3944;
wire      [7:0] n3945;
wire      [7:0] n3946;
wire      [7:0] n3947;
wire      [7:0] n3948;
wire      [7:0] n3949;
wire      [7:0] n395;
wire      [7:0] n3950;
wire      [7:0] n3951;
wire      [7:0] n3952;
wire      [7:0] n3953;
wire      [7:0] n3954;
wire      [7:0] n3955;
wire      [7:0] n3956;
wire      [7:0] n3957;
wire      [7:0] n3958;
wire      [7:0] n3959;
wire      [7:0] n3960;
wire      [7:0] n3961;
wire      [7:0] n3962;
wire      [7:0] n3963;
wire      [7:0] n3964;
wire      [7:0] n3965;
wire      [7:0] n3966;
wire      [7:0] n3967;
wire      [7:0] n3968;
wire      [7:0] n3969;
wire            n397;
wire      [7:0] n3970;
wire      [7:0] n3971;
wire      [7:0] n3972;
wire      [7:0] n3973;
wire      [7:0] n3974;
wire      [7:0] n3975;
wire      [7:0] n3976;
wire      [7:0] n3977;
wire      [7:0] n3978;
wire      [7:0] n3979;
wire      [7:0] n3980;
wire      [7:0] n3981;
wire      [7:0] n3982;
wire      [7:0] n3983;
wire      [7:0] n3984;
wire      [7:0] n3985;
wire      [7:0] n3986;
wire      [7:0] n3987;
wire      [7:0] n3988;
wire      [7:0] n3989;
wire      [7:0] n399;
wire      [7:0] n3990;
wire      [7:0] n3991;
wire      [7:0] n3992;
wire      [7:0] n3993;
wire      [7:0] n3994;
wire      [7:0] n3995;
wire      [7:0] n3996;
wire      [7:0] n3997;
wire      [7:0] n3998;
wire      [7:0] n3999;
wire      [7:0] n4;
wire      [7:0] n40;
wire            n400;
wire      [7:0] n4000;
wire      [7:0] n4001;
wire      [7:0] n4002;
wire      [7:0] n4003;
wire      [7:0] n4004;
wire      [7:0] n4005;
wire      [7:0] n4006;
wire      [7:0] n4007;
wire      [7:0] n4008;
wire      [7:0] n4009;
wire      [7:0] n4010;
wire      [7:0] n4011;
wire      [7:0] n4012;
wire      [7:0] n4013;
wire      [7:0] n4014;
wire      [7:0] n4015;
wire      [7:0] n4016;
wire      [7:0] n4017;
wire      [7:0] n4018;
wire      [7:0] n4019;
wire      [7:0] n402;
wire      [7:0] n4020;
wire      [7:0] n4021;
wire      [7:0] n4022;
wire      [7:0] n4023;
wire      [7:0] n4024;
wire      [7:0] n4025;
wire      [7:0] n4026;
wire      [7:0] n4027;
wire      [7:0] n4028;
wire      [7:0] n4029;
wire            n403;
wire      [7:0] n4030;
wire      [7:0] n4031;
wire      [7:0] n4032;
wire      [7:0] n4033;
wire      [7:0] n4034;
wire      [7:0] n4035;
wire      [7:0] n4036;
wire      [7:0] n4037;
wire      [7:0] n4038;
wire      [7:0] n4039;
wire      [7:0] n4040;
wire      [7:0] n4041;
wire      [7:0] n4042;
wire      [7:0] n4043;
wire      [7:0] n4044;
wire      [7:0] n4045;
wire      [7:0] n4046;
wire      [7:0] n4047;
wire      [7:0] n4048;
wire      [7:0] n4049;
wire      [7:0] n405;
wire      [7:0] n4050;
wire      [7:0] n4051;
wire      [7:0] n4052;
wire      [7:0] n4053;
wire      [7:0] n4054;
wire      [7:0] n4055;
wire      [7:0] n4056;
wire      [7:0] n4057;
wire      [7:0] n4058;
wire      [7:0] n4059;
wire      [7:0] n4060;
wire      [7:0] n4061;
wire      [7:0] n4062;
wire      [7:0] n4063;
wire      [7:0] n4064;
wire      [7:0] n4065;
wire      [7:0] n4066;
wire      [7:0] n4067;
wire      [7:0] n4068;
wire      [7:0] n4069;
wire            n407;
wire      [7:0] n4070;
wire      [7:0] n4071;
wire      [7:0] n4072;
wire      [7:0] n4073;
wire      [7:0] n4074;
wire      [7:0] n4075;
wire      [7:0] n4076;
wire      [7:0] n4077;
wire      [7:0] n4078;
wire      [7:0] n4079;
wire      [7:0] n4080;
wire      [7:0] n4081;
wire      [7:0] n4082;
wire      [7:0] n4083;
wire      [7:0] n4084;
wire      [7:0] n4085;
wire      [7:0] n4086;
wire      [7:0] n4087;
wire      [7:0] n4088;
wire      [7:0] n4089;
wire      [7:0] n409;
wire      [7:0] n4090;
wire      [7:0] n4091;
wire      [7:0] n4092;
wire      [7:0] n4093;
wire      [7:0] n4094;
wire      [7:0] n4095;
wire      [7:0] n4096;
wire      [7:0] n4097;
wire      [7:0] n4098;
wire      [7:0] n4099;
wire            n410;
wire      [7:0] n4100;
wire      [7:0] n4101;
wire      [7:0] n4102;
wire      [7:0] n4103;
wire      [7:0] n4104;
wire      [7:0] n4105;
wire      [7:0] n4106;
wire      [7:0] n4107;
wire      [7:0] n4108;
wire      [7:0] n4109;
wire      [7:0] n4110;
wire      [7:0] n4111;
wire      [7:0] n4112;
wire      [7:0] n4113;
wire      [7:0] n4114;
wire      [7:0] n4115;
wire      [7:0] n4116;
wire      [7:0] n4117;
wire      [7:0] n4118;
wire      [7:0] n4119;
wire      [7:0] n412;
wire      [7:0] n4120;
wire      [7:0] n4121;
wire      [7:0] n4122;
wire      [7:0] n4123;
wire      [7:0] n4124;
wire      [7:0] n4125;
wire      [7:0] n4126;
wire      [7:0] n4127;
wire      [7:0] n4128;
wire      [7:0] n4129;
wire            n413;
wire      [7:0] n4130;
wire      [7:0] n4131;
wire      [7:0] n4132;
wire      [7:0] n4133;
wire      [7:0] n4134;
wire      [7:0] n4135;
wire      [7:0] n4136;
wire      [7:0] n4137;
wire      [7:0] n4138;
wire      [7:0] n4139;
wire      [7:0] n4140;
wire      [7:0] n4141;
wire      [7:0] n4142;
wire      [7:0] n4143;
wire      [7:0] n4144;
wire      [7:0] n4145;
wire      [7:0] n4146;
wire      [7:0] n4147;
wire      [7:0] n4148;
wire      [7:0] n4149;
wire      [7:0] n415;
wire      [7:0] n4150;
wire      [7:0] n4151;
wire      [7:0] n4152;
wire      [7:0] n4153;
wire      [7:0] n4154;
wire      [7:0] n4155;
wire      [7:0] n4156;
wire      [7:0] n4157;
wire      [7:0] n4158;
wire      [7:0] n4159;
wire            n416;
wire      [7:0] n4160;
wire      [7:0] n4161;
wire      [7:0] n4162;
wire      [7:0] n4163;
wire      [7:0] n4164;
wire      [7:0] n4165;
wire      [7:0] n4166;
wire      [7:0] n4167;
wire      [7:0] n4168;
wire      [7:0] n4169;
wire      [7:0] n4170;
wire      [7:0] n4171;
wire      [7:0] n4172;
wire      [7:0] n4173;
wire      [7:0] n4174;
wire      [7:0] n4175;
wire      [7:0] n4176;
wire      [7:0] n4177;
wire      [7:0] n4178;
wire      [7:0] n4179;
wire      [7:0] n418;
wire      [7:0] n4180;
wire      [7:0] n4181;
wire      [7:0] n4182;
wire      [7:0] n4183;
wire      [7:0] n4184;
wire      [7:0] n4185;
wire      [7:0] n4186;
wire      [7:0] n4187;
wire      [7:0] n4188;
wire      [7:0] n4189;
wire            n419;
wire      [7:0] n4190;
wire      [7:0] n4191;
wire      [7:0] n4192;
wire      [7:0] n4193;
wire      [7:0] n4194;
wire      [7:0] n4195;
wire      [7:0] n4196;
wire      [7:0] n4197;
wire      [7:0] n4198;
wire      [7:0] n4199;
wire            n42;
wire      [7:0] n4200;
wire      [7:0] n4201;
wire      [7:0] n4202;
wire            n4203;
wire      [7:0] n4204;
wire            n4205;
wire      [7:0] n4206;
wire            n4207;
wire      [7:0] n4208;
wire            n4209;
wire      [7:0] n421;
wire      [7:0] n4210;
wire            n4211;
wire      [7:0] n4212;
wire            n4213;
wire      [7:0] n4214;
wire            n4215;
wire      [7:0] n4216;
wire            n4217;
wire      [7:0] n4218;
wire            n4219;
wire            n422;
wire      [7:0] n4220;
wire            n4221;
wire      [7:0] n4222;
wire            n4223;
wire      [7:0] n4224;
wire            n4225;
wire      [7:0] n4226;
wire            n4227;
wire      [7:0] n4228;
wire            n4229;
wire      [7:0] n4230;
wire            n4231;
wire      [7:0] n4232;
wire            n4233;
wire      [7:0] n4234;
wire            n4235;
wire      [7:0] n4236;
wire            n4237;
wire      [7:0] n4238;
wire            n4239;
wire      [7:0] n424;
wire      [7:0] n4240;
wire            n4241;
wire      [7:0] n4242;
wire            n4243;
wire      [7:0] n4244;
wire            n4245;
wire      [7:0] n4246;
wire            n4247;
wire      [7:0] n4248;
wire            n4249;
wire            n425;
wire      [7:0] n4250;
wire            n4251;
wire      [7:0] n4252;
wire            n4253;
wire      [7:0] n4254;
wire            n4255;
wire      [7:0] n4256;
wire            n4257;
wire      [7:0] n4258;
wire            n4259;
wire      [7:0] n426;
wire      [7:0] n4260;
wire            n4261;
wire      [7:0] n4262;
wire            n4263;
wire      [7:0] n4264;
wire            n4265;
wire      [7:0] n4266;
wire            n4267;
wire      [7:0] n4268;
wire            n4269;
wire            n427;
wire      [7:0] n4270;
wire            n4271;
wire      [7:0] n4272;
wire            n4273;
wire      [7:0] n4274;
wire            n4275;
wire      [7:0] n4276;
wire            n4277;
wire      [7:0] n4278;
wire            n4279;
wire      [7:0] n428;
wire      [7:0] n4280;
wire            n4281;
wire      [7:0] n4282;
wire            n4283;
wire      [7:0] n4284;
wire            n4285;
wire      [7:0] n4286;
wire            n4287;
wire      [7:0] n4288;
wire            n4289;
wire            n429;
wire      [7:0] n4290;
wire            n4291;
wire      [7:0] n4292;
wire            n4293;
wire      [7:0] n4294;
wire            n4295;
wire      [7:0] n4296;
wire            n4297;
wire      [7:0] n4298;
wire            n4299;
wire      [7:0] n4300;
wire            n4301;
wire      [7:0] n4302;
wire            n4303;
wire      [7:0] n4304;
wire            n4305;
wire      [7:0] n4306;
wire            n4307;
wire      [7:0] n4308;
wire            n4309;
wire      [7:0] n431;
wire      [7:0] n4310;
wire            n4311;
wire      [7:0] n4312;
wire            n4313;
wire      [7:0] n4314;
wire            n4315;
wire      [7:0] n4316;
wire            n4317;
wire      [7:0] n4318;
wire            n4319;
wire            n432;
wire      [7:0] n4320;
wire            n4321;
wire      [7:0] n4322;
wire            n4323;
wire      [7:0] n4324;
wire            n4325;
wire      [7:0] n4326;
wire            n4327;
wire      [7:0] n4328;
wire            n4329;
wire      [7:0] n4330;
wire            n4331;
wire      [7:0] n4332;
wire            n4333;
wire      [7:0] n4334;
wire            n4335;
wire      [7:0] n4336;
wire            n4337;
wire      [7:0] n4338;
wire            n4339;
wire      [7:0] n434;
wire      [7:0] n4340;
wire            n4341;
wire      [7:0] n4342;
wire            n4343;
wire      [7:0] n4344;
wire            n4345;
wire      [7:0] n4346;
wire            n4347;
wire      [7:0] n4348;
wire            n4349;
wire      [7:0] n4350;
wire            n4351;
wire      [7:0] n4352;
wire            n4353;
wire      [7:0] n4354;
wire            n4355;
wire      [7:0] n4356;
wire            n4357;
wire      [7:0] n4358;
wire            n4359;
wire            n436;
wire      [7:0] n4360;
wire            n4361;
wire      [7:0] n4362;
wire            n4363;
wire      [7:0] n4364;
wire            n4365;
wire      [7:0] n4366;
wire            n4367;
wire      [7:0] n4368;
wire            n4369;
wire      [7:0] n437;
wire      [7:0] n4370;
wire            n4371;
wire      [7:0] n4372;
wire            n4373;
wire      [7:0] n4374;
wire            n4375;
wire      [7:0] n4376;
wire            n4377;
wire      [7:0] n4378;
wire            n4379;
wire      [7:0] n4380;
wire            n4381;
wire      [7:0] n4382;
wire            n4383;
wire      [7:0] n4384;
wire            n4385;
wire      [7:0] n4386;
wire            n4387;
wire      [7:0] n4388;
wire            n4389;
wire            n439;
wire      [7:0] n4390;
wire            n4391;
wire      [7:0] n4392;
wire            n4393;
wire      [7:0] n4394;
wire            n4395;
wire      [7:0] n4396;
wire            n4397;
wire      [7:0] n4398;
wire            n4399;
wire      [7:0] n44;
wire      [7:0] n4400;
wire            n4401;
wire      [7:0] n4402;
wire            n4403;
wire      [7:0] n4404;
wire            n4405;
wire      [7:0] n4406;
wire            n4407;
wire      [7:0] n4408;
wire            n4409;
wire      [7:0] n441;
wire      [7:0] n4410;
wire            n4411;
wire      [7:0] n4412;
wire            n4413;
wire      [7:0] n4414;
wire            n4415;
wire      [7:0] n4416;
wire            n4417;
wire      [7:0] n4418;
wire            n4419;
wire      [7:0] n4420;
wire            n4421;
wire      [7:0] n4422;
wire            n4423;
wire      [7:0] n4424;
wire            n4425;
wire      [7:0] n4426;
wire            n4427;
wire      [7:0] n4428;
wire            n4429;
wire            n443;
wire      [7:0] n4430;
wire            n4431;
wire      [7:0] n4432;
wire            n4433;
wire      [7:0] n4434;
wire            n4435;
wire      [7:0] n4436;
wire            n4437;
wire      [7:0] n4438;
wire            n4439;
wire      [7:0] n444;
wire      [7:0] n4440;
wire            n4441;
wire      [7:0] n4442;
wire            n4443;
wire      [7:0] n4444;
wire            n4445;
wire      [7:0] n4446;
wire            n4447;
wire      [7:0] n4448;
wire            n4449;
wire      [7:0] n4450;
wire            n4451;
wire      [7:0] n4452;
wire            n4453;
wire      [7:0] n4454;
wire            n4455;
wire      [7:0] n4456;
wire            n4457;
wire      [7:0] n4458;
wire            n4459;
wire            n446;
wire      [7:0] n4460;
wire            n4461;
wire      [7:0] n4462;
wire            n4463;
wire      [7:0] n4464;
wire            n4465;
wire      [7:0] n4466;
wire            n4467;
wire      [7:0] n4468;
wire            n4469;
wire      [7:0] n4470;
wire            n4471;
wire      [7:0] n4472;
wire            n4473;
wire      [7:0] n4474;
wire            n4475;
wire      [7:0] n4476;
wire            n4477;
wire      [7:0] n4478;
wire            n4479;
wire      [7:0] n448;
wire      [7:0] n4480;
wire            n4481;
wire      [7:0] n4482;
wire            n4483;
wire      [7:0] n4484;
wire            n4485;
wire      [7:0] n4486;
wire            n4487;
wire      [7:0] n4488;
wire            n4489;
wire            n449;
wire      [7:0] n4490;
wire            n4491;
wire      [7:0] n4492;
wire            n4493;
wire      [7:0] n4494;
wire            n4495;
wire      [7:0] n4496;
wire            n4497;
wire      [7:0] n4498;
wire            n4499;
wire      [7:0] n4500;
wire            n4501;
wire      [7:0] n4502;
wire            n4503;
wire      [7:0] n4504;
wire            n4505;
wire      [7:0] n4506;
wire            n4507;
wire      [7:0] n4508;
wire            n4509;
wire      [7:0] n451;
wire      [7:0] n4510;
wire            n4511;
wire      [7:0] n4512;
wire            n4513;
wire      [7:0] n4514;
wire            n4515;
wire      [7:0] n4516;
wire            n4517;
wire      [7:0] n4518;
wire            n4519;
wire      [7:0] n4520;
wire            n4521;
wire      [7:0] n4522;
wire            n4523;
wire      [7:0] n4524;
wire            n4525;
wire      [7:0] n4526;
wire            n4527;
wire      [7:0] n4528;
wire            n4529;
wire            n453;
wire      [7:0] n4530;
wire            n4531;
wire      [7:0] n4532;
wire            n4533;
wire      [7:0] n4534;
wire            n4535;
wire      [7:0] n4536;
wire            n4537;
wire      [7:0] n4538;
wire            n4539;
wire      [7:0] n454;
wire      [7:0] n4540;
wire            n4541;
wire      [7:0] n4542;
wire            n4543;
wire      [7:0] n4544;
wire            n4545;
wire      [7:0] n4546;
wire            n4547;
wire      [7:0] n4548;
wire            n4549;
wire      [7:0] n4550;
wire            n4551;
wire      [7:0] n4552;
wire            n4553;
wire      [7:0] n4554;
wire            n4555;
wire      [7:0] n4556;
wire            n4557;
wire      [7:0] n4558;
wire            n4559;
wire            n456;
wire      [7:0] n4560;
wire            n4561;
wire      [7:0] n4562;
wire            n4563;
wire      [7:0] n4564;
wire            n4565;
wire      [7:0] n4566;
wire            n4567;
wire      [7:0] n4568;
wire            n4569;
wire      [7:0] n457;
wire      [7:0] n4570;
wire            n4571;
wire      [7:0] n4572;
wire            n4573;
wire      [7:0] n4574;
wire            n4575;
wire      [7:0] n4576;
wire            n4577;
wire      [7:0] n4578;
wire            n4579;
wire            n458;
wire      [7:0] n4580;
wire            n4581;
wire      [7:0] n4582;
wire            n4583;
wire      [7:0] n4584;
wire            n4585;
wire      [7:0] n4586;
wire            n4587;
wire      [7:0] n4588;
wire            n4589;
wire      [7:0] n459;
wire      [7:0] n4590;
wire            n4591;
wire      [7:0] n4592;
wire            n4593;
wire      [7:0] n4594;
wire            n4595;
wire      [7:0] n4596;
wire            n4597;
wire      [7:0] n4598;
wire            n4599;
wire            n46;
wire      [7:0] n4600;
wire            n4601;
wire      [7:0] n4602;
wire            n4603;
wire      [7:0] n4604;
wire            n4605;
wire      [7:0] n4606;
wire            n4607;
wire      [7:0] n4608;
wire            n4609;
wire            n461;
wire      [7:0] n4610;
wire            n4611;
wire      [7:0] n4612;
wire            n4613;
wire      [7:0] n4614;
wire            n4615;
wire      [7:0] n4616;
wire            n4617;
wire      [7:0] n4618;
wire            n4619;
wire      [7:0] n462;
wire      [7:0] n4620;
wire            n4621;
wire      [7:0] n4622;
wire            n4623;
wire      [7:0] n4624;
wire            n4625;
wire      [7:0] n4626;
wire            n4627;
wire      [7:0] n4628;
wire            n4629;
wire      [7:0] n4630;
wire            n4631;
wire      [7:0] n4632;
wire            n4633;
wire      [7:0] n4634;
wire            n4635;
wire      [7:0] n4636;
wire            n4637;
wire      [7:0] n4638;
wire            n4639;
wire            n464;
wire      [7:0] n4640;
wire            n4641;
wire      [7:0] n4642;
wire            n4643;
wire      [7:0] n4644;
wire            n4645;
wire      [7:0] n4646;
wire            n4647;
wire      [7:0] n4648;
wire            n4649;
wire      [7:0] n4650;
wire            n4651;
wire      [7:0] n4652;
wire            n4653;
wire      [7:0] n4654;
wire            n4655;
wire      [7:0] n4656;
wire            n4657;
wire      [7:0] n4658;
wire            n4659;
wire      [7:0] n466;
wire      [7:0] n4660;
wire            n4661;
wire      [7:0] n4662;
wire            n4663;
wire      [7:0] n4664;
wire            n4665;
wire      [7:0] n4666;
wire            n4667;
wire      [7:0] n4668;
wire            n4669;
wire      [7:0] n4670;
wire            n4671;
wire      [7:0] n4672;
wire            n4673;
wire      [7:0] n4674;
wire            n4675;
wire      [7:0] n4676;
wire            n4677;
wire      [7:0] n4678;
wire            n4679;
wire            n468;
wire      [7:0] n4680;
wire            n4681;
wire      [7:0] n4682;
wire            n4683;
wire      [7:0] n4684;
wire            n4685;
wire      [7:0] n4686;
wire            n4687;
wire      [7:0] n4688;
wire            n4689;
wire      [7:0] n4690;
wire            n4691;
wire      [7:0] n4692;
wire            n4693;
wire      [7:0] n4694;
wire            n4695;
wire      [7:0] n4696;
wire            n4697;
wire      [7:0] n4698;
wire            n4699;
wire      [7:0] n470;
wire      [7:0] n4700;
wire            n4701;
wire      [7:0] n4702;
wire            n4703;
wire      [7:0] n4704;
wire            n4705;
wire      [7:0] n4706;
wire            n4707;
wire      [7:0] n4708;
wire            n4709;
wire            n471;
wire      [7:0] n4710;
wire            n4711;
wire      [7:0] n4712;
wire            n4713;
wire      [7:0] n4714;
wire      [7:0] n4715;
wire      [7:0] n4716;
wire      [7:0] n4717;
wire      [7:0] n4718;
wire      [7:0] n4719;
wire      [7:0] n472;
wire      [7:0] n4720;
wire      [7:0] n4721;
wire      [7:0] n4722;
wire      [7:0] n4723;
wire      [7:0] n4724;
wire      [7:0] n4725;
wire      [7:0] n4726;
wire      [7:0] n4727;
wire      [7:0] n4728;
wire      [7:0] n4729;
wire            n473;
wire      [7:0] n4730;
wire      [7:0] n4731;
wire      [7:0] n4732;
wire      [7:0] n4733;
wire      [7:0] n4734;
wire      [7:0] n4735;
wire      [7:0] n4736;
wire      [7:0] n4737;
wire      [7:0] n4738;
wire      [7:0] n4739;
wire      [7:0] n474;
wire      [7:0] n4740;
wire      [7:0] n4741;
wire      [7:0] n4742;
wire      [7:0] n4743;
wire      [7:0] n4744;
wire      [7:0] n4745;
wire      [7:0] n4746;
wire      [7:0] n4747;
wire      [7:0] n4748;
wire      [7:0] n4749;
wire            n475;
wire      [7:0] n4750;
wire      [7:0] n4751;
wire      [7:0] n4752;
wire      [7:0] n4753;
wire      [7:0] n4754;
wire      [7:0] n4755;
wire      [7:0] n4756;
wire      [7:0] n4757;
wire      [7:0] n4758;
wire      [7:0] n4759;
wire      [7:0] n476;
wire      [7:0] n4760;
wire      [7:0] n4761;
wire      [7:0] n4762;
wire      [7:0] n4763;
wire      [7:0] n4764;
wire      [7:0] n4765;
wire      [7:0] n4766;
wire      [7:0] n4767;
wire      [7:0] n4768;
wire      [7:0] n4769;
wire      [7:0] n4770;
wire      [7:0] n4771;
wire      [7:0] n4772;
wire      [7:0] n4773;
wire      [7:0] n4774;
wire      [7:0] n4775;
wire      [7:0] n4776;
wire      [7:0] n4777;
wire      [7:0] n4778;
wire      [7:0] n4779;
wire            n478;
wire      [7:0] n4780;
wire      [7:0] n4781;
wire      [7:0] n4782;
wire      [7:0] n4783;
wire      [7:0] n4784;
wire      [7:0] n4785;
wire      [7:0] n4786;
wire      [7:0] n4787;
wire      [7:0] n4788;
wire      [7:0] n4789;
wire      [7:0] n479;
wire      [7:0] n4790;
wire      [7:0] n4791;
wire      [7:0] n4792;
wire      [7:0] n4793;
wire      [7:0] n4794;
wire      [7:0] n4795;
wire      [7:0] n4796;
wire      [7:0] n4797;
wire      [7:0] n4798;
wire      [7:0] n4799;
wire      [7:0] n48;
wire      [7:0] n4800;
wire      [7:0] n4801;
wire      [7:0] n4802;
wire      [7:0] n4803;
wire      [7:0] n4804;
wire      [7:0] n4805;
wire      [7:0] n4806;
wire      [7:0] n4807;
wire      [7:0] n4808;
wire      [7:0] n4809;
wire            n481;
wire      [7:0] n4810;
wire      [7:0] n4811;
wire      [7:0] n4812;
wire      [7:0] n4813;
wire      [7:0] n4814;
wire      [7:0] n4815;
wire      [7:0] n4816;
wire      [7:0] n4817;
wire      [7:0] n4818;
wire      [7:0] n4819;
wire      [7:0] n4820;
wire      [7:0] n4821;
wire      [7:0] n4822;
wire      [7:0] n4823;
wire      [7:0] n4824;
wire      [7:0] n4825;
wire      [7:0] n4826;
wire      [7:0] n4827;
wire      [7:0] n4828;
wire      [7:0] n4829;
wire      [7:0] n483;
wire      [7:0] n4830;
wire      [7:0] n4831;
wire      [7:0] n4832;
wire      [7:0] n4833;
wire      [7:0] n4834;
wire      [7:0] n4835;
wire      [7:0] n4836;
wire      [7:0] n4837;
wire      [7:0] n4838;
wire      [7:0] n4839;
wire      [7:0] n4840;
wire      [7:0] n4841;
wire      [7:0] n4842;
wire      [7:0] n4843;
wire      [7:0] n4844;
wire      [7:0] n4845;
wire      [7:0] n4846;
wire      [7:0] n4847;
wire      [7:0] n4848;
wire      [7:0] n4849;
wire            n485;
wire      [7:0] n4850;
wire      [7:0] n4851;
wire      [7:0] n4852;
wire      [7:0] n4853;
wire      [7:0] n4854;
wire      [7:0] n4855;
wire      [7:0] n4856;
wire      [7:0] n4857;
wire      [7:0] n4858;
wire      [7:0] n4859;
wire      [7:0] n486;
wire      [7:0] n4860;
wire      [7:0] n4861;
wire      [7:0] n4862;
wire      [7:0] n4863;
wire      [7:0] n4864;
wire      [7:0] n4865;
wire      [7:0] n4866;
wire      [7:0] n4867;
wire      [7:0] n4868;
wire      [7:0] n4869;
wire            n487;
wire      [7:0] n4870;
wire      [7:0] n4871;
wire      [7:0] n4872;
wire      [7:0] n4873;
wire      [7:0] n4874;
wire      [7:0] n4875;
wire      [7:0] n4876;
wire      [7:0] n4877;
wire      [7:0] n4878;
wire      [7:0] n4879;
wire      [7:0] n488;
wire      [7:0] n4880;
wire      [7:0] n4881;
wire      [7:0] n4882;
wire      [7:0] n4883;
wire      [7:0] n4884;
wire      [7:0] n4885;
wire      [7:0] n4886;
wire      [7:0] n4887;
wire      [7:0] n4888;
wire      [7:0] n4889;
wire            n489;
wire      [7:0] n4890;
wire      [7:0] n4891;
wire      [7:0] n4892;
wire      [7:0] n4893;
wire      [7:0] n4894;
wire      [7:0] n4895;
wire      [7:0] n4896;
wire      [7:0] n4897;
wire      [7:0] n4898;
wire      [7:0] n4899;
wire      [7:0] n490;
wire      [7:0] n4900;
wire      [7:0] n4901;
wire      [7:0] n4902;
wire      [7:0] n4903;
wire      [7:0] n4904;
wire      [7:0] n4905;
wire      [7:0] n4906;
wire      [7:0] n4907;
wire      [7:0] n4908;
wire      [7:0] n4909;
wire      [7:0] n4910;
wire      [7:0] n4911;
wire      [7:0] n4912;
wire      [7:0] n4913;
wire      [7:0] n4914;
wire      [7:0] n4915;
wire      [7:0] n4916;
wire      [7:0] n4917;
wire      [7:0] n4918;
wire      [7:0] n4919;
wire            n492;
wire      [7:0] n4920;
wire      [7:0] n4921;
wire      [7:0] n4922;
wire      [7:0] n4923;
wire      [7:0] n4924;
wire      [7:0] n4925;
wire      [7:0] n4926;
wire      [7:0] n4927;
wire      [7:0] n4928;
wire      [7:0] n4929;
wire      [7:0] n4930;
wire      [7:0] n4931;
wire      [7:0] n4932;
wire      [7:0] n4933;
wire      [7:0] n4934;
wire      [7:0] n4935;
wire      [7:0] n4936;
wire      [7:0] n4937;
wire      [7:0] n4938;
wire      [7:0] n4939;
wire      [7:0] n494;
wire      [7:0] n4940;
wire      [7:0] n4941;
wire      [7:0] n4942;
wire      [7:0] n4943;
wire      [7:0] n4944;
wire      [7:0] n4945;
wire      [7:0] n4946;
wire      [7:0] n4947;
wire      [7:0] n4948;
wire      [7:0] n4949;
wire      [7:0] n4950;
wire      [7:0] n4951;
wire      [7:0] n4952;
wire      [7:0] n4953;
wire      [7:0] n4954;
wire      [7:0] n4955;
wire      [7:0] n4956;
wire      [7:0] n4957;
wire      [7:0] n4958;
wire      [7:0] n4959;
wire            n496;
wire      [7:0] n4960;
wire      [7:0] n4961;
wire      [7:0] n4962;
wire      [7:0] n4963;
wire      [7:0] n4964;
wire      [7:0] n4965;
wire      [7:0] n4966;
wire      [7:0] n4967;
wire      [7:0] n4968;
wire      [7:0] n4969;
wire      [7:0] n497;
wire      [7:0] n4970;
wire     [15:0] n4971;
wire      [7:0] n4972;
wire      [7:0] n4973;
wire            n4974;
wire      [7:0] n4975;
wire            n4976;
wire      [7:0] n4977;
wire            n4978;
wire      [7:0] n4979;
wire            n498;
wire            n4980;
wire      [7:0] n4981;
wire            n4982;
wire      [7:0] n4983;
wire            n4984;
wire      [7:0] n4985;
wire            n4986;
wire      [7:0] n4987;
wire            n4988;
wire      [7:0] n4989;
wire            n4990;
wire      [7:0] n4991;
wire            n4992;
wire      [7:0] n4993;
wire            n4994;
wire      [7:0] n4995;
wire            n4996;
wire      [7:0] n4997;
wire            n4998;
wire      [7:0] n4999;
wire            n50;
wire      [7:0] n500;
wire            n5000;
wire      [7:0] n5001;
wire            n5002;
wire      [7:0] n5003;
wire            n5004;
wire      [7:0] n5005;
wire            n5006;
wire      [7:0] n5007;
wire            n5008;
wire      [7:0] n5009;
wire            n5010;
wire      [7:0] n5011;
wire            n5012;
wire      [7:0] n5013;
wire            n5014;
wire      [7:0] n5015;
wire            n5016;
wire      [7:0] n5017;
wire            n5018;
wire      [7:0] n5019;
wire            n502;
wire            n5020;
wire      [7:0] n5021;
wire            n5022;
wire      [7:0] n5023;
wire            n5024;
wire      [7:0] n5025;
wire            n5026;
wire      [7:0] n5027;
wire            n5028;
wire      [7:0] n5029;
wire      [7:0] n503;
wire            n5030;
wire      [7:0] n5031;
wire            n5032;
wire      [7:0] n5033;
wire            n5034;
wire      [7:0] n5035;
wire            n5036;
wire      [7:0] n5037;
wire            n5038;
wire      [7:0] n5039;
wire            n5040;
wire      [7:0] n5041;
wire            n5042;
wire      [7:0] n5043;
wire            n5044;
wire      [7:0] n5045;
wire            n5046;
wire      [7:0] n5047;
wire            n5048;
wire      [7:0] n5049;
wire            n505;
wire            n5050;
wire      [7:0] n5051;
wire            n5052;
wire      [7:0] n5053;
wire            n5054;
wire      [7:0] n5055;
wire            n5056;
wire      [7:0] n5057;
wire            n5058;
wire      [7:0] n5059;
wire      [7:0] n506;
wire            n5060;
wire      [7:0] n5061;
wire            n5062;
wire      [7:0] n5063;
wire            n5064;
wire      [7:0] n5065;
wire            n5066;
wire      [7:0] n5067;
wire            n5068;
wire      [7:0] n5069;
wire            n507;
wire            n5070;
wire      [7:0] n5071;
wire            n5072;
wire      [7:0] n5073;
wire            n5074;
wire      [7:0] n5075;
wire            n5076;
wire      [7:0] n5077;
wire            n5078;
wire      [7:0] n5079;
wire            n5080;
wire      [7:0] n5081;
wire            n5082;
wire      [7:0] n5083;
wire            n5084;
wire      [7:0] n5085;
wire            n5086;
wire      [7:0] n5087;
wire            n5088;
wire      [7:0] n5089;
wire      [7:0] n509;
wire            n5090;
wire      [7:0] n5091;
wire            n5092;
wire      [7:0] n5093;
wire            n5094;
wire      [7:0] n5095;
wire            n5096;
wire      [7:0] n5097;
wire            n5098;
wire      [7:0] n5099;
wire            n510;
wire            n5100;
wire      [7:0] n5101;
wire            n5102;
wire      [7:0] n5103;
wire            n5104;
wire      [7:0] n5105;
wire            n5106;
wire      [7:0] n5107;
wire            n5108;
wire      [7:0] n5109;
wire            n5110;
wire      [7:0] n5111;
wire            n5112;
wire      [7:0] n5113;
wire            n5114;
wire      [7:0] n5115;
wire            n5116;
wire      [7:0] n5117;
wire            n5118;
wire      [7:0] n5119;
wire      [7:0] n512;
wire            n5120;
wire      [7:0] n5121;
wire            n5122;
wire      [7:0] n5123;
wire            n5124;
wire      [7:0] n5125;
wire            n5126;
wire      [7:0] n5127;
wire            n5128;
wire      [7:0] n5129;
wire            n5130;
wire      [7:0] n5131;
wire            n5132;
wire      [7:0] n5133;
wire            n5134;
wire      [7:0] n5135;
wire            n5136;
wire      [7:0] n5137;
wire            n5138;
wire      [7:0] n5139;
wire            n514;
wire            n5140;
wire      [7:0] n5141;
wire            n5142;
wire      [7:0] n5143;
wire            n5144;
wire      [7:0] n5145;
wire            n5146;
wire      [7:0] n5147;
wire            n5148;
wire      [7:0] n5149;
wire      [7:0] n515;
wire            n5150;
wire      [7:0] n5151;
wire            n5152;
wire      [7:0] n5153;
wire            n5154;
wire      [7:0] n5155;
wire            n5156;
wire      [7:0] n5157;
wire            n5158;
wire      [7:0] n5159;
wire            n5160;
wire      [7:0] n5161;
wire            n5162;
wire      [7:0] n5163;
wire            n5164;
wire      [7:0] n5165;
wire            n5166;
wire      [7:0] n5167;
wire            n5168;
wire      [7:0] n5169;
wire            n517;
wire            n5170;
wire      [7:0] n5171;
wire            n5172;
wire      [7:0] n5173;
wire            n5174;
wire      [7:0] n5175;
wire            n5176;
wire      [7:0] n5177;
wire            n5178;
wire      [7:0] n5179;
wire            n5180;
wire      [7:0] n5181;
wire            n5182;
wire      [7:0] n5183;
wire            n5184;
wire      [7:0] n5185;
wire            n5186;
wire      [7:0] n5187;
wire            n5188;
wire      [7:0] n5189;
wire      [7:0] n519;
wire            n5190;
wire      [7:0] n5191;
wire            n5192;
wire      [7:0] n5193;
wire            n5194;
wire      [7:0] n5195;
wire            n5196;
wire      [7:0] n5197;
wire            n5198;
wire      [7:0] n5199;
wire      [7:0] n52;
wire            n520;
wire            n5200;
wire      [7:0] n5201;
wire            n5202;
wire      [7:0] n5203;
wire            n5204;
wire      [7:0] n5205;
wire            n5206;
wire      [7:0] n5207;
wire            n5208;
wire      [7:0] n5209;
wire      [7:0] n521;
wire            n5210;
wire      [7:0] n5211;
wire            n5212;
wire      [7:0] n5213;
wire            n5214;
wire      [7:0] n5215;
wire            n5216;
wire      [7:0] n5217;
wire            n5218;
wire      [7:0] n5219;
wire            n522;
wire            n5220;
wire      [7:0] n5221;
wire            n5222;
wire      [7:0] n5223;
wire            n5224;
wire      [7:0] n5225;
wire            n5226;
wire      [7:0] n5227;
wire            n5228;
wire      [7:0] n5229;
wire            n5230;
wire      [7:0] n5231;
wire            n5232;
wire      [7:0] n5233;
wire            n5234;
wire      [7:0] n5235;
wire            n5236;
wire      [7:0] n5237;
wire            n5238;
wire      [7:0] n5239;
wire      [7:0] n524;
wire            n5240;
wire      [7:0] n5241;
wire            n5242;
wire      [7:0] n5243;
wire            n5244;
wire      [7:0] n5245;
wire            n5246;
wire      [7:0] n5247;
wire            n5248;
wire      [7:0] n5249;
wire            n5250;
wire      [7:0] n5251;
wire            n5252;
wire      [7:0] n5253;
wire            n5254;
wire      [7:0] n5255;
wire            n5256;
wire      [7:0] n5257;
wire            n5258;
wire      [7:0] n5259;
wire            n526;
wire            n5260;
wire      [7:0] n5261;
wire            n5262;
wire      [7:0] n5263;
wire            n5264;
wire      [7:0] n5265;
wire            n5266;
wire      [7:0] n5267;
wire            n5268;
wire      [7:0] n5269;
wire      [7:0] n527;
wire            n5270;
wire      [7:0] n5271;
wire            n5272;
wire      [7:0] n5273;
wire            n5274;
wire      [7:0] n5275;
wire            n5276;
wire      [7:0] n5277;
wire            n5278;
wire      [7:0] n5279;
wire            n528;
wire            n5280;
wire      [7:0] n5281;
wire            n5282;
wire      [7:0] n5283;
wire            n5284;
wire      [7:0] n5285;
wire            n5286;
wire      [7:0] n5287;
wire            n5288;
wire      [7:0] n5289;
wire            n5290;
wire      [7:0] n5291;
wire            n5292;
wire      [7:0] n5293;
wire            n5294;
wire      [7:0] n5295;
wire            n5296;
wire      [7:0] n5297;
wire            n5298;
wire      [7:0] n5299;
wire      [7:0] n530;
wire            n5300;
wire      [7:0] n5301;
wire            n5302;
wire      [7:0] n5303;
wire            n5304;
wire      [7:0] n5305;
wire            n5306;
wire      [7:0] n5307;
wire            n5308;
wire      [7:0] n5309;
wire            n531;
wire            n5310;
wire      [7:0] n5311;
wire            n5312;
wire      [7:0] n5313;
wire            n5314;
wire      [7:0] n5315;
wire            n5316;
wire      [7:0] n5317;
wire            n5318;
wire      [7:0] n5319;
wire            n5320;
wire      [7:0] n5321;
wire            n5322;
wire      [7:0] n5323;
wire            n5324;
wire      [7:0] n5325;
wire            n5326;
wire      [7:0] n5327;
wire            n5328;
wire      [7:0] n5329;
wire      [7:0] n533;
wire            n5330;
wire      [7:0] n5331;
wire            n5332;
wire      [7:0] n5333;
wire            n5334;
wire      [7:0] n5335;
wire            n5336;
wire      [7:0] n5337;
wire            n5338;
wire      [7:0] n5339;
wire            n534;
wire            n5340;
wire      [7:0] n5341;
wire            n5342;
wire      [7:0] n5343;
wire            n5344;
wire      [7:0] n5345;
wire            n5346;
wire      [7:0] n5347;
wire            n5348;
wire      [7:0] n5349;
wire            n5350;
wire      [7:0] n5351;
wire            n5352;
wire      [7:0] n5353;
wire            n5354;
wire      [7:0] n5355;
wire            n5356;
wire      [7:0] n5357;
wire            n5358;
wire      [7:0] n5359;
wire      [7:0] n536;
wire            n5360;
wire      [7:0] n5361;
wire            n5362;
wire      [7:0] n5363;
wire            n5364;
wire      [7:0] n5365;
wire            n5366;
wire      [7:0] n5367;
wire            n5368;
wire      [7:0] n5369;
wire            n5370;
wire      [7:0] n5371;
wire            n5372;
wire      [7:0] n5373;
wire            n5374;
wire      [7:0] n5375;
wire            n5376;
wire      [7:0] n5377;
wire            n5378;
wire      [7:0] n5379;
wire            n538;
wire            n5380;
wire      [7:0] n5381;
wire            n5382;
wire      [7:0] n5383;
wire            n5384;
wire      [7:0] n5385;
wire            n5386;
wire      [7:0] n5387;
wire            n5388;
wire      [7:0] n5389;
wire      [7:0] n539;
wire            n5390;
wire      [7:0] n5391;
wire            n5392;
wire      [7:0] n5393;
wire            n5394;
wire      [7:0] n5395;
wire            n5396;
wire      [7:0] n5397;
wire            n5398;
wire      [7:0] n5399;
wire            n54;
wire            n540;
wire            n5400;
wire      [7:0] n5401;
wire            n5402;
wire      [7:0] n5403;
wire            n5404;
wire      [7:0] n5405;
wire            n5406;
wire      [7:0] n5407;
wire            n5408;
wire      [7:0] n5409;
wire      [7:0] n541;
wire            n5410;
wire      [7:0] n5411;
wire            n5412;
wire      [7:0] n5413;
wire            n5414;
wire      [7:0] n5415;
wire            n5416;
wire      [7:0] n5417;
wire            n5418;
wire      [7:0] n5419;
wire            n542;
wire            n5420;
wire      [7:0] n5421;
wire            n5422;
wire      [7:0] n5423;
wire            n5424;
wire      [7:0] n5425;
wire            n5426;
wire      [7:0] n5427;
wire            n5428;
wire      [7:0] n5429;
wire      [7:0] n543;
wire            n5430;
wire      [7:0] n5431;
wire            n5432;
wire      [7:0] n5433;
wire            n5434;
wire      [7:0] n5435;
wire            n5436;
wire      [7:0] n5437;
wire            n5438;
wire      [7:0] n5439;
wire            n544;
wire            n5440;
wire      [7:0] n5441;
wire            n5442;
wire      [7:0] n5443;
wire            n5444;
wire      [7:0] n5445;
wire            n5446;
wire      [7:0] n5447;
wire            n5448;
wire      [7:0] n5449;
wire      [7:0] n545;
wire            n5450;
wire      [7:0] n5451;
wire            n5452;
wire      [7:0] n5453;
wire            n5454;
wire      [7:0] n5455;
wire            n5456;
wire      [7:0] n5457;
wire            n5458;
wire      [7:0] n5459;
wire            n546;
wire            n5460;
wire      [7:0] n5461;
wire            n5462;
wire      [7:0] n5463;
wire            n5464;
wire      [7:0] n5465;
wire            n5466;
wire      [7:0] n5467;
wire            n5468;
wire      [7:0] n5469;
wire      [7:0] n547;
wire            n5470;
wire      [7:0] n5471;
wire            n5472;
wire      [7:0] n5473;
wire            n5474;
wire      [7:0] n5475;
wire            n5476;
wire      [7:0] n5477;
wire            n5478;
wire      [7:0] n5479;
wire            n548;
wire            n5480;
wire      [7:0] n5481;
wire            n5482;
wire      [7:0] n5483;
wire            n5484;
wire      [7:0] n5485;
wire      [7:0] n5486;
wire      [7:0] n5487;
wire      [7:0] n5488;
wire      [7:0] n5489;
wire      [7:0] n5490;
wire      [7:0] n5491;
wire      [7:0] n5492;
wire      [7:0] n5493;
wire      [7:0] n5494;
wire      [7:0] n5495;
wire      [7:0] n5496;
wire      [7:0] n5497;
wire      [7:0] n5498;
wire      [7:0] n5499;
wire      [7:0] n550;
wire      [7:0] n5500;
wire      [7:0] n5501;
wire      [7:0] n5502;
wire      [7:0] n5503;
wire      [7:0] n5504;
wire      [7:0] n5505;
wire      [7:0] n5506;
wire      [7:0] n5507;
wire      [7:0] n5508;
wire      [7:0] n5509;
wire            n551;
wire      [7:0] n5510;
wire      [7:0] n5511;
wire      [7:0] n5512;
wire      [7:0] n5513;
wire      [7:0] n5514;
wire      [7:0] n5515;
wire      [7:0] n5516;
wire      [7:0] n5517;
wire      [7:0] n5518;
wire      [7:0] n5519;
wire      [7:0] n5520;
wire      [7:0] n5521;
wire      [7:0] n5522;
wire      [7:0] n5523;
wire      [7:0] n5524;
wire      [7:0] n5525;
wire      [7:0] n5526;
wire      [7:0] n5527;
wire      [7:0] n5528;
wire      [7:0] n5529;
wire      [7:0] n553;
wire      [7:0] n5530;
wire      [7:0] n5531;
wire      [7:0] n5532;
wire      [7:0] n5533;
wire      [7:0] n5534;
wire      [7:0] n5535;
wire      [7:0] n5536;
wire      [7:0] n5537;
wire      [7:0] n5538;
wire      [7:0] n5539;
wire            n554;
wire      [7:0] n5540;
wire      [7:0] n5541;
wire      [7:0] n5542;
wire      [7:0] n5543;
wire      [7:0] n5544;
wire      [7:0] n5545;
wire      [7:0] n5546;
wire      [7:0] n5547;
wire      [7:0] n5548;
wire      [7:0] n5549;
wire      [7:0] n5550;
wire      [7:0] n5551;
wire      [7:0] n5552;
wire      [7:0] n5553;
wire      [7:0] n5554;
wire      [7:0] n5555;
wire      [7:0] n5556;
wire      [7:0] n5557;
wire      [7:0] n5558;
wire      [7:0] n5559;
wire      [7:0] n556;
wire      [7:0] n5560;
wire      [7:0] n5561;
wire      [7:0] n5562;
wire      [7:0] n5563;
wire      [7:0] n5564;
wire      [7:0] n5565;
wire      [7:0] n5566;
wire      [7:0] n5567;
wire      [7:0] n5568;
wire      [7:0] n5569;
wire      [7:0] n5570;
wire      [7:0] n5571;
wire      [7:0] n5572;
wire      [7:0] n5573;
wire      [7:0] n5574;
wire      [7:0] n5575;
wire      [7:0] n5576;
wire      [7:0] n5577;
wire      [7:0] n5578;
wire      [7:0] n5579;
wire            n558;
wire      [7:0] n5580;
wire      [7:0] n5581;
wire      [7:0] n5582;
wire      [7:0] n5583;
wire      [7:0] n5584;
wire      [7:0] n5585;
wire      [7:0] n5586;
wire      [7:0] n5587;
wire      [7:0] n5588;
wire      [7:0] n5589;
wire      [7:0] n5590;
wire      [7:0] n5591;
wire      [7:0] n5592;
wire      [7:0] n5593;
wire      [7:0] n5594;
wire      [7:0] n5595;
wire      [7:0] n5596;
wire      [7:0] n5597;
wire      [7:0] n5598;
wire      [7:0] n5599;
wire      [7:0] n56;
wire      [7:0] n560;
wire      [7:0] n5600;
wire      [7:0] n5601;
wire      [7:0] n5602;
wire      [7:0] n5603;
wire      [7:0] n5604;
wire      [7:0] n5605;
wire      [7:0] n5606;
wire      [7:0] n5607;
wire      [7:0] n5608;
wire      [7:0] n5609;
wire      [7:0] n5610;
wire      [7:0] n5611;
wire      [7:0] n5612;
wire      [7:0] n5613;
wire      [7:0] n5614;
wire      [7:0] n5615;
wire      [7:0] n5616;
wire      [7:0] n5617;
wire      [7:0] n5618;
wire      [7:0] n5619;
wire            n562;
wire      [7:0] n5620;
wire      [7:0] n5621;
wire      [7:0] n5622;
wire      [7:0] n5623;
wire      [7:0] n5624;
wire      [7:0] n5625;
wire      [7:0] n5626;
wire      [7:0] n5627;
wire      [7:0] n5628;
wire      [7:0] n5629;
wire      [7:0] n563;
wire      [7:0] n5630;
wire      [7:0] n5631;
wire      [7:0] n5632;
wire      [7:0] n5633;
wire      [7:0] n5634;
wire      [7:0] n5635;
wire      [7:0] n5636;
wire      [7:0] n5637;
wire      [7:0] n5638;
wire      [7:0] n5639;
wire      [7:0] n5640;
wire      [7:0] n5641;
wire      [7:0] n5642;
wire      [7:0] n5643;
wire      [7:0] n5644;
wire      [7:0] n5645;
wire      [7:0] n5646;
wire      [7:0] n5647;
wire      [7:0] n5648;
wire      [7:0] n5649;
wire            n565;
wire      [7:0] n5650;
wire      [7:0] n5651;
wire      [7:0] n5652;
wire      [7:0] n5653;
wire      [7:0] n5654;
wire      [7:0] n5655;
wire      [7:0] n5656;
wire      [7:0] n5657;
wire      [7:0] n5658;
wire      [7:0] n5659;
wire      [7:0] n566;
wire      [7:0] n5660;
wire      [7:0] n5661;
wire      [7:0] n5662;
wire      [7:0] n5663;
wire      [7:0] n5664;
wire      [7:0] n5665;
wire      [7:0] n5666;
wire      [7:0] n5667;
wire      [7:0] n5668;
wire      [7:0] n5669;
wire            n567;
wire      [7:0] n5670;
wire      [7:0] n5671;
wire      [7:0] n5672;
wire      [7:0] n5673;
wire      [7:0] n5674;
wire      [7:0] n5675;
wire      [7:0] n5676;
wire      [7:0] n5677;
wire      [7:0] n5678;
wire      [7:0] n5679;
wire      [7:0] n568;
wire      [7:0] n5680;
wire      [7:0] n5681;
wire      [7:0] n5682;
wire      [7:0] n5683;
wire      [7:0] n5684;
wire      [7:0] n5685;
wire      [7:0] n5686;
wire      [7:0] n5687;
wire      [7:0] n5688;
wire      [7:0] n5689;
wire            n569;
wire      [7:0] n5690;
wire      [7:0] n5691;
wire      [7:0] n5692;
wire      [7:0] n5693;
wire      [7:0] n5694;
wire      [7:0] n5695;
wire      [7:0] n5696;
wire      [7:0] n5697;
wire      [7:0] n5698;
wire      [7:0] n5699;
wire      [7:0] n570;
wire      [7:0] n5700;
wire      [7:0] n5701;
wire      [7:0] n5702;
wire      [7:0] n5703;
wire      [7:0] n5704;
wire      [7:0] n5705;
wire      [7:0] n5706;
wire      [7:0] n5707;
wire      [7:0] n5708;
wire      [7:0] n5709;
wire            n571;
wire      [7:0] n5710;
wire      [7:0] n5711;
wire      [7:0] n5712;
wire      [7:0] n5713;
wire      [7:0] n5714;
wire      [7:0] n5715;
wire      [7:0] n5716;
wire      [7:0] n5717;
wire      [7:0] n5718;
wire      [7:0] n5719;
wire      [7:0] n572;
wire      [7:0] n5720;
wire      [7:0] n5721;
wire      [7:0] n5722;
wire      [7:0] n5723;
wire      [7:0] n5724;
wire      [7:0] n5725;
wire      [7:0] n5726;
wire      [7:0] n5727;
wire      [7:0] n5728;
wire      [7:0] n5729;
wire            n573;
wire      [7:0] n5730;
wire      [7:0] n5731;
wire      [7:0] n5732;
wire      [7:0] n5733;
wire      [7:0] n5734;
wire      [7:0] n5735;
wire      [7:0] n5736;
wire      [7:0] n5737;
wire      [7:0] n5738;
wire      [7:0] n5739;
wire      [7:0] n574;
wire      [7:0] n5740;
wire      [7:0] n5741;
wire     [23:0] n5742;
wire      [7:0] n5743;
wire      [7:0] n5744;
wire            n5745;
wire      [7:0] n5746;
wire            n5747;
wire      [7:0] n5748;
wire            n5749;
wire            n575;
wire      [7:0] n5750;
wire            n5751;
wire      [7:0] n5752;
wire            n5753;
wire      [7:0] n5754;
wire            n5755;
wire      [7:0] n5756;
wire            n5757;
wire      [7:0] n5758;
wire            n5759;
wire      [7:0] n5760;
wire            n5761;
wire      [7:0] n5762;
wire            n5763;
wire      [7:0] n5764;
wire            n5765;
wire      [7:0] n5766;
wire            n5767;
wire      [7:0] n5768;
wire            n5769;
wire      [7:0] n577;
wire      [7:0] n5770;
wire            n5771;
wire      [7:0] n5772;
wire            n5773;
wire      [7:0] n5774;
wire            n5775;
wire      [7:0] n5776;
wire            n5777;
wire      [7:0] n5778;
wire            n5779;
wire      [7:0] n5780;
wire            n5781;
wire      [7:0] n5782;
wire            n5783;
wire      [7:0] n5784;
wire            n5785;
wire      [7:0] n5786;
wire            n5787;
wire      [7:0] n5788;
wire            n5789;
wire            n579;
wire      [7:0] n5790;
wire            n5791;
wire      [7:0] n5792;
wire            n5793;
wire      [7:0] n5794;
wire            n5795;
wire      [7:0] n5796;
wire            n5797;
wire      [7:0] n5798;
wire            n5799;
wire            n58;
wire      [7:0] n580;
wire      [7:0] n5800;
wire            n5801;
wire      [7:0] n5802;
wire            n5803;
wire      [7:0] n5804;
wire            n5805;
wire      [7:0] n5806;
wire            n5807;
wire      [7:0] n5808;
wire            n5809;
wire      [7:0] n5810;
wire            n5811;
wire      [7:0] n5812;
wire            n5813;
wire      [7:0] n5814;
wire            n5815;
wire      [7:0] n5816;
wire            n5817;
wire      [7:0] n5818;
wire            n5819;
wire            n582;
wire      [7:0] n5820;
wire            n5821;
wire      [7:0] n5822;
wire            n5823;
wire      [7:0] n5824;
wire            n5825;
wire      [7:0] n5826;
wire            n5827;
wire      [7:0] n5828;
wire            n5829;
wire      [7:0] n5830;
wire            n5831;
wire      [7:0] n5832;
wire            n5833;
wire      [7:0] n5834;
wire            n5835;
wire      [7:0] n5836;
wire            n5837;
wire      [7:0] n5838;
wire            n5839;
wire      [7:0] n584;
wire      [7:0] n5840;
wire            n5841;
wire      [7:0] n5842;
wire            n5843;
wire      [7:0] n5844;
wire            n5845;
wire      [7:0] n5846;
wire            n5847;
wire      [7:0] n5848;
wire            n5849;
wire            n585;
wire      [7:0] n5850;
wire            n5851;
wire      [7:0] n5852;
wire            n5853;
wire      [7:0] n5854;
wire            n5855;
wire      [7:0] n5856;
wire            n5857;
wire      [7:0] n5858;
wire            n5859;
wire      [7:0] n586;
wire      [7:0] n5860;
wire            n5861;
wire      [7:0] n5862;
wire            n5863;
wire      [7:0] n5864;
wire            n5865;
wire      [7:0] n5866;
wire            n5867;
wire      [7:0] n5868;
wire            n5869;
wire            n587;
wire      [7:0] n5870;
wire            n5871;
wire      [7:0] n5872;
wire            n5873;
wire      [7:0] n5874;
wire            n5875;
wire      [7:0] n5876;
wire            n5877;
wire      [7:0] n5878;
wire            n5879;
wire      [7:0] n588;
wire      [7:0] n5880;
wire            n5881;
wire      [7:0] n5882;
wire            n5883;
wire      [7:0] n5884;
wire            n5885;
wire      [7:0] n5886;
wire            n5887;
wire      [7:0] n5888;
wire            n5889;
wire            n589;
wire      [7:0] n5890;
wire            n5891;
wire      [7:0] n5892;
wire            n5893;
wire      [7:0] n5894;
wire            n5895;
wire      [7:0] n5896;
wire            n5897;
wire      [7:0] n5898;
wire            n5899;
wire      [7:0] n590;
wire      [7:0] n5900;
wire            n5901;
wire      [7:0] n5902;
wire            n5903;
wire      [7:0] n5904;
wire            n5905;
wire      [7:0] n5906;
wire            n5907;
wire      [7:0] n5908;
wire            n5909;
wire            n591;
wire      [7:0] n5910;
wire            n5911;
wire      [7:0] n5912;
wire            n5913;
wire      [7:0] n5914;
wire            n5915;
wire      [7:0] n5916;
wire            n5917;
wire      [7:0] n5918;
wire            n5919;
wire      [7:0] n5920;
wire            n5921;
wire      [7:0] n5922;
wire            n5923;
wire      [7:0] n5924;
wire            n5925;
wire      [7:0] n5926;
wire            n5927;
wire      [7:0] n5928;
wire            n5929;
wire      [7:0] n593;
wire      [7:0] n5930;
wire            n5931;
wire      [7:0] n5932;
wire            n5933;
wire      [7:0] n5934;
wire            n5935;
wire      [7:0] n5936;
wire            n5937;
wire      [7:0] n5938;
wire            n5939;
wire            n594;
wire      [7:0] n5940;
wire            n5941;
wire      [7:0] n5942;
wire            n5943;
wire      [7:0] n5944;
wire            n5945;
wire      [7:0] n5946;
wire            n5947;
wire      [7:0] n5948;
wire            n5949;
wire      [7:0] n595;
wire      [7:0] n5950;
wire            n5951;
wire      [7:0] n5952;
wire            n5953;
wire      [7:0] n5954;
wire            n5955;
wire      [7:0] n5956;
wire            n5957;
wire      [7:0] n5958;
wire            n5959;
wire            n596;
wire      [7:0] n5960;
wire            n5961;
wire      [7:0] n5962;
wire            n5963;
wire      [7:0] n5964;
wire            n5965;
wire      [7:0] n5966;
wire            n5967;
wire      [7:0] n5968;
wire            n5969;
wire      [7:0] n5970;
wire            n5971;
wire      [7:0] n5972;
wire            n5973;
wire      [7:0] n5974;
wire            n5975;
wire      [7:0] n5976;
wire            n5977;
wire      [7:0] n5978;
wire            n5979;
wire      [7:0] n598;
wire      [7:0] n5980;
wire            n5981;
wire      [7:0] n5982;
wire            n5983;
wire      [7:0] n5984;
wire            n5985;
wire      [7:0] n5986;
wire            n5987;
wire      [7:0] n5988;
wire            n5989;
wire            n599;
wire      [7:0] n5990;
wire            n5991;
wire      [7:0] n5992;
wire            n5993;
wire      [7:0] n5994;
wire            n5995;
wire      [7:0] n5996;
wire            n5997;
wire      [7:0] n5998;
wire            n5999;
wire            n6;
wire      [7:0] n60;
wire      [7:0] n600;
wire      [7:0] n6000;
wire            n6001;
wire      [7:0] n6002;
wire            n6003;
wire      [7:0] n6004;
wire            n6005;
wire      [7:0] n6006;
wire            n6007;
wire      [7:0] n6008;
wire            n6009;
wire            n601;
wire      [7:0] n6010;
wire            n6011;
wire      [7:0] n6012;
wire            n6013;
wire      [7:0] n6014;
wire            n6015;
wire      [7:0] n6016;
wire            n6017;
wire      [7:0] n6018;
wire            n6019;
wire      [7:0] n602;
wire      [7:0] n6020;
wire            n6021;
wire      [7:0] n6022;
wire            n6023;
wire      [7:0] n6024;
wire            n6025;
wire      [7:0] n6026;
wire            n6027;
wire      [7:0] n6028;
wire            n6029;
wire            n603;
wire      [7:0] n6030;
wire            n6031;
wire      [7:0] n6032;
wire            n6033;
wire      [7:0] n6034;
wire            n6035;
wire      [7:0] n6036;
wire            n6037;
wire      [7:0] n6038;
wire            n6039;
wire      [7:0] n6040;
wire            n6041;
wire      [7:0] n6042;
wire            n6043;
wire      [7:0] n6044;
wire            n6045;
wire      [7:0] n6046;
wire            n6047;
wire      [7:0] n6048;
wire            n6049;
wire      [7:0] n605;
wire      [7:0] n6050;
wire            n6051;
wire      [7:0] n6052;
wire            n6053;
wire      [7:0] n6054;
wire            n6055;
wire      [7:0] n6056;
wire            n6057;
wire      [7:0] n6058;
wire            n6059;
wire            n606;
wire      [7:0] n6060;
wire            n6061;
wire      [7:0] n6062;
wire            n6063;
wire      [7:0] n6064;
wire            n6065;
wire      [7:0] n6066;
wire            n6067;
wire      [7:0] n6068;
wire            n6069;
wire      [7:0] n607;
wire      [7:0] n6070;
wire            n6071;
wire      [7:0] n6072;
wire            n6073;
wire      [7:0] n6074;
wire            n6075;
wire      [7:0] n6076;
wire            n6077;
wire      [7:0] n6078;
wire            n6079;
wire      [7:0] n6080;
wire            n6081;
wire      [7:0] n6082;
wire            n6083;
wire      [7:0] n6084;
wire            n6085;
wire      [7:0] n6086;
wire            n6087;
wire      [7:0] n6088;
wire            n6089;
wire            n609;
wire      [7:0] n6090;
wire            n6091;
wire      [7:0] n6092;
wire            n6093;
wire      [7:0] n6094;
wire            n6095;
wire      [7:0] n6096;
wire            n6097;
wire      [7:0] n6098;
wire            n6099;
wire      [7:0] n610;
wire      [7:0] n6100;
wire            n6101;
wire      [7:0] n6102;
wire            n6103;
wire      [7:0] n6104;
wire            n6105;
wire      [7:0] n6106;
wire            n6107;
wire      [7:0] n6108;
wire            n6109;
wire            n611;
wire      [7:0] n6110;
wire            n6111;
wire      [7:0] n6112;
wire            n6113;
wire      [7:0] n6114;
wire            n6115;
wire      [7:0] n6116;
wire            n6117;
wire      [7:0] n6118;
wire            n6119;
wire      [7:0] n612;
wire      [7:0] n6120;
wire            n6121;
wire      [7:0] n6122;
wire            n6123;
wire      [7:0] n6124;
wire            n6125;
wire      [7:0] n6126;
wire            n6127;
wire      [7:0] n6128;
wire            n6129;
wire            n613;
wire      [7:0] n6130;
wire            n6131;
wire      [7:0] n6132;
wire            n6133;
wire      [7:0] n6134;
wire            n6135;
wire      [7:0] n6136;
wire            n6137;
wire      [7:0] n6138;
wire            n6139;
wire      [7:0] n614;
wire      [7:0] n6140;
wire            n6141;
wire      [7:0] n6142;
wire            n6143;
wire      [7:0] n6144;
wire            n6145;
wire      [7:0] n6146;
wire            n6147;
wire      [7:0] n6148;
wire            n6149;
wire            n615;
wire      [7:0] n6150;
wire            n6151;
wire      [7:0] n6152;
wire            n6153;
wire      [7:0] n6154;
wire            n6155;
wire      [7:0] n6156;
wire            n6157;
wire      [7:0] n6158;
wire            n6159;
wire      [7:0] n6160;
wire            n6161;
wire      [7:0] n6162;
wire            n6163;
wire      [7:0] n6164;
wire            n6165;
wire      [7:0] n6166;
wire            n6167;
wire      [7:0] n6168;
wire            n6169;
wire      [7:0] n617;
wire      [7:0] n6170;
wire            n6171;
wire      [7:0] n6172;
wire            n6173;
wire      [7:0] n6174;
wire            n6175;
wire      [7:0] n6176;
wire            n6177;
wire      [7:0] n6178;
wire            n6179;
wire            n618;
wire      [7:0] n6180;
wire            n6181;
wire      [7:0] n6182;
wire            n6183;
wire      [7:0] n6184;
wire            n6185;
wire      [7:0] n6186;
wire            n6187;
wire      [7:0] n6188;
wire            n6189;
wire      [7:0] n6190;
wire            n6191;
wire      [7:0] n6192;
wire            n6193;
wire      [7:0] n6194;
wire            n6195;
wire      [7:0] n6196;
wire            n6197;
wire      [7:0] n6198;
wire            n6199;
wire            n62;
wire      [7:0] n620;
wire      [7:0] n6200;
wire            n6201;
wire      [7:0] n6202;
wire            n6203;
wire      [7:0] n6204;
wire            n6205;
wire      [7:0] n6206;
wire            n6207;
wire      [7:0] n6208;
wire            n6209;
wire            n621;
wire      [7:0] n6210;
wire            n6211;
wire      [7:0] n6212;
wire            n6213;
wire      [7:0] n6214;
wire            n6215;
wire      [7:0] n6216;
wire            n6217;
wire      [7:0] n6218;
wire            n6219;
wire      [7:0] n6220;
wire            n6221;
wire      [7:0] n6222;
wire            n6223;
wire      [7:0] n6224;
wire            n6225;
wire      [7:0] n6226;
wire            n6227;
wire      [7:0] n6228;
wire            n6229;
wire      [7:0] n623;
wire      [7:0] n6230;
wire            n6231;
wire      [7:0] n6232;
wire            n6233;
wire      [7:0] n6234;
wire            n6235;
wire      [7:0] n6236;
wire            n6237;
wire      [7:0] n6238;
wire            n6239;
wire            n624;
wire      [7:0] n6240;
wire            n6241;
wire      [7:0] n6242;
wire            n6243;
wire      [7:0] n6244;
wire            n6245;
wire      [7:0] n6246;
wire            n6247;
wire      [7:0] n6248;
wire            n6249;
wire      [7:0] n625;
wire      [7:0] n6250;
wire            n6251;
wire      [7:0] n6252;
wire            n6253;
wire      [7:0] n6254;
wire            n6255;
wire      [7:0] n6256;
wire      [7:0] n6257;
wire      [7:0] n6258;
wire      [7:0] n6259;
wire            n626;
wire      [7:0] n6260;
wire      [7:0] n6261;
wire      [7:0] n6262;
wire      [7:0] n6263;
wire      [7:0] n6264;
wire      [7:0] n6265;
wire      [7:0] n6266;
wire      [7:0] n6267;
wire      [7:0] n6268;
wire      [7:0] n6269;
wire      [7:0] n6270;
wire      [7:0] n6271;
wire      [7:0] n6272;
wire      [7:0] n6273;
wire      [7:0] n6274;
wire      [7:0] n6275;
wire      [7:0] n6276;
wire      [7:0] n6277;
wire      [7:0] n6278;
wire      [7:0] n6279;
wire      [7:0] n628;
wire      [7:0] n6280;
wire      [7:0] n6281;
wire      [7:0] n6282;
wire      [7:0] n6283;
wire      [7:0] n6284;
wire      [7:0] n6285;
wire      [7:0] n6286;
wire      [7:0] n6287;
wire      [7:0] n6288;
wire      [7:0] n6289;
wire      [7:0] n6290;
wire      [7:0] n6291;
wire      [7:0] n6292;
wire      [7:0] n6293;
wire      [7:0] n6294;
wire      [7:0] n6295;
wire      [7:0] n6296;
wire      [7:0] n6297;
wire      [7:0] n6298;
wire      [7:0] n6299;
wire            n630;
wire      [7:0] n6300;
wire      [7:0] n6301;
wire      [7:0] n6302;
wire      [7:0] n6303;
wire      [7:0] n6304;
wire      [7:0] n6305;
wire      [7:0] n6306;
wire      [7:0] n6307;
wire      [7:0] n6308;
wire      [7:0] n6309;
wire      [7:0] n631;
wire      [7:0] n6310;
wire      [7:0] n6311;
wire      [7:0] n6312;
wire      [7:0] n6313;
wire      [7:0] n6314;
wire      [7:0] n6315;
wire      [7:0] n6316;
wire      [7:0] n6317;
wire      [7:0] n6318;
wire      [7:0] n6319;
wire            n632;
wire      [7:0] n6320;
wire      [7:0] n6321;
wire      [7:0] n6322;
wire      [7:0] n6323;
wire      [7:0] n6324;
wire      [7:0] n6325;
wire      [7:0] n6326;
wire      [7:0] n6327;
wire      [7:0] n6328;
wire      [7:0] n6329;
wire      [7:0] n633;
wire      [7:0] n6330;
wire      [7:0] n6331;
wire      [7:0] n6332;
wire      [7:0] n6333;
wire      [7:0] n6334;
wire      [7:0] n6335;
wire      [7:0] n6336;
wire      [7:0] n6337;
wire      [7:0] n6338;
wire      [7:0] n6339;
wire            n634;
wire      [7:0] n6340;
wire      [7:0] n6341;
wire      [7:0] n6342;
wire      [7:0] n6343;
wire      [7:0] n6344;
wire      [7:0] n6345;
wire      [7:0] n6346;
wire      [7:0] n6347;
wire      [7:0] n6348;
wire      [7:0] n6349;
wire      [7:0] n6350;
wire      [7:0] n6351;
wire      [7:0] n6352;
wire      [7:0] n6353;
wire      [7:0] n6354;
wire      [7:0] n6355;
wire      [7:0] n6356;
wire      [7:0] n6357;
wire      [7:0] n6358;
wire      [7:0] n6359;
wire      [7:0] n636;
wire      [7:0] n6360;
wire      [7:0] n6361;
wire      [7:0] n6362;
wire      [7:0] n6363;
wire      [7:0] n6364;
wire      [7:0] n6365;
wire      [7:0] n6366;
wire      [7:0] n6367;
wire      [7:0] n6368;
wire      [7:0] n6369;
wire            n637;
wire      [7:0] n6370;
wire      [7:0] n6371;
wire      [7:0] n6372;
wire      [7:0] n6373;
wire      [7:0] n6374;
wire      [7:0] n6375;
wire      [7:0] n6376;
wire      [7:0] n6377;
wire      [7:0] n6378;
wire      [7:0] n6379;
wire      [7:0] n638;
wire      [7:0] n6380;
wire      [7:0] n6381;
wire      [7:0] n6382;
wire      [7:0] n6383;
wire      [7:0] n6384;
wire      [7:0] n6385;
wire      [7:0] n6386;
wire      [7:0] n6387;
wire      [7:0] n6388;
wire      [7:0] n6389;
wire            n639;
wire      [7:0] n6390;
wire      [7:0] n6391;
wire      [7:0] n6392;
wire      [7:0] n6393;
wire      [7:0] n6394;
wire      [7:0] n6395;
wire      [7:0] n6396;
wire      [7:0] n6397;
wire      [7:0] n6398;
wire      [7:0] n6399;
wire      [7:0] n64;
wire      [7:0] n640;
wire      [7:0] n6400;
wire      [7:0] n6401;
wire      [7:0] n6402;
wire      [7:0] n6403;
wire      [7:0] n6404;
wire      [7:0] n6405;
wire      [7:0] n6406;
wire      [7:0] n6407;
wire      [7:0] n6408;
wire      [7:0] n6409;
wire            n641;
wire      [7:0] n6410;
wire      [7:0] n6411;
wire      [7:0] n6412;
wire      [7:0] n6413;
wire      [7:0] n6414;
wire      [7:0] n6415;
wire      [7:0] n6416;
wire      [7:0] n6417;
wire      [7:0] n6418;
wire      [7:0] n6419;
wire      [7:0] n642;
wire      [7:0] n6420;
wire      [7:0] n6421;
wire      [7:0] n6422;
wire      [7:0] n6423;
wire      [7:0] n6424;
wire      [7:0] n6425;
wire      [7:0] n6426;
wire      [7:0] n6427;
wire      [7:0] n6428;
wire      [7:0] n6429;
wire            n643;
wire      [7:0] n6430;
wire      [7:0] n6431;
wire      [7:0] n6432;
wire      [7:0] n6433;
wire      [7:0] n6434;
wire      [7:0] n6435;
wire      [7:0] n6436;
wire      [7:0] n6437;
wire      [7:0] n6438;
wire      [7:0] n6439;
wire      [7:0] n6440;
wire      [7:0] n6441;
wire      [7:0] n6442;
wire      [7:0] n6443;
wire      [7:0] n6444;
wire      [7:0] n6445;
wire      [7:0] n6446;
wire      [7:0] n6447;
wire      [7:0] n6448;
wire      [7:0] n6449;
wire      [7:0] n645;
wire      [7:0] n6450;
wire      [7:0] n6451;
wire      [7:0] n6452;
wire      [7:0] n6453;
wire      [7:0] n6454;
wire      [7:0] n6455;
wire      [7:0] n6456;
wire      [7:0] n6457;
wire      [7:0] n6458;
wire      [7:0] n6459;
wire            n646;
wire      [7:0] n6460;
wire      [7:0] n6461;
wire      [7:0] n6462;
wire      [7:0] n6463;
wire      [7:0] n6464;
wire      [7:0] n6465;
wire      [7:0] n6466;
wire      [7:0] n6467;
wire      [7:0] n6468;
wire      [7:0] n6469;
wire      [7:0] n6470;
wire      [7:0] n6471;
wire      [7:0] n6472;
wire      [7:0] n6473;
wire      [7:0] n6474;
wire      [7:0] n6475;
wire      [7:0] n6476;
wire      [7:0] n6477;
wire      [7:0] n6478;
wire      [7:0] n6479;
wire      [7:0] n648;
wire      [7:0] n6480;
wire      [7:0] n6481;
wire      [7:0] n6482;
wire      [7:0] n6483;
wire      [7:0] n6484;
wire      [7:0] n6485;
wire      [7:0] n6486;
wire      [7:0] n6487;
wire      [7:0] n6488;
wire      [7:0] n6489;
wire            n649;
wire      [7:0] n6490;
wire      [7:0] n6491;
wire      [7:0] n6492;
wire      [7:0] n6493;
wire      [7:0] n6494;
wire      [7:0] n6495;
wire      [7:0] n6496;
wire      [7:0] n6497;
wire      [7:0] n6498;
wire      [7:0] n6499;
wire      [7:0] n650;
wire      [7:0] n6500;
wire      [7:0] n6501;
wire      [7:0] n6502;
wire      [7:0] n6503;
wire      [7:0] n6504;
wire      [7:0] n6505;
wire      [7:0] n6506;
wire      [7:0] n6507;
wire      [7:0] n6508;
wire      [7:0] n6509;
wire      [7:0] n6510;
wire      [7:0] n6511;
wire      [7:0] n6512;
wire     [31:0] n6513;
wire      [7:0] n6514;
wire      [7:0] n6515;
wire      [7:0] n6516;
wire      [7:0] n6517;
wire      [7:0] n6518;
wire     [39:0] n6519;
wire            n652;
wire      [7:0] n6520;
wire      [7:0] n6521;
wire      [7:0] n6522;
wire      [7:0] n6523;
wire     [47:0] n6524;
wire      [7:0] n6525;
wire      [7:0] n6526;
wire      [7:0] n6527;
wire      [7:0] n6528;
wire     [55:0] n6529;
wire      [7:0] n6530;
wire      [7:0] n6531;
wire      [7:0] n6532;
wire      [7:0] n6533;
wire     [63:0] n6534;
wire      [7:0] n6535;
wire      [7:0] n6536;
wire      [7:0] n6537;
wire      [7:0] n6538;
wire      [7:0] n6539;
wire      [7:0] n654;
wire      [7:0] n6540;
wire      [7:0] n6541;
wire     [71:0] n6542;
wire      [7:0] n6543;
wire      [7:0] n6544;
wire      [7:0] n6545;
wire      [7:0] n6546;
wire      [7:0] n6547;
wire      [7:0] n6548;
wire     [79:0] n6549;
wire            n655;
wire      [7:0] n6550;
wire      [7:0] n6551;
wire      [7:0] n6552;
wire      [7:0] n6553;
wire      [7:0] n6554;
wire      [7:0] n6555;
wire     [87:0] n6556;
wire      [7:0] n6557;
wire      [7:0] n6558;
wire      [7:0] n6559;
wire      [7:0] n656;
wire      [7:0] n6560;
wire      [7:0] n6561;
wire      [7:0] n6562;
wire     [95:0] n6563;
wire      [7:0] n6564;
wire      [7:0] n6565;
wire      [7:0] n6566;
wire      [7:0] n6567;
wire      [7:0] n6568;
wire      [7:0] n6569;
wire      [7:0] n6570;
wire      [7:0] n6571;
wire      [7:0] n6572;
wire    [103:0] n6573;
wire      [7:0] n6574;
wire      [7:0] n6575;
wire      [7:0] n6576;
wire      [7:0] n6577;
wire      [7:0] n6578;
wire      [7:0] n6579;
wire            n658;
wire      [7:0] n6580;
wire      [7:0] n6581;
wire    [111:0] n6582;
wire      [7:0] n6583;
wire      [7:0] n6584;
wire      [7:0] n6585;
wire      [7:0] n6586;
wire      [7:0] n6587;
wire      [7:0] n6588;
wire      [7:0] n6589;
wire      [7:0] n6590;
wire    [119:0] n6591;
wire      [7:0] n6592;
wire      [7:0] n6593;
wire      [7:0] n6594;
wire      [7:0] n6595;
wire      [7:0] n6596;
wire      [7:0] n6597;
wire      [7:0] n6598;
wire      [7:0] n6599;
wire            n66;
wire      [7:0] n660;
wire    [127:0] n6600;
wire    [127:0] n6601;
wire            n661;
wire      [7:0] n662;
wire            n663;
wire      [7:0] n665;
wire            n667;
wire      [7:0] n668;
wire            n670;
wire      [7:0] n672;
wire            n673;
wire      [7:0] n675;
wire            n676;
wire      [7:0] n677;
wire            n678;
wire      [7:0] n679;
wire      [7:0] n68;
wire            n680;
wire      [7:0] n681;
wire            n683;
wire      [7:0] n684;
wire            n685;
wire      [7:0] n686;
wire            n687;
wire      [7:0] n688;
wire            n689;
wire      [7:0] n690;
wire            n691;
wire      [7:0] n692;
wire            n694;
wire      [7:0] n695;
wire            n696;
wire      [7:0] n697;
wire            n698;
wire      [7:0] n699;
wire            n70;
wire            n700;
wire      [7:0] n701;
wire            n702;
wire      [7:0] n703;
wire            n704;
wire      [7:0] n705;
wire            n706;
wire      [7:0] n707;
wire            n708;
wire      [7:0] n709;
wire            n710;
wire      [7:0] n711;
wire            n712;
wire      [7:0] n713;
wire            n714;
wire      [7:0] n715;
wire            n716;
wire      [7:0] n717;
wire            n718;
wire      [7:0] n719;
wire      [7:0] n72;
wire            n720;
wire      [7:0] n721;
wire            n722;
wire      [7:0] n723;
wire            n724;
wire      [7:0] n725;
wire            n726;
wire      [7:0] n727;
wire            n728;
wire      [7:0] n729;
wire            n730;
wire      [7:0] n731;
wire            n732;
wire      [7:0] n733;
wire            n734;
wire      [7:0] n735;
wire            n736;
wire      [7:0] n737;
wire            n738;
wire      [7:0] n739;
wire            n74;
wire            n740;
wire      [7:0] n741;
wire            n742;
wire      [7:0] n743;
wire            n744;
wire      [7:0] n745;
wire            n746;
wire      [7:0] n747;
wire            n748;
wire      [7:0] n749;
wire            n750;
wire      [7:0] n751;
wire            n752;
wire      [7:0] n754;
wire            n755;
wire      [7:0] n756;
wire            n757;
wire      [7:0] n758;
wire            n759;
wire      [7:0] n76;
wire      [7:0] n760;
wire            n761;
wire      [7:0] n762;
wire            n763;
wire      [7:0] n764;
wire            n765;
wire      [7:0] n766;
wire            n767;
wire      [7:0] n768;
wire            n769;
wire      [7:0] n770;
wire            n771;
wire      [7:0] n772;
wire      [7:0] n773;
wire      [7:0] n774;
wire      [7:0] n775;
wire      [7:0] n776;
wire      [7:0] n777;
wire      [7:0] n778;
wire      [7:0] n779;
wire            n78;
wire      [7:0] n780;
wire      [7:0] n781;
wire      [7:0] n782;
wire      [7:0] n783;
wire      [7:0] n784;
wire      [7:0] n785;
wire      [7:0] n786;
wire      [7:0] n787;
wire      [7:0] n788;
wire      [7:0] n789;
wire      [7:0] n790;
wire      [7:0] n791;
wire      [7:0] n792;
wire      [7:0] n793;
wire      [7:0] n794;
wire      [7:0] n795;
wire      [7:0] n796;
wire      [7:0] n797;
wire      [7:0] n798;
wire      [7:0] n799;
wire      [7:0] n8;
wire      [7:0] n80;
wire      [7:0] n800;
wire      [7:0] n801;
wire      [7:0] n802;
wire      [7:0] n803;
wire      [7:0] n804;
wire      [7:0] n805;
wire      [7:0] n806;
wire      [7:0] n807;
wire      [7:0] n808;
wire      [7:0] n809;
wire      [7:0] n810;
wire      [7:0] n811;
wire      [7:0] n812;
wire      [7:0] n813;
wire      [7:0] n814;
wire      [7:0] n815;
wire      [7:0] n816;
wire      [7:0] n817;
wire      [7:0] n818;
wire      [7:0] n819;
wire            n82;
wire      [7:0] n820;
wire      [7:0] n821;
wire      [7:0] n822;
wire      [7:0] n823;
wire      [7:0] n824;
wire      [7:0] n825;
wire      [7:0] n826;
wire      [7:0] n827;
wire      [7:0] n828;
wire      [7:0] n829;
wire      [7:0] n830;
wire      [7:0] n831;
wire      [7:0] n832;
wire      [7:0] n833;
wire      [7:0] n834;
wire      [7:0] n835;
wire      [7:0] n836;
wire      [7:0] n837;
wire      [7:0] n838;
wire      [7:0] n839;
wire      [7:0] n84;
wire      [7:0] n840;
wire      [7:0] n841;
wire      [7:0] n842;
wire      [7:0] n843;
wire      [7:0] n844;
wire      [7:0] n845;
wire      [7:0] n846;
wire      [7:0] n847;
wire      [7:0] n848;
wire      [7:0] n849;
wire      [7:0] n850;
wire      [7:0] n851;
wire      [7:0] n852;
wire      [7:0] n853;
wire      [7:0] n854;
wire      [7:0] n855;
wire      [7:0] n856;
wire      [7:0] n857;
wire      [7:0] n858;
wire      [7:0] n859;
wire            n86;
wire      [7:0] n860;
wire      [7:0] n861;
wire      [7:0] n862;
wire      [7:0] n863;
wire      [7:0] n864;
wire      [7:0] n865;
wire      [7:0] n866;
wire      [7:0] n867;
wire      [7:0] n868;
wire      [7:0] n869;
wire      [7:0] n870;
wire      [7:0] n871;
wire      [7:0] n872;
wire      [7:0] n873;
wire      [7:0] n874;
wire      [7:0] n875;
wire      [7:0] n876;
wire      [7:0] n877;
wire      [7:0] n878;
wire      [7:0] n879;
wire      [7:0] n88;
wire      [7:0] n880;
wire      [7:0] n881;
wire      [7:0] n882;
wire      [7:0] n883;
wire      [7:0] n884;
wire      [7:0] n885;
wire      [7:0] n886;
wire      [7:0] n887;
wire      [7:0] n888;
wire      [7:0] n889;
wire      [7:0] n890;
wire      [7:0] n891;
wire      [7:0] n892;
wire      [7:0] n893;
wire      [7:0] n894;
wire      [7:0] n895;
wire      [7:0] n896;
wire      [7:0] n897;
wire      [7:0] n898;
wire      [7:0] n899;
wire            n90;
wire      [7:0] n900;
wire      [7:0] n901;
wire      [7:0] n902;
wire      [7:0] n903;
wire      [7:0] n904;
wire      [7:0] n905;
wire      [7:0] n906;
wire      [7:0] n907;
wire      [7:0] n908;
wire      [7:0] n909;
wire      [7:0] n910;
wire      [7:0] n911;
wire      [7:0] n912;
wire      [7:0] n913;
wire      [7:0] n914;
wire      [7:0] n915;
wire      [7:0] n916;
wire      [7:0] n917;
wire      [7:0] n918;
wire      [7:0] n919;
wire      [7:0] n92;
wire      [7:0] n920;
wire      [7:0] n921;
wire      [7:0] n922;
wire      [7:0] n923;
wire      [7:0] n924;
wire      [7:0] n925;
wire      [7:0] n926;
wire      [7:0] n927;
wire      [7:0] n928;
wire      [7:0] n929;
wire            n93;
wire      [7:0] n930;
wire      [7:0] n931;
wire      [7:0] n932;
wire      [7:0] n933;
wire      [7:0] n934;
wire      [7:0] n935;
wire      [7:0] n936;
wire      [7:0] n937;
wire      [7:0] n938;
wire      [7:0] n939;
wire      [7:0] n940;
wire      [7:0] n941;
wire      [7:0] n942;
wire      [7:0] n943;
wire      [7:0] n944;
wire      [7:0] n945;
wire      [7:0] n946;
wire      [7:0] n947;
wire      [7:0] n948;
wire      [7:0] n949;
wire      [7:0] n95;
wire      [7:0] n950;
wire      [7:0] n951;
wire      [7:0] n952;
wire      [7:0] n953;
wire      [7:0] n954;
wire      [7:0] n955;
wire      [7:0] n956;
wire      [7:0] n957;
wire      [7:0] n958;
wire      [7:0] n959;
wire      [7:0] n960;
wire      [7:0] n961;
wire      [7:0] n962;
wire      [7:0] n963;
wire      [7:0] n964;
wire      [7:0] n965;
wire      [7:0] n966;
wire      [7:0] n967;
wire      [7:0] n968;
wire      [7:0] n969;
wire            n97;
wire      [7:0] n970;
wire      [7:0] n971;
wire      [7:0] n972;
wire      [7:0] n973;
wire      [7:0] n974;
wire      [7:0] n975;
wire      [7:0] n976;
wire      [7:0] n977;
wire      [7:0] n978;
wire      [7:0] n979;
wire      [7:0] n980;
wire      [7:0] n981;
wire      [7:0] n982;
wire      [7:0] n983;
wire      [7:0] n984;
wire      [7:0] n985;
wire      [7:0] n986;
wire      [7:0] n987;
wire      [7:0] n988;
wire      [7:0] n989;
wire      [7:0] n99;
wire      [7:0] n990;
wire      [7:0] n991;
wire      [7:0] n992;
wire      [7:0] n993;
wire      [7:0] n994;
wire      [7:0] n995;
wire      [7:0] n996;
wire      [7:0] n997;
wire      [7:0] n998;
wire      [7:0] n999;
(* keep *) wire    [127:0] out_1_randinit;
(* keep *) wire    [127:0] out_2_randinit;
(* keep *) wire      [7:0] rcon_randinit;
wire            rst;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign bv_128_0_n1 = 128'h0 ;
assign n2 = in[127:120] ;
assign n3 =  ( n2 ) ^ ( rcon )  ;
assign n4 = in[23:16] ;
assign bv_8_255_n5 = 8'hff ;
assign n6 =  ( n4 ) == ( bv_8_255_n5 )  ;
assign bv_8_22_n7 = 8'h16 ;
assign n8 = in[23:16] ;
assign bv_8_254_n9 = 8'hfe ;
assign n10 =  ( n8 ) == ( bv_8_254_n9 )  ;
assign bv_8_187_n11 = 8'hbb ;
assign n12 = in[23:16] ;
assign bv_8_253_n13 = 8'hfd ;
assign n14 =  ( n12 ) == ( bv_8_253_n13 )  ;
assign bv_8_84_n15 = 8'h54 ;
assign n16 = in[23:16] ;
assign bv_8_252_n17 = 8'hfc ;
assign n18 =  ( n16 ) == ( bv_8_252_n17 )  ;
assign bv_8_176_n19 = 8'hb0 ;
assign n20 = in[23:16] ;
assign bv_8_251_n21 = 8'hfb ;
assign n22 =  ( n20 ) == ( bv_8_251_n21 )  ;
assign bv_8_15_n23 = 8'hf ;
assign n24 = in[23:16] ;
assign bv_8_250_n25 = 8'hfa ;
assign n26 =  ( n24 ) == ( bv_8_250_n25 )  ;
assign bv_8_45_n27 = 8'h2d ;
assign n28 = in[23:16] ;
assign bv_8_249_n29 = 8'hf9 ;
assign n30 =  ( n28 ) == ( bv_8_249_n29 )  ;
assign bv_8_153_n31 = 8'h99 ;
assign n32 = in[23:16] ;
assign bv_8_248_n33 = 8'hf8 ;
assign n34 =  ( n32 ) == ( bv_8_248_n33 )  ;
assign bv_8_65_n35 = 8'h41 ;
assign n36 = in[23:16] ;
assign bv_8_247_n37 = 8'hf7 ;
assign n38 =  ( n36 ) == ( bv_8_247_n37 )  ;
assign bv_8_104_n39 = 8'h68 ;
assign n40 = in[23:16] ;
assign bv_8_246_n41 = 8'hf6 ;
assign n42 =  ( n40 ) == ( bv_8_246_n41 )  ;
assign bv_8_66_n43 = 8'h42 ;
assign n44 = in[23:16] ;
assign bv_8_245_n45 = 8'hf5 ;
assign n46 =  ( n44 ) == ( bv_8_245_n45 )  ;
assign bv_8_230_n47 = 8'he6 ;
assign n48 = in[23:16] ;
assign bv_8_244_n49 = 8'hf4 ;
assign n50 =  ( n48 ) == ( bv_8_244_n49 )  ;
assign bv_8_191_n51 = 8'hbf ;
assign n52 = in[23:16] ;
assign bv_8_243_n53 = 8'hf3 ;
assign n54 =  ( n52 ) == ( bv_8_243_n53 )  ;
assign bv_8_13_n55 = 8'hd ;
assign n56 = in[23:16] ;
assign bv_8_242_n57 = 8'hf2 ;
assign n58 =  ( n56 ) == ( bv_8_242_n57 )  ;
assign bv_8_137_n59 = 8'h89 ;
assign n60 = in[23:16] ;
assign bv_8_241_n61 = 8'hf1 ;
assign n62 =  ( n60 ) == ( bv_8_241_n61 )  ;
assign bv_8_161_n63 = 8'ha1 ;
assign n64 = in[23:16] ;
assign bv_8_240_n65 = 8'hf0 ;
assign n66 =  ( n64 ) == ( bv_8_240_n65 )  ;
assign bv_8_140_n67 = 8'h8c ;
assign n68 = in[23:16] ;
assign bv_8_239_n69 = 8'hef ;
assign n70 =  ( n68 ) == ( bv_8_239_n69 )  ;
assign bv_8_223_n71 = 8'hdf ;
assign n72 = in[23:16] ;
assign bv_8_238_n73 = 8'hee ;
assign n74 =  ( n72 ) == ( bv_8_238_n73 )  ;
assign bv_8_40_n75 = 8'h28 ;
assign n76 = in[23:16] ;
assign bv_8_237_n77 = 8'hed ;
assign n78 =  ( n76 ) == ( bv_8_237_n77 )  ;
assign bv_8_85_n79 = 8'h55 ;
assign n80 = in[23:16] ;
assign bv_8_236_n81 = 8'hec ;
assign n82 =  ( n80 ) == ( bv_8_236_n81 )  ;
assign bv_8_206_n83 = 8'hce ;
assign n84 = in[23:16] ;
assign bv_8_235_n85 = 8'heb ;
assign n86 =  ( n84 ) == ( bv_8_235_n85 )  ;
assign bv_8_233_n87 = 8'he9 ;
assign n88 = in[23:16] ;
assign bv_8_234_n89 = 8'hea ;
assign n90 =  ( n88 ) == ( bv_8_234_n89 )  ;
assign bv_8_135_n91 = 8'h87 ;
assign n92 = in[23:16] ;
assign n93 =  ( n92 ) == ( bv_8_233_n87 )  ;
assign bv_8_30_n94 = 8'h1e ;
assign n95 = in[23:16] ;
assign bv_8_232_n96 = 8'he8 ;
assign n97 =  ( n95 ) == ( bv_8_232_n96 )  ;
assign bv_8_155_n98 = 8'h9b ;
assign n99 = in[23:16] ;
assign bv_8_231_n100 = 8'he7 ;
assign n101 =  ( n99 ) == ( bv_8_231_n100 )  ;
assign bv_8_148_n102 = 8'h94 ;
assign n103 = in[23:16] ;
assign n104 =  ( n103 ) == ( bv_8_230_n47 )  ;
assign bv_8_142_n105 = 8'h8e ;
assign n106 = in[23:16] ;
assign bv_8_229_n107 = 8'he5 ;
assign n108 =  ( n106 ) == ( bv_8_229_n107 )  ;
assign bv_8_217_n109 = 8'hd9 ;
assign n110 = in[23:16] ;
assign bv_8_228_n111 = 8'he4 ;
assign n112 =  ( n110 ) == ( bv_8_228_n111 )  ;
assign bv_8_105_n113 = 8'h69 ;
assign n114 = in[23:16] ;
assign bv_8_227_n115 = 8'he3 ;
assign n116 =  ( n114 ) == ( bv_8_227_n115 )  ;
assign bv_8_17_n117 = 8'h11 ;
assign n118 = in[23:16] ;
assign bv_8_226_n119 = 8'he2 ;
assign n120 =  ( n118 ) == ( bv_8_226_n119 )  ;
assign bv_8_152_n121 = 8'h98 ;
assign n122 = in[23:16] ;
assign bv_8_225_n123 = 8'he1 ;
assign n124 =  ( n122 ) == ( bv_8_225_n123 )  ;
assign n125 = in[23:16] ;
assign bv_8_224_n126 = 8'he0 ;
assign n127 =  ( n125 ) == ( bv_8_224_n126 )  ;
assign n128 = in[23:16] ;
assign n129 =  ( n128 ) == ( bv_8_223_n71 )  ;
assign bv_8_158_n130 = 8'h9e ;
assign n131 = in[23:16] ;
assign bv_8_222_n132 = 8'hde ;
assign n133 =  ( n131 ) == ( bv_8_222_n132 )  ;
assign bv_8_29_n134 = 8'h1d ;
assign n135 = in[23:16] ;
assign bv_8_221_n136 = 8'hdd ;
assign n137 =  ( n135 ) == ( bv_8_221_n136 )  ;
assign bv_8_193_n138 = 8'hc1 ;
assign n139 = in[23:16] ;
assign bv_8_220_n140 = 8'hdc ;
assign n141 =  ( n139 ) == ( bv_8_220_n140 )  ;
assign bv_8_134_n142 = 8'h86 ;
assign n143 = in[23:16] ;
assign bv_8_219_n144 = 8'hdb ;
assign n145 =  ( n143 ) == ( bv_8_219_n144 )  ;
assign bv_8_185_n146 = 8'hb9 ;
assign n147 = in[23:16] ;
assign bv_8_218_n148 = 8'hda ;
assign n149 =  ( n147 ) == ( bv_8_218_n148 )  ;
assign bv_8_87_n150 = 8'h57 ;
assign n151 = in[23:16] ;
assign n152 =  ( n151 ) == ( bv_8_217_n109 )  ;
assign bv_8_53_n153 = 8'h35 ;
assign n154 = in[23:16] ;
assign bv_8_216_n155 = 8'hd8 ;
assign n156 =  ( n154 ) == ( bv_8_216_n155 )  ;
assign bv_8_97_n157 = 8'h61 ;
assign n158 = in[23:16] ;
assign bv_8_215_n159 = 8'hd7 ;
assign n160 =  ( n158 ) == ( bv_8_215_n159 )  ;
assign bv_8_14_n161 = 8'he ;
assign n162 = in[23:16] ;
assign bv_8_214_n163 = 8'hd6 ;
assign n164 =  ( n162 ) == ( bv_8_214_n163 )  ;
assign n165 = in[23:16] ;
assign bv_8_213_n166 = 8'hd5 ;
assign n167 =  ( n165 ) == ( bv_8_213_n166 )  ;
assign bv_8_3_n168 = 8'h3 ;
assign n169 = in[23:16] ;
assign bv_8_212_n170 = 8'hd4 ;
assign n171 =  ( n169 ) == ( bv_8_212_n170 )  ;
assign bv_8_72_n172 = 8'h48 ;
assign n173 = in[23:16] ;
assign bv_8_211_n174 = 8'hd3 ;
assign n175 =  ( n173 ) == ( bv_8_211_n174 )  ;
assign bv_8_102_n176 = 8'h66 ;
assign n177 = in[23:16] ;
assign bv_8_210_n178 = 8'hd2 ;
assign n179 =  ( n177 ) == ( bv_8_210_n178 )  ;
assign bv_8_181_n180 = 8'hb5 ;
assign n181 = in[23:16] ;
assign bv_8_209_n182 = 8'hd1 ;
assign n183 =  ( n181 ) == ( bv_8_209_n182 )  ;
assign bv_8_62_n184 = 8'h3e ;
assign n185 = in[23:16] ;
assign bv_8_208_n186 = 8'hd0 ;
assign n187 =  ( n185 ) == ( bv_8_208_n186 )  ;
assign bv_8_112_n188 = 8'h70 ;
assign n189 = in[23:16] ;
assign bv_8_207_n190 = 8'hcf ;
assign n191 =  ( n189 ) == ( bv_8_207_n190 )  ;
assign bv_8_138_n192 = 8'h8a ;
assign n193 = in[23:16] ;
assign n194 =  ( n193 ) == ( bv_8_206_n83 )  ;
assign bv_8_139_n195 = 8'h8b ;
assign n196 = in[23:16] ;
assign bv_8_205_n197 = 8'hcd ;
assign n198 =  ( n196 ) == ( bv_8_205_n197 )  ;
assign bv_8_189_n199 = 8'hbd ;
assign n200 = in[23:16] ;
assign bv_8_204_n201 = 8'hcc ;
assign n202 =  ( n200 ) == ( bv_8_204_n201 )  ;
assign bv_8_75_n203 = 8'h4b ;
assign n204 = in[23:16] ;
assign bv_8_203_n205 = 8'hcb ;
assign n206 =  ( n204 ) == ( bv_8_203_n205 )  ;
assign bv_8_31_n207 = 8'h1f ;
assign n208 = in[23:16] ;
assign bv_8_202_n209 = 8'hca ;
assign n210 =  ( n208 ) == ( bv_8_202_n209 )  ;
assign bv_8_116_n211 = 8'h74 ;
assign n212 = in[23:16] ;
assign bv_8_201_n213 = 8'hc9 ;
assign n214 =  ( n212 ) == ( bv_8_201_n213 )  ;
assign n215 = in[23:16] ;
assign bv_8_200_n216 = 8'hc8 ;
assign n217 =  ( n215 ) == ( bv_8_200_n216 )  ;
assign n218 = in[23:16] ;
assign bv_8_199_n219 = 8'hc7 ;
assign n220 =  ( n218 ) == ( bv_8_199_n219 )  ;
assign bv_8_198_n221 = 8'hc6 ;
assign n222 = in[23:16] ;
assign n223 =  ( n222 ) == ( bv_8_198_n221 )  ;
assign bv_8_180_n224 = 8'hb4 ;
assign n225 = in[23:16] ;
assign bv_8_197_n226 = 8'hc5 ;
assign n227 =  ( n225 ) == ( bv_8_197_n226 )  ;
assign bv_8_166_n228 = 8'ha6 ;
assign n229 = in[23:16] ;
assign bv_8_196_n230 = 8'hc4 ;
assign n231 =  ( n229 ) == ( bv_8_196_n230 )  ;
assign bv_8_28_n232 = 8'h1c ;
assign n233 = in[23:16] ;
assign bv_8_195_n234 = 8'hc3 ;
assign n235 =  ( n233 ) == ( bv_8_195_n234 )  ;
assign bv_8_46_n236 = 8'h2e ;
assign n237 = in[23:16] ;
assign bv_8_194_n238 = 8'hc2 ;
assign n239 =  ( n237 ) == ( bv_8_194_n238 )  ;
assign bv_8_37_n240 = 8'h25 ;
assign n241 = in[23:16] ;
assign n242 =  ( n241 ) == ( bv_8_193_n138 )  ;
assign bv_8_120_n243 = 8'h78 ;
assign n244 = in[23:16] ;
assign bv_8_192_n245 = 8'hc0 ;
assign n246 =  ( n244 ) == ( bv_8_192_n245 )  ;
assign bv_8_186_n247 = 8'hba ;
assign n248 = in[23:16] ;
assign n249 =  ( n248 ) == ( bv_8_191_n51 )  ;
assign bv_8_8_n250 = 8'h8 ;
assign n251 = in[23:16] ;
assign bv_8_190_n252 = 8'hbe ;
assign n253 =  ( n251 ) == ( bv_8_190_n252 )  ;
assign bv_8_174_n254 = 8'hae ;
assign n255 = in[23:16] ;
assign n256 =  ( n255 ) == ( bv_8_189_n199 )  ;
assign bv_8_122_n257 = 8'h7a ;
assign n258 = in[23:16] ;
assign bv_8_188_n259 = 8'hbc ;
assign n260 =  ( n258 ) == ( bv_8_188_n259 )  ;
assign bv_8_101_n261 = 8'h65 ;
assign n262 = in[23:16] ;
assign n263 =  ( n262 ) == ( bv_8_187_n11 )  ;
assign n264 = in[23:16] ;
assign n265 =  ( n264 ) == ( bv_8_186_n247 )  ;
assign n266 = in[23:16] ;
assign n267 =  ( n266 ) == ( bv_8_185_n146 )  ;
assign bv_8_86_n268 = 8'h56 ;
assign n269 = in[23:16] ;
assign bv_8_184_n270 = 8'hb8 ;
assign n271 =  ( n269 ) == ( bv_8_184_n270 )  ;
assign bv_8_108_n272 = 8'h6c ;
assign n273 = in[23:16] ;
assign bv_8_183_n274 = 8'hb7 ;
assign n275 =  ( n273 ) == ( bv_8_183_n274 )  ;
assign bv_8_169_n276 = 8'ha9 ;
assign n277 = in[23:16] ;
assign bv_8_182_n278 = 8'hb6 ;
assign n279 =  ( n277 ) == ( bv_8_182_n278 )  ;
assign bv_8_78_n280 = 8'h4e ;
assign n281 = in[23:16] ;
assign n282 =  ( n281 ) == ( bv_8_181_n180 )  ;
assign n283 = in[23:16] ;
assign n284 =  ( n283 ) == ( bv_8_180_n224 )  ;
assign bv_8_141_n285 = 8'h8d ;
assign n286 = in[23:16] ;
assign bv_8_179_n287 = 8'hb3 ;
assign n288 =  ( n286 ) == ( bv_8_179_n287 )  ;
assign bv_8_109_n289 = 8'h6d ;
assign n290 = in[23:16] ;
assign bv_8_178_n291 = 8'hb2 ;
assign n292 =  ( n290 ) == ( bv_8_178_n291 )  ;
assign bv_8_55_n293 = 8'h37 ;
assign n294 = in[23:16] ;
assign bv_8_177_n295 = 8'hb1 ;
assign n296 =  ( n294 ) == ( bv_8_177_n295 )  ;
assign n297 = in[23:16] ;
assign n298 =  ( n297 ) == ( bv_8_176_n19 )  ;
assign n299 = in[23:16] ;
assign bv_8_175_n300 = 8'haf ;
assign n301 =  ( n299 ) == ( bv_8_175_n300 )  ;
assign bv_8_121_n302 = 8'h79 ;
assign n303 = in[23:16] ;
assign n304 =  ( n303 ) == ( bv_8_174_n254 )  ;
assign n305 = in[23:16] ;
assign bv_8_173_n306 = 8'had ;
assign n307 =  ( n305 ) == ( bv_8_173_n306 )  ;
assign bv_8_149_n308 = 8'h95 ;
assign n309 = in[23:16] ;
assign bv_8_172_n310 = 8'hac ;
assign n311 =  ( n309 ) == ( bv_8_172_n310 )  ;
assign bv_8_145_n312 = 8'h91 ;
assign n313 = in[23:16] ;
assign bv_8_171_n314 = 8'hab ;
assign n315 =  ( n313 ) == ( bv_8_171_n314 )  ;
assign bv_8_98_n316 = 8'h62 ;
assign n317 = in[23:16] ;
assign bv_8_170_n318 = 8'haa ;
assign n319 =  ( n317 ) == ( bv_8_170_n318 )  ;
assign n320 = in[23:16] ;
assign n321 =  ( n320 ) == ( bv_8_169_n276 )  ;
assign n322 = in[23:16] ;
assign bv_8_168_n323 = 8'ha8 ;
assign n324 =  ( n322 ) == ( bv_8_168_n323 )  ;
assign n325 = in[23:16] ;
assign bv_8_167_n326 = 8'ha7 ;
assign n327 =  ( n325 ) == ( bv_8_167_n326 )  ;
assign bv_8_92_n328 = 8'h5c ;
assign n329 = in[23:16] ;
assign n330 =  ( n329 ) == ( bv_8_166_n228 )  ;
assign bv_8_36_n331 = 8'h24 ;
assign n332 = in[23:16] ;
assign bv_8_165_n333 = 8'ha5 ;
assign n334 =  ( n332 ) == ( bv_8_165_n333 )  ;
assign bv_8_6_n335 = 8'h6 ;
assign n336 = in[23:16] ;
assign bv_8_164_n337 = 8'ha4 ;
assign n338 =  ( n336 ) == ( bv_8_164_n337 )  ;
assign bv_8_73_n339 = 8'h49 ;
assign n340 = in[23:16] ;
assign bv_8_163_n341 = 8'ha3 ;
assign n342 =  ( n340 ) == ( bv_8_163_n341 )  ;
assign bv_8_10_n343 = 8'ha ;
assign n344 = in[23:16] ;
assign bv_8_162_n345 = 8'ha2 ;
assign n346 =  ( n344 ) == ( bv_8_162_n345 )  ;
assign bv_8_58_n347 = 8'h3a ;
assign n348 = in[23:16] ;
assign n349 =  ( n348 ) == ( bv_8_161_n63 )  ;
assign bv_8_50_n350 = 8'h32 ;
assign n351 = in[23:16] ;
assign bv_8_160_n352 = 8'ha0 ;
assign n353 =  ( n351 ) == ( bv_8_160_n352 )  ;
assign n354 = in[23:16] ;
assign bv_8_159_n355 = 8'h9f ;
assign n356 =  ( n354 ) == ( bv_8_159_n355 )  ;
assign n357 = in[23:16] ;
assign n358 =  ( n357 ) == ( bv_8_158_n130 )  ;
assign bv_8_11_n359 = 8'hb ;
assign n360 = in[23:16] ;
assign bv_8_157_n361 = 8'h9d ;
assign n362 =  ( n360 ) == ( bv_8_157_n361 )  ;
assign bv_8_94_n363 = 8'h5e ;
assign n364 = in[23:16] ;
assign bv_8_156_n365 = 8'h9c ;
assign n366 =  ( n364 ) == ( bv_8_156_n365 )  ;
assign n367 = in[23:16] ;
assign n368 =  ( n367 ) == ( bv_8_155_n98 )  ;
assign bv_8_20_n369 = 8'h14 ;
assign n370 = in[23:16] ;
assign bv_8_154_n371 = 8'h9a ;
assign n372 =  ( n370 ) == ( bv_8_154_n371 )  ;
assign n373 = in[23:16] ;
assign n374 =  ( n373 ) == ( bv_8_153_n31 )  ;
assign n375 = in[23:16] ;
assign n376 =  ( n375 ) == ( bv_8_152_n121 )  ;
assign bv_8_70_n377 = 8'h46 ;
assign n378 = in[23:16] ;
assign bv_8_151_n379 = 8'h97 ;
assign n380 =  ( n378 ) == ( bv_8_151_n379 )  ;
assign bv_8_136_n381 = 8'h88 ;
assign n382 = in[23:16] ;
assign bv_8_150_n383 = 8'h96 ;
assign n384 =  ( n382 ) == ( bv_8_150_n383 )  ;
assign bv_8_144_n385 = 8'h90 ;
assign n386 = in[23:16] ;
assign n387 =  ( n386 ) == ( bv_8_149_n308 )  ;
assign bv_8_42_n388 = 8'h2a ;
assign n389 = in[23:16] ;
assign n390 =  ( n389 ) == ( bv_8_148_n102 )  ;
assign bv_8_34_n391 = 8'h22 ;
assign n392 = in[23:16] ;
assign bv_8_147_n393 = 8'h93 ;
assign n394 =  ( n392 ) == ( bv_8_147_n393 )  ;
assign n395 = in[23:16] ;
assign bv_8_146_n396 = 8'h92 ;
assign n397 =  ( n395 ) == ( bv_8_146_n396 )  ;
assign bv_8_79_n398 = 8'h4f ;
assign n399 = in[23:16] ;
assign n400 =  ( n399 ) == ( bv_8_145_n312 )  ;
assign bv_8_129_n401 = 8'h81 ;
assign n402 = in[23:16] ;
assign n403 =  ( n402 ) == ( bv_8_144_n385 )  ;
assign bv_8_96_n404 = 8'h60 ;
assign n405 = in[23:16] ;
assign bv_8_143_n406 = 8'h8f ;
assign n407 =  ( n405 ) == ( bv_8_143_n406 )  ;
assign bv_8_115_n408 = 8'h73 ;
assign n409 = in[23:16] ;
assign n410 =  ( n409 ) == ( bv_8_142_n105 )  ;
assign bv_8_25_n411 = 8'h19 ;
assign n412 = in[23:16] ;
assign n413 =  ( n412 ) == ( bv_8_141_n285 )  ;
assign bv_8_93_n414 = 8'h5d ;
assign n415 = in[23:16] ;
assign n416 =  ( n415 ) == ( bv_8_140_n67 )  ;
assign bv_8_100_n417 = 8'h64 ;
assign n418 = in[23:16] ;
assign n419 =  ( n418 ) == ( bv_8_139_n195 )  ;
assign bv_8_61_n420 = 8'h3d ;
assign n421 = in[23:16] ;
assign n422 =  ( n421 ) == ( bv_8_138_n192 )  ;
assign bv_8_126_n423 = 8'h7e ;
assign n424 = in[23:16] ;
assign n425 =  ( n424 ) == ( bv_8_137_n59 )  ;
assign n426 = in[23:16] ;
assign n427 =  ( n426 ) == ( bv_8_136_n381 )  ;
assign n428 = in[23:16] ;
assign n429 =  ( n428 ) == ( bv_8_135_n91 )  ;
assign bv_8_23_n430 = 8'h17 ;
assign n431 = in[23:16] ;
assign n432 =  ( n431 ) == ( bv_8_134_n142 )  ;
assign bv_8_68_n433 = 8'h44 ;
assign n434 = in[23:16] ;
assign bv_8_133_n435 = 8'h85 ;
assign n436 =  ( n434 ) == ( bv_8_133_n435 )  ;
assign n437 = in[23:16] ;
assign bv_8_132_n438 = 8'h84 ;
assign n439 =  ( n437 ) == ( bv_8_132_n438 )  ;
assign bv_8_95_n440 = 8'h5f ;
assign n441 = in[23:16] ;
assign bv_8_131_n442 = 8'h83 ;
assign n443 =  ( n441 ) == ( bv_8_131_n442 )  ;
assign n444 = in[23:16] ;
assign bv_8_130_n445 = 8'h82 ;
assign n446 =  ( n444 ) == ( bv_8_130_n445 )  ;
assign bv_8_19_n447 = 8'h13 ;
assign n448 = in[23:16] ;
assign n449 =  ( n448 ) == ( bv_8_129_n401 )  ;
assign bv_8_12_n450 = 8'hc ;
assign n451 = in[23:16] ;
assign bv_8_128_n452 = 8'h80 ;
assign n453 =  ( n451 ) == ( bv_8_128_n452 )  ;
assign n454 = in[23:16] ;
assign bv_8_127_n455 = 8'h7f ;
assign n456 =  ( n454 ) == ( bv_8_127_n455 )  ;
assign n457 = in[23:16] ;
assign n458 =  ( n457 ) == ( bv_8_126_n423 )  ;
assign n459 = in[23:16] ;
assign bv_8_125_n460 = 8'h7d ;
assign n461 =  ( n459 ) == ( bv_8_125_n460 )  ;
assign n462 = in[23:16] ;
assign bv_8_124_n463 = 8'h7c ;
assign n464 =  ( n462 ) == ( bv_8_124_n463 )  ;
assign bv_8_16_n465 = 8'h10 ;
assign n466 = in[23:16] ;
assign bv_8_123_n467 = 8'h7b ;
assign n468 =  ( n466 ) == ( bv_8_123_n467 )  ;
assign bv_8_33_n469 = 8'h21 ;
assign n470 = in[23:16] ;
assign n471 =  ( n470 ) == ( bv_8_122_n257 )  ;
assign n472 = in[23:16] ;
assign n473 =  ( n472 ) == ( bv_8_121_n302 )  ;
assign n474 = in[23:16] ;
assign n475 =  ( n474 ) == ( bv_8_120_n243 )  ;
assign n476 = in[23:16] ;
assign bv_8_119_n477 = 8'h77 ;
assign n478 =  ( n476 ) == ( bv_8_119_n477 )  ;
assign n479 = in[23:16] ;
assign bv_8_118_n480 = 8'h76 ;
assign n481 =  ( n479 ) == ( bv_8_118_n480 )  ;
assign bv_8_56_n482 = 8'h38 ;
assign n483 = in[23:16] ;
assign bv_8_117_n484 = 8'h75 ;
assign n485 =  ( n483 ) == ( bv_8_117_n484 )  ;
assign n486 = in[23:16] ;
assign n487 =  ( n486 ) == ( bv_8_116_n211 )  ;
assign n488 = in[23:16] ;
assign n489 =  ( n488 ) == ( bv_8_115_n408 )  ;
assign n490 = in[23:16] ;
assign bv_8_114_n491 = 8'h72 ;
assign n492 =  ( n490 ) == ( bv_8_114_n491 )  ;
assign bv_8_64_n493 = 8'h40 ;
assign n494 = in[23:16] ;
assign bv_8_113_n495 = 8'h71 ;
assign n496 =  ( n494 ) == ( bv_8_113_n495 )  ;
assign n497 = in[23:16] ;
assign n498 =  ( n497 ) == ( bv_8_112_n188 )  ;
assign bv_8_81_n499 = 8'h51 ;
assign n500 = in[23:16] ;
assign bv_8_111_n501 = 8'h6f ;
assign n502 =  ( n500 ) == ( bv_8_111_n501 )  ;
assign n503 = in[23:16] ;
assign bv_8_110_n504 = 8'h6e ;
assign n505 =  ( n503 ) == ( bv_8_110_n504 )  ;
assign n506 = in[23:16] ;
assign n507 =  ( n506 ) == ( bv_8_109_n289 )  ;
assign bv_8_60_n508 = 8'h3c ;
assign n509 = in[23:16] ;
assign n510 =  ( n509 ) == ( bv_8_108_n272 )  ;
assign bv_8_80_n511 = 8'h50 ;
assign n512 = in[23:16] ;
assign bv_8_107_n513 = 8'h6b ;
assign n514 =  ( n512 ) == ( bv_8_107_n513 )  ;
assign n515 = in[23:16] ;
assign bv_8_106_n516 = 8'h6a ;
assign n517 =  ( n515 ) == ( bv_8_106_n516 )  ;
assign bv_8_2_n518 = 8'h2 ;
assign n519 = in[23:16] ;
assign n520 =  ( n519 ) == ( bv_8_105_n113 )  ;
assign n521 = in[23:16] ;
assign n522 =  ( n521 ) == ( bv_8_104_n39 )  ;
assign bv_8_69_n523 = 8'h45 ;
assign n524 = in[23:16] ;
assign bv_8_103_n525 = 8'h67 ;
assign n526 =  ( n524 ) == ( bv_8_103_n525 )  ;
assign n527 = in[23:16] ;
assign n528 =  ( n527 ) == ( bv_8_102_n176 )  ;
assign bv_8_51_n529 = 8'h33 ;
assign n530 = in[23:16] ;
assign n531 =  ( n530 ) == ( bv_8_101_n261 )  ;
assign bv_8_77_n532 = 8'h4d ;
assign n533 = in[23:16] ;
assign n534 =  ( n533 ) == ( bv_8_100_n417 )  ;
assign bv_8_67_n535 = 8'h43 ;
assign n536 = in[23:16] ;
assign bv_8_99_n537 = 8'h63 ;
assign n538 =  ( n536 ) == ( bv_8_99_n537 )  ;
assign n539 = in[23:16] ;
assign n540 =  ( n539 ) == ( bv_8_98_n316 )  ;
assign n541 = in[23:16] ;
assign n542 =  ( n541 ) == ( bv_8_97_n157 )  ;
assign n543 = in[23:16] ;
assign n544 =  ( n543 ) == ( bv_8_96_n404 )  ;
assign n545 = in[23:16] ;
assign n546 =  ( n545 ) == ( bv_8_95_n440 )  ;
assign n547 = in[23:16] ;
assign n548 =  ( n547 ) == ( bv_8_94_n363 )  ;
assign bv_8_88_n549 = 8'h58 ;
assign n550 = in[23:16] ;
assign n551 =  ( n550 ) == ( bv_8_93_n414 )  ;
assign bv_8_76_n552 = 8'h4c ;
assign n553 = in[23:16] ;
assign n554 =  ( n553 ) == ( bv_8_92_n328 )  ;
assign bv_8_74_n555 = 8'h4a ;
assign n556 = in[23:16] ;
assign bv_8_91_n557 = 8'h5b ;
assign n558 =  ( n556 ) == ( bv_8_91_n557 )  ;
assign bv_8_57_n559 = 8'h39 ;
assign n560 = in[23:16] ;
assign bv_8_90_n561 = 8'h5a ;
assign n562 =  ( n560 ) == ( bv_8_90_n561 )  ;
assign n563 = in[23:16] ;
assign bv_8_89_n564 = 8'h59 ;
assign n565 =  ( n563 ) == ( bv_8_89_n564 )  ;
assign n566 = in[23:16] ;
assign n567 =  ( n566 ) == ( bv_8_88_n549 )  ;
assign n568 = in[23:16] ;
assign n569 =  ( n568 ) == ( bv_8_87_n150 )  ;
assign n570 = in[23:16] ;
assign n571 =  ( n570 ) == ( bv_8_86_n268 )  ;
assign n572 = in[23:16] ;
assign n573 =  ( n572 ) == ( bv_8_85_n79 )  ;
assign n574 = in[23:16] ;
assign n575 =  ( n574 ) == ( bv_8_84_n15 )  ;
assign bv_8_32_n576 = 8'h20 ;
assign n577 = in[23:16] ;
assign bv_8_83_n578 = 8'h53 ;
assign n579 =  ( n577 ) == ( bv_8_83_n578 )  ;
assign n580 = in[23:16] ;
assign bv_8_82_n581 = 8'h52 ;
assign n582 =  ( n580 ) == ( bv_8_82_n581 )  ;
assign bv_8_0_n583 = 8'h0 ;
assign n584 = in[23:16] ;
assign n585 =  ( n584 ) == ( bv_8_81_n499 )  ;
assign n586 = in[23:16] ;
assign n587 =  ( n586 ) == ( bv_8_80_n511 )  ;
assign n588 = in[23:16] ;
assign n589 =  ( n588 ) == ( bv_8_79_n398 )  ;
assign n590 = in[23:16] ;
assign n591 =  ( n590 ) == ( bv_8_78_n280 )  ;
assign bv_8_47_n592 = 8'h2f ;
assign n593 = in[23:16] ;
assign n594 =  ( n593 ) == ( bv_8_77_n532 )  ;
assign n595 = in[23:16] ;
assign n596 =  ( n595 ) == ( bv_8_76_n552 )  ;
assign bv_8_41_n597 = 8'h29 ;
assign n598 = in[23:16] ;
assign n599 =  ( n598 ) == ( bv_8_75_n203 )  ;
assign n600 = in[23:16] ;
assign n601 =  ( n600 ) == ( bv_8_74_n555 )  ;
assign n602 = in[23:16] ;
assign n603 =  ( n602 ) == ( bv_8_73_n339 )  ;
assign bv_8_59_n604 = 8'h3b ;
assign n605 = in[23:16] ;
assign n606 =  ( n605 ) == ( bv_8_72_n172 )  ;
assign n607 = in[23:16] ;
assign bv_8_71_n608 = 8'h47 ;
assign n609 =  ( n607 ) == ( bv_8_71_n608 )  ;
assign n610 = in[23:16] ;
assign n611 =  ( n610 ) == ( bv_8_70_n377 )  ;
assign n612 = in[23:16] ;
assign n613 =  ( n612 ) == ( bv_8_69_n523 )  ;
assign n614 = in[23:16] ;
assign n615 =  ( n614 ) == ( bv_8_68_n433 )  ;
assign bv_8_27_n616 = 8'h1b ;
assign n617 = in[23:16] ;
assign n618 =  ( n617 ) == ( bv_8_67_n535 )  ;
assign bv_8_26_n619 = 8'h1a ;
assign n620 = in[23:16] ;
assign n621 =  ( n620 ) == ( bv_8_66_n43 )  ;
assign bv_8_44_n622 = 8'h2c ;
assign n623 = in[23:16] ;
assign n624 =  ( n623 ) == ( bv_8_65_n35 )  ;
assign n625 = in[23:16] ;
assign n626 =  ( n625 ) == ( bv_8_64_n493 )  ;
assign bv_8_9_n627 = 8'h9 ;
assign n628 = in[23:16] ;
assign bv_8_63_n629 = 8'h3f ;
assign n630 =  ( n628 ) == ( bv_8_63_n629 )  ;
assign n631 = in[23:16] ;
assign n632 =  ( n631 ) == ( bv_8_62_n184 )  ;
assign n633 = in[23:16] ;
assign n634 =  ( n633 ) == ( bv_8_61_n420 )  ;
assign bv_8_39_n635 = 8'h27 ;
assign n636 = in[23:16] ;
assign n637 =  ( n636 ) == ( bv_8_60_n508 )  ;
assign n638 = in[23:16] ;
assign n639 =  ( n638 ) == ( bv_8_59_n604 )  ;
assign n640 = in[23:16] ;
assign n641 =  ( n640 ) == ( bv_8_58_n347 )  ;
assign n642 = in[23:16] ;
assign n643 =  ( n642 ) == ( bv_8_57_n559 )  ;
assign bv_8_18_n644 = 8'h12 ;
assign n645 = in[23:16] ;
assign n646 =  ( n645 ) == ( bv_8_56_n482 )  ;
assign bv_8_7_n647 = 8'h7 ;
assign n648 = in[23:16] ;
assign n649 =  ( n648 ) == ( bv_8_55_n293 )  ;
assign n650 = in[23:16] ;
assign bv_8_54_n651 = 8'h36 ;
assign n652 =  ( n650 ) == ( bv_8_54_n651 )  ;
assign bv_8_5_n653 = 8'h5 ;
assign n654 = in[23:16] ;
assign n655 =  ( n654 ) == ( bv_8_53_n153 )  ;
assign n656 = in[23:16] ;
assign bv_8_52_n657 = 8'h34 ;
assign n658 =  ( n656 ) == ( bv_8_52_n657 )  ;
assign bv_8_24_n659 = 8'h18 ;
assign n660 = in[23:16] ;
assign n661 =  ( n660 ) == ( bv_8_51_n529 )  ;
assign n662 = in[23:16] ;
assign n663 =  ( n662 ) == ( bv_8_50_n350 )  ;
assign bv_8_35_n664 = 8'h23 ;
assign n665 = in[23:16] ;
assign bv_8_49_n666 = 8'h31 ;
assign n667 =  ( n665 ) == ( bv_8_49_n666 )  ;
assign n668 = in[23:16] ;
assign bv_8_48_n669 = 8'h30 ;
assign n670 =  ( n668 ) == ( bv_8_48_n669 )  ;
assign bv_8_4_n671 = 8'h4 ;
assign n672 = in[23:16] ;
assign n673 =  ( n672 ) == ( bv_8_47_n592 )  ;
assign bv_8_21_n674 = 8'h15 ;
assign n675 = in[23:16] ;
assign n676 =  ( n675 ) == ( bv_8_46_n236 )  ;
assign n677 = in[23:16] ;
assign n678 =  ( n677 ) == ( bv_8_45_n27 )  ;
assign n679 = in[23:16] ;
assign n680 =  ( n679 ) == ( bv_8_44_n622 )  ;
assign n681 = in[23:16] ;
assign bv_8_43_n682 = 8'h2b ;
assign n683 =  ( n681 ) == ( bv_8_43_n682 )  ;
assign n684 = in[23:16] ;
assign n685 =  ( n684 ) == ( bv_8_42_n388 )  ;
assign n686 = in[23:16] ;
assign n687 =  ( n686 ) == ( bv_8_41_n597 )  ;
assign n688 = in[23:16] ;
assign n689 =  ( n688 ) == ( bv_8_40_n75 )  ;
assign n690 = in[23:16] ;
assign n691 =  ( n690 ) == ( bv_8_39_n635 )  ;
assign n692 = in[23:16] ;
assign bv_8_38_n693 = 8'h26 ;
assign n694 =  ( n692 ) == ( bv_8_38_n693 )  ;
assign n695 = in[23:16] ;
assign n696 =  ( n695 ) == ( bv_8_37_n240 )  ;
assign n697 = in[23:16] ;
assign n698 =  ( n697 ) == ( bv_8_36_n331 )  ;
assign n699 = in[23:16] ;
assign n700 =  ( n699 ) == ( bv_8_35_n664 )  ;
assign n701 = in[23:16] ;
assign n702 =  ( n701 ) == ( bv_8_34_n391 )  ;
assign n703 = in[23:16] ;
assign n704 =  ( n703 ) == ( bv_8_33_n469 )  ;
assign n705 = in[23:16] ;
assign n706 =  ( n705 ) == ( bv_8_32_n576 )  ;
assign n707 = in[23:16] ;
assign n708 =  ( n707 ) == ( bv_8_31_n207 )  ;
assign n709 = in[23:16] ;
assign n710 =  ( n709 ) == ( bv_8_30_n94 )  ;
assign n711 = in[23:16] ;
assign n712 =  ( n711 ) == ( bv_8_29_n134 )  ;
assign n713 = in[23:16] ;
assign n714 =  ( n713 ) == ( bv_8_28_n232 )  ;
assign n715 = in[23:16] ;
assign n716 =  ( n715 ) == ( bv_8_27_n616 )  ;
assign n717 = in[23:16] ;
assign n718 =  ( n717 ) == ( bv_8_26_n619 )  ;
assign n719 = in[23:16] ;
assign n720 =  ( n719 ) == ( bv_8_25_n411 )  ;
assign n721 = in[23:16] ;
assign n722 =  ( n721 ) == ( bv_8_24_n659 )  ;
assign n723 = in[23:16] ;
assign n724 =  ( n723 ) == ( bv_8_23_n430 )  ;
assign n725 = in[23:16] ;
assign n726 =  ( n725 ) == ( bv_8_22_n7 )  ;
assign n727 = in[23:16] ;
assign n728 =  ( n727 ) == ( bv_8_21_n674 )  ;
assign n729 = in[23:16] ;
assign n730 =  ( n729 ) == ( bv_8_20_n369 )  ;
assign n731 = in[23:16] ;
assign n732 =  ( n731 ) == ( bv_8_19_n447 )  ;
assign n733 = in[23:16] ;
assign n734 =  ( n733 ) == ( bv_8_18_n644 )  ;
assign n735 = in[23:16] ;
assign n736 =  ( n735 ) == ( bv_8_17_n117 )  ;
assign n737 = in[23:16] ;
assign n738 =  ( n737 ) == ( bv_8_16_n465 )  ;
assign n739 = in[23:16] ;
assign n740 =  ( n739 ) == ( bv_8_15_n23 )  ;
assign n741 = in[23:16] ;
assign n742 =  ( n741 ) == ( bv_8_14_n161 )  ;
assign n743 = in[23:16] ;
assign n744 =  ( n743 ) == ( bv_8_13_n55 )  ;
assign n745 = in[23:16] ;
assign n746 =  ( n745 ) == ( bv_8_12_n450 )  ;
assign n747 = in[23:16] ;
assign n748 =  ( n747 ) == ( bv_8_11_n359 )  ;
assign n749 = in[23:16] ;
assign n750 =  ( n749 ) == ( bv_8_10_n343 )  ;
assign n751 = in[23:16] ;
assign n752 =  ( n751 ) == ( bv_8_9_n627 )  ;
assign bv_8_1_n753 = 8'h1 ;
assign n754 = in[23:16] ;
assign n755 =  ( n754 ) == ( bv_8_8_n250 )  ;
assign n756 = in[23:16] ;
assign n757 =  ( n756 ) == ( bv_8_7_n647 )  ;
assign n758 = in[23:16] ;
assign n759 =  ( n758 ) == ( bv_8_6_n335 )  ;
assign n760 = in[23:16] ;
assign n761 =  ( n760 ) == ( bv_8_5_n653 )  ;
assign n762 = in[23:16] ;
assign n763 =  ( n762 ) == ( bv_8_4_n671 )  ;
assign n764 = in[23:16] ;
assign n765 =  ( n764 ) == ( bv_8_3_n168 )  ;
assign n766 = in[23:16] ;
assign n767 =  ( n766 ) == ( bv_8_2_n518 )  ;
assign n768 = in[23:16] ;
assign n769 =  ( n768 ) == ( bv_8_1_n753 )  ;
assign n770 = in[23:16] ;
assign n771 =  ( n770 ) == ( bv_8_0_n583 )  ;
assign n772 =  ( n771 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n773 =  ( n769 ) ? ( bv_8_124_n463 ) : ( n772 ) ;
assign n774 =  ( n767 ) ? ( bv_8_119_n477 ) : ( n773 ) ;
assign n775 =  ( n765 ) ? ( bv_8_123_n467 ) : ( n774 ) ;
assign n776 =  ( n763 ) ? ( bv_8_242_n57 ) : ( n775 ) ;
assign n777 =  ( n761 ) ? ( bv_8_107_n513 ) : ( n776 ) ;
assign n778 =  ( n759 ) ? ( bv_8_111_n501 ) : ( n777 ) ;
assign n779 =  ( n757 ) ? ( bv_8_197_n226 ) : ( n778 ) ;
assign n780 =  ( n755 ) ? ( bv_8_48_n669 ) : ( n779 ) ;
assign n781 =  ( n752 ) ? ( bv_8_1_n753 ) : ( n780 ) ;
assign n782 =  ( n750 ) ? ( bv_8_103_n525 ) : ( n781 ) ;
assign n783 =  ( n748 ) ? ( bv_8_43_n682 ) : ( n782 ) ;
assign n784 =  ( n746 ) ? ( bv_8_254_n9 ) : ( n783 ) ;
assign n785 =  ( n744 ) ? ( bv_8_215_n159 ) : ( n784 ) ;
assign n786 =  ( n742 ) ? ( bv_8_171_n314 ) : ( n785 ) ;
assign n787 =  ( n740 ) ? ( bv_8_118_n480 ) : ( n786 ) ;
assign n788 =  ( n738 ) ? ( bv_8_202_n209 ) : ( n787 ) ;
assign n789 =  ( n736 ) ? ( bv_8_130_n445 ) : ( n788 ) ;
assign n790 =  ( n734 ) ? ( bv_8_201_n213 ) : ( n789 ) ;
assign n791 =  ( n732 ) ? ( bv_8_125_n460 ) : ( n790 ) ;
assign n792 =  ( n730 ) ? ( bv_8_250_n25 ) : ( n791 ) ;
assign n793 =  ( n728 ) ? ( bv_8_89_n564 ) : ( n792 ) ;
assign n794 =  ( n726 ) ? ( bv_8_71_n608 ) : ( n793 ) ;
assign n795 =  ( n724 ) ? ( bv_8_240_n65 ) : ( n794 ) ;
assign n796 =  ( n722 ) ? ( bv_8_173_n306 ) : ( n795 ) ;
assign n797 =  ( n720 ) ? ( bv_8_212_n170 ) : ( n796 ) ;
assign n798 =  ( n718 ) ? ( bv_8_162_n345 ) : ( n797 ) ;
assign n799 =  ( n716 ) ? ( bv_8_175_n300 ) : ( n798 ) ;
assign n800 =  ( n714 ) ? ( bv_8_156_n365 ) : ( n799 ) ;
assign n801 =  ( n712 ) ? ( bv_8_164_n337 ) : ( n800 ) ;
assign n802 =  ( n710 ) ? ( bv_8_114_n491 ) : ( n801 ) ;
assign n803 =  ( n708 ) ? ( bv_8_192_n245 ) : ( n802 ) ;
assign n804 =  ( n706 ) ? ( bv_8_183_n274 ) : ( n803 ) ;
assign n805 =  ( n704 ) ? ( bv_8_253_n13 ) : ( n804 ) ;
assign n806 =  ( n702 ) ? ( bv_8_147_n393 ) : ( n805 ) ;
assign n807 =  ( n700 ) ? ( bv_8_38_n693 ) : ( n806 ) ;
assign n808 =  ( n698 ) ? ( bv_8_54_n651 ) : ( n807 ) ;
assign n809 =  ( n696 ) ? ( bv_8_63_n629 ) : ( n808 ) ;
assign n810 =  ( n694 ) ? ( bv_8_247_n37 ) : ( n809 ) ;
assign n811 =  ( n691 ) ? ( bv_8_204_n201 ) : ( n810 ) ;
assign n812 =  ( n689 ) ? ( bv_8_52_n657 ) : ( n811 ) ;
assign n813 =  ( n687 ) ? ( bv_8_165_n333 ) : ( n812 ) ;
assign n814 =  ( n685 ) ? ( bv_8_229_n107 ) : ( n813 ) ;
assign n815 =  ( n683 ) ? ( bv_8_241_n61 ) : ( n814 ) ;
assign n816 =  ( n680 ) ? ( bv_8_113_n495 ) : ( n815 ) ;
assign n817 =  ( n678 ) ? ( bv_8_216_n155 ) : ( n816 ) ;
assign n818 =  ( n676 ) ? ( bv_8_49_n666 ) : ( n817 ) ;
assign n819 =  ( n673 ) ? ( bv_8_21_n674 ) : ( n818 ) ;
assign n820 =  ( n670 ) ? ( bv_8_4_n671 ) : ( n819 ) ;
assign n821 =  ( n667 ) ? ( bv_8_199_n219 ) : ( n820 ) ;
assign n822 =  ( n663 ) ? ( bv_8_35_n664 ) : ( n821 ) ;
assign n823 =  ( n661 ) ? ( bv_8_195_n234 ) : ( n822 ) ;
assign n824 =  ( n658 ) ? ( bv_8_24_n659 ) : ( n823 ) ;
assign n825 =  ( n655 ) ? ( bv_8_150_n383 ) : ( n824 ) ;
assign n826 =  ( n652 ) ? ( bv_8_5_n653 ) : ( n825 ) ;
assign n827 =  ( n649 ) ? ( bv_8_154_n371 ) : ( n826 ) ;
assign n828 =  ( n646 ) ? ( bv_8_7_n647 ) : ( n827 ) ;
assign n829 =  ( n643 ) ? ( bv_8_18_n644 ) : ( n828 ) ;
assign n830 =  ( n641 ) ? ( bv_8_128_n452 ) : ( n829 ) ;
assign n831 =  ( n639 ) ? ( bv_8_226_n119 ) : ( n830 ) ;
assign n832 =  ( n637 ) ? ( bv_8_235_n85 ) : ( n831 ) ;
assign n833 =  ( n634 ) ? ( bv_8_39_n635 ) : ( n832 ) ;
assign n834 =  ( n632 ) ? ( bv_8_178_n291 ) : ( n833 ) ;
assign n835 =  ( n630 ) ? ( bv_8_117_n484 ) : ( n834 ) ;
assign n836 =  ( n626 ) ? ( bv_8_9_n627 ) : ( n835 ) ;
assign n837 =  ( n624 ) ? ( bv_8_131_n442 ) : ( n836 ) ;
assign n838 =  ( n621 ) ? ( bv_8_44_n622 ) : ( n837 ) ;
assign n839 =  ( n618 ) ? ( bv_8_26_n619 ) : ( n838 ) ;
assign n840 =  ( n615 ) ? ( bv_8_27_n616 ) : ( n839 ) ;
assign n841 =  ( n613 ) ? ( bv_8_110_n504 ) : ( n840 ) ;
assign n842 =  ( n611 ) ? ( bv_8_90_n561 ) : ( n841 ) ;
assign n843 =  ( n609 ) ? ( bv_8_160_n352 ) : ( n842 ) ;
assign n844 =  ( n606 ) ? ( bv_8_82_n581 ) : ( n843 ) ;
assign n845 =  ( n603 ) ? ( bv_8_59_n604 ) : ( n844 ) ;
assign n846 =  ( n601 ) ? ( bv_8_214_n163 ) : ( n845 ) ;
assign n847 =  ( n599 ) ? ( bv_8_179_n287 ) : ( n846 ) ;
assign n848 =  ( n596 ) ? ( bv_8_41_n597 ) : ( n847 ) ;
assign n849 =  ( n594 ) ? ( bv_8_227_n115 ) : ( n848 ) ;
assign n850 =  ( n591 ) ? ( bv_8_47_n592 ) : ( n849 ) ;
assign n851 =  ( n589 ) ? ( bv_8_132_n438 ) : ( n850 ) ;
assign n852 =  ( n587 ) ? ( bv_8_83_n578 ) : ( n851 ) ;
assign n853 =  ( n585 ) ? ( bv_8_209_n182 ) : ( n852 ) ;
assign n854 =  ( n582 ) ? ( bv_8_0_n583 ) : ( n853 ) ;
assign n855 =  ( n579 ) ? ( bv_8_237_n77 ) : ( n854 ) ;
assign n856 =  ( n575 ) ? ( bv_8_32_n576 ) : ( n855 ) ;
assign n857 =  ( n573 ) ? ( bv_8_252_n17 ) : ( n856 ) ;
assign n858 =  ( n571 ) ? ( bv_8_177_n295 ) : ( n857 ) ;
assign n859 =  ( n569 ) ? ( bv_8_91_n557 ) : ( n858 ) ;
assign n860 =  ( n567 ) ? ( bv_8_106_n516 ) : ( n859 ) ;
assign n861 =  ( n565 ) ? ( bv_8_203_n205 ) : ( n860 ) ;
assign n862 =  ( n562 ) ? ( bv_8_190_n252 ) : ( n861 ) ;
assign n863 =  ( n558 ) ? ( bv_8_57_n559 ) : ( n862 ) ;
assign n864 =  ( n554 ) ? ( bv_8_74_n555 ) : ( n863 ) ;
assign n865 =  ( n551 ) ? ( bv_8_76_n552 ) : ( n864 ) ;
assign n866 =  ( n548 ) ? ( bv_8_88_n549 ) : ( n865 ) ;
assign n867 =  ( n546 ) ? ( bv_8_207_n190 ) : ( n866 ) ;
assign n868 =  ( n544 ) ? ( bv_8_208_n186 ) : ( n867 ) ;
assign n869 =  ( n542 ) ? ( bv_8_239_n69 ) : ( n868 ) ;
assign n870 =  ( n540 ) ? ( bv_8_170_n318 ) : ( n869 ) ;
assign n871 =  ( n538 ) ? ( bv_8_251_n21 ) : ( n870 ) ;
assign n872 =  ( n534 ) ? ( bv_8_67_n535 ) : ( n871 ) ;
assign n873 =  ( n531 ) ? ( bv_8_77_n532 ) : ( n872 ) ;
assign n874 =  ( n528 ) ? ( bv_8_51_n529 ) : ( n873 ) ;
assign n875 =  ( n526 ) ? ( bv_8_133_n435 ) : ( n874 ) ;
assign n876 =  ( n522 ) ? ( bv_8_69_n523 ) : ( n875 ) ;
assign n877 =  ( n520 ) ? ( bv_8_249_n29 ) : ( n876 ) ;
assign n878 =  ( n517 ) ? ( bv_8_2_n518 ) : ( n877 ) ;
assign n879 =  ( n514 ) ? ( bv_8_127_n455 ) : ( n878 ) ;
assign n880 =  ( n510 ) ? ( bv_8_80_n511 ) : ( n879 ) ;
assign n881 =  ( n507 ) ? ( bv_8_60_n508 ) : ( n880 ) ;
assign n882 =  ( n505 ) ? ( bv_8_159_n355 ) : ( n881 ) ;
assign n883 =  ( n502 ) ? ( bv_8_168_n323 ) : ( n882 ) ;
assign n884 =  ( n498 ) ? ( bv_8_81_n499 ) : ( n883 ) ;
assign n885 =  ( n496 ) ? ( bv_8_163_n341 ) : ( n884 ) ;
assign n886 =  ( n492 ) ? ( bv_8_64_n493 ) : ( n885 ) ;
assign n887 =  ( n489 ) ? ( bv_8_143_n406 ) : ( n886 ) ;
assign n888 =  ( n487 ) ? ( bv_8_146_n396 ) : ( n887 ) ;
assign n889 =  ( n485 ) ? ( bv_8_157_n361 ) : ( n888 ) ;
assign n890 =  ( n481 ) ? ( bv_8_56_n482 ) : ( n889 ) ;
assign n891 =  ( n478 ) ? ( bv_8_245_n45 ) : ( n890 ) ;
assign n892 =  ( n475 ) ? ( bv_8_188_n259 ) : ( n891 ) ;
assign n893 =  ( n473 ) ? ( bv_8_182_n278 ) : ( n892 ) ;
assign n894 =  ( n471 ) ? ( bv_8_218_n148 ) : ( n893 ) ;
assign n895 =  ( n468 ) ? ( bv_8_33_n469 ) : ( n894 ) ;
assign n896 =  ( n464 ) ? ( bv_8_16_n465 ) : ( n895 ) ;
assign n897 =  ( n461 ) ? ( bv_8_255_n5 ) : ( n896 ) ;
assign n898 =  ( n458 ) ? ( bv_8_243_n53 ) : ( n897 ) ;
assign n899 =  ( n456 ) ? ( bv_8_210_n178 ) : ( n898 ) ;
assign n900 =  ( n453 ) ? ( bv_8_205_n197 ) : ( n899 ) ;
assign n901 =  ( n449 ) ? ( bv_8_12_n450 ) : ( n900 ) ;
assign n902 =  ( n446 ) ? ( bv_8_19_n447 ) : ( n901 ) ;
assign n903 =  ( n443 ) ? ( bv_8_236_n81 ) : ( n902 ) ;
assign n904 =  ( n439 ) ? ( bv_8_95_n440 ) : ( n903 ) ;
assign n905 =  ( n436 ) ? ( bv_8_151_n379 ) : ( n904 ) ;
assign n906 =  ( n432 ) ? ( bv_8_68_n433 ) : ( n905 ) ;
assign n907 =  ( n429 ) ? ( bv_8_23_n430 ) : ( n906 ) ;
assign n908 =  ( n427 ) ? ( bv_8_196_n230 ) : ( n907 ) ;
assign n909 =  ( n425 ) ? ( bv_8_167_n326 ) : ( n908 ) ;
assign n910 =  ( n422 ) ? ( bv_8_126_n423 ) : ( n909 ) ;
assign n911 =  ( n419 ) ? ( bv_8_61_n420 ) : ( n910 ) ;
assign n912 =  ( n416 ) ? ( bv_8_100_n417 ) : ( n911 ) ;
assign n913 =  ( n413 ) ? ( bv_8_93_n414 ) : ( n912 ) ;
assign n914 =  ( n410 ) ? ( bv_8_25_n411 ) : ( n913 ) ;
assign n915 =  ( n407 ) ? ( bv_8_115_n408 ) : ( n914 ) ;
assign n916 =  ( n403 ) ? ( bv_8_96_n404 ) : ( n915 ) ;
assign n917 =  ( n400 ) ? ( bv_8_129_n401 ) : ( n916 ) ;
assign n918 =  ( n397 ) ? ( bv_8_79_n398 ) : ( n917 ) ;
assign n919 =  ( n394 ) ? ( bv_8_220_n140 ) : ( n918 ) ;
assign n920 =  ( n390 ) ? ( bv_8_34_n391 ) : ( n919 ) ;
assign n921 =  ( n387 ) ? ( bv_8_42_n388 ) : ( n920 ) ;
assign n922 =  ( n384 ) ? ( bv_8_144_n385 ) : ( n921 ) ;
assign n923 =  ( n380 ) ? ( bv_8_136_n381 ) : ( n922 ) ;
assign n924 =  ( n376 ) ? ( bv_8_70_n377 ) : ( n923 ) ;
assign n925 =  ( n374 ) ? ( bv_8_238_n73 ) : ( n924 ) ;
assign n926 =  ( n372 ) ? ( bv_8_184_n270 ) : ( n925 ) ;
assign n927 =  ( n368 ) ? ( bv_8_20_n369 ) : ( n926 ) ;
assign n928 =  ( n366 ) ? ( bv_8_222_n132 ) : ( n927 ) ;
assign n929 =  ( n362 ) ? ( bv_8_94_n363 ) : ( n928 ) ;
assign n930 =  ( n358 ) ? ( bv_8_11_n359 ) : ( n929 ) ;
assign n931 =  ( n356 ) ? ( bv_8_219_n144 ) : ( n930 ) ;
assign n932 =  ( n353 ) ? ( bv_8_224_n126 ) : ( n931 ) ;
assign n933 =  ( n349 ) ? ( bv_8_50_n350 ) : ( n932 ) ;
assign n934 =  ( n346 ) ? ( bv_8_58_n347 ) : ( n933 ) ;
assign n935 =  ( n342 ) ? ( bv_8_10_n343 ) : ( n934 ) ;
assign n936 =  ( n338 ) ? ( bv_8_73_n339 ) : ( n935 ) ;
assign n937 =  ( n334 ) ? ( bv_8_6_n335 ) : ( n936 ) ;
assign n938 =  ( n330 ) ? ( bv_8_36_n331 ) : ( n937 ) ;
assign n939 =  ( n327 ) ? ( bv_8_92_n328 ) : ( n938 ) ;
assign n940 =  ( n324 ) ? ( bv_8_194_n238 ) : ( n939 ) ;
assign n941 =  ( n321 ) ? ( bv_8_211_n174 ) : ( n940 ) ;
assign n942 =  ( n319 ) ? ( bv_8_172_n310 ) : ( n941 ) ;
assign n943 =  ( n315 ) ? ( bv_8_98_n316 ) : ( n942 ) ;
assign n944 =  ( n311 ) ? ( bv_8_145_n312 ) : ( n943 ) ;
assign n945 =  ( n307 ) ? ( bv_8_149_n308 ) : ( n944 ) ;
assign n946 =  ( n304 ) ? ( bv_8_228_n111 ) : ( n945 ) ;
assign n947 =  ( n301 ) ? ( bv_8_121_n302 ) : ( n946 ) ;
assign n948 =  ( n298 ) ? ( bv_8_231_n100 ) : ( n947 ) ;
assign n949 =  ( n296 ) ? ( bv_8_200_n216 ) : ( n948 ) ;
assign n950 =  ( n292 ) ? ( bv_8_55_n293 ) : ( n949 ) ;
assign n951 =  ( n288 ) ? ( bv_8_109_n289 ) : ( n950 ) ;
assign n952 =  ( n284 ) ? ( bv_8_141_n285 ) : ( n951 ) ;
assign n953 =  ( n282 ) ? ( bv_8_213_n166 ) : ( n952 ) ;
assign n954 =  ( n279 ) ? ( bv_8_78_n280 ) : ( n953 ) ;
assign n955 =  ( n275 ) ? ( bv_8_169_n276 ) : ( n954 ) ;
assign n956 =  ( n271 ) ? ( bv_8_108_n272 ) : ( n955 ) ;
assign n957 =  ( n267 ) ? ( bv_8_86_n268 ) : ( n956 ) ;
assign n958 =  ( n265 ) ? ( bv_8_244_n49 ) : ( n957 ) ;
assign n959 =  ( n263 ) ? ( bv_8_234_n89 ) : ( n958 ) ;
assign n960 =  ( n260 ) ? ( bv_8_101_n261 ) : ( n959 ) ;
assign n961 =  ( n256 ) ? ( bv_8_122_n257 ) : ( n960 ) ;
assign n962 =  ( n253 ) ? ( bv_8_174_n254 ) : ( n961 ) ;
assign n963 =  ( n249 ) ? ( bv_8_8_n250 ) : ( n962 ) ;
assign n964 =  ( n246 ) ? ( bv_8_186_n247 ) : ( n963 ) ;
assign n965 =  ( n242 ) ? ( bv_8_120_n243 ) : ( n964 ) ;
assign n966 =  ( n239 ) ? ( bv_8_37_n240 ) : ( n965 ) ;
assign n967 =  ( n235 ) ? ( bv_8_46_n236 ) : ( n966 ) ;
assign n968 =  ( n231 ) ? ( bv_8_28_n232 ) : ( n967 ) ;
assign n969 =  ( n227 ) ? ( bv_8_166_n228 ) : ( n968 ) ;
assign n970 =  ( n223 ) ? ( bv_8_180_n224 ) : ( n969 ) ;
assign n971 =  ( n220 ) ? ( bv_8_198_n221 ) : ( n970 ) ;
assign n972 =  ( n217 ) ? ( bv_8_232_n96 ) : ( n971 ) ;
assign n973 =  ( n214 ) ? ( bv_8_221_n136 ) : ( n972 ) ;
assign n974 =  ( n210 ) ? ( bv_8_116_n211 ) : ( n973 ) ;
assign n975 =  ( n206 ) ? ( bv_8_31_n207 ) : ( n974 ) ;
assign n976 =  ( n202 ) ? ( bv_8_75_n203 ) : ( n975 ) ;
assign n977 =  ( n198 ) ? ( bv_8_189_n199 ) : ( n976 ) ;
assign n978 =  ( n194 ) ? ( bv_8_139_n195 ) : ( n977 ) ;
assign n979 =  ( n191 ) ? ( bv_8_138_n192 ) : ( n978 ) ;
assign n980 =  ( n187 ) ? ( bv_8_112_n188 ) : ( n979 ) ;
assign n981 =  ( n183 ) ? ( bv_8_62_n184 ) : ( n980 ) ;
assign n982 =  ( n179 ) ? ( bv_8_181_n180 ) : ( n981 ) ;
assign n983 =  ( n175 ) ? ( bv_8_102_n176 ) : ( n982 ) ;
assign n984 =  ( n171 ) ? ( bv_8_72_n172 ) : ( n983 ) ;
assign n985 =  ( n167 ) ? ( bv_8_3_n168 ) : ( n984 ) ;
assign n986 =  ( n164 ) ? ( bv_8_246_n41 ) : ( n985 ) ;
assign n987 =  ( n160 ) ? ( bv_8_14_n161 ) : ( n986 ) ;
assign n988 =  ( n156 ) ? ( bv_8_97_n157 ) : ( n987 ) ;
assign n989 =  ( n152 ) ? ( bv_8_53_n153 ) : ( n988 ) ;
assign n990 =  ( n149 ) ? ( bv_8_87_n150 ) : ( n989 ) ;
assign n991 =  ( n145 ) ? ( bv_8_185_n146 ) : ( n990 ) ;
assign n992 =  ( n141 ) ? ( bv_8_134_n142 ) : ( n991 ) ;
assign n993 =  ( n137 ) ? ( bv_8_193_n138 ) : ( n992 ) ;
assign n994 =  ( n133 ) ? ( bv_8_29_n134 ) : ( n993 ) ;
assign n995 =  ( n129 ) ? ( bv_8_158_n130 ) : ( n994 ) ;
assign n996 =  ( n127 ) ? ( bv_8_225_n123 ) : ( n995 ) ;
assign n997 =  ( n124 ) ? ( bv_8_248_n33 ) : ( n996 ) ;
assign n998 =  ( n120 ) ? ( bv_8_152_n121 ) : ( n997 ) ;
assign n999 =  ( n116 ) ? ( bv_8_17_n117 ) : ( n998 ) ;
assign n1000 =  ( n112 ) ? ( bv_8_105_n113 ) : ( n999 ) ;
assign n1001 =  ( n108 ) ? ( bv_8_217_n109 ) : ( n1000 ) ;
assign n1002 =  ( n104 ) ? ( bv_8_142_n105 ) : ( n1001 ) ;
assign n1003 =  ( n101 ) ? ( bv_8_148_n102 ) : ( n1002 ) ;
assign n1004 =  ( n97 ) ? ( bv_8_155_n98 ) : ( n1003 ) ;
assign n1005 =  ( n93 ) ? ( bv_8_30_n94 ) : ( n1004 ) ;
assign n1006 =  ( n90 ) ? ( bv_8_135_n91 ) : ( n1005 ) ;
assign n1007 =  ( n86 ) ? ( bv_8_233_n87 ) : ( n1006 ) ;
assign n1008 =  ( n82 ) ? ( bv_8_206_n83 ) : ( n1007 ) ;
assign n1009 =  ( n78 ) ? ( bv_8_85_n79 ) : ( n1008 ) ;
assign n1010 =  ( n74 ) ? ( bv_8_40_n75 ) : ( n1009 ) ;
assign n1011 =  ( n70 ) ? ( bv_8_223_n71 ) : ( n1010 ) ;
assign n1012 =  ( n66 ) ? ( bv_8_140_n67 ) : ( n1011 ) ;
assign n1013 =  ( n62 ) ? ( bv_8_161_n63 ) : ( n1012 ) ;
assign n1014 =  ( n58 ) ? ( bv_8_137_n59 ) : ( n1013 ) ;
assign n1015 =  ( n54 ) ? ( bv_8_13_n55 ) : ( n1014 ) ;
assign n1016 =  ( n50 ) ? ( bv_8_191_n51 ) : ( n1015 ) ;
assign n1017 =  ( n46 ) ? ( bv_8_230_n47 ) : ( n1016 ) ;
assign n1018 =  ( n42 ) ? ( bv_8_66_n43 ) : ( n1017 ) ;
assign n1019 =  ( n38 ) ? ( bv_8_104_n39 ) : ( n1018 ) ;
assign n1020 =  ( n34 ) ? ( bv_8_65_n35 ) : ( n1019 ) ;
assign n1021 =  ( n30 ) ? ( bv_8_153_n31 ) : ( n1020 ) ;
assign n1022 =  ( n26 ) ? ( bv_8_45_n27 ) : ( n1021 ) ;
assign n1023 =  ( n22 ) ? ( bv_8_15_n23 ) : ( n1022 ) ;
assign n1024 =  ( n18 ) ? ( bv_8_176_n19 ) : ( n1023 ) ;
assign n1025 =  ( n14 ) ? ( bv_8_84_n15 ) : ( n1024 ) ;
assign n1026 =  ( n10 ) ? ( bv_8_187_n11 ) : ( n1025 ) ;
assign n1027 =  ( n6 ) ? ( bv_8_22_n7 ) : ( n1026 ) ;
assign n1028 =  ( n3 ) ^ ( n1027 )  ;
assign n1029 = in[119:112] ;
assign n1030 = in[15:8] ;
assign n1031 =  ( n1030 ) == ( bv_8_255_n5 )  ;
assign n1032 = in[15:8] ;
assign n1033 =  ( n1032 ) == ( bv_8_254_n9 )  ;
assign n1034 = in[15:8] ;
assign n1035 =  ( n1034 ) == ( bv_8_253_n13 )  ;
assign n1036 = in[15:8] ;
assign n1037 =  ( n1036 ) == ( bv_8_252_n17 )  ;
assign n1038 = in[15:8] ;
assign n1039 =  ( n1038 ) == ( bv_8_251_n21 )  ;
assign n1040 = in[15:8] ;
assign n1041 =  ( n1040 ) == ( bv_8_250_n25 )  ;
assign n1042 = in[15:8] ;
assign n1043 =  ( n1042 ) == ( bv_8_249_n29 )  ;
assign n1044 = in[15:8] ;
assign n1045 =  ( n1044 ) == ( bv_8_248_n33 )  ;
assign n1046 = in[15:8] ;
assign n1047 =  ( n1046 ) == ( bv_8_247_n37 )  ;
assign n1048 = in[15:8] ;
assign n1049 =  ( n1048 ) == ( bv_8_246_n41 )  ;
assign n1050 = in[15:8] ;
assign n1051 =  ( n1050 ) == ( bv_8_245_n45 )  ;
assign n1052 = in[15:8] ;
assign n1053 =  ( n1052 ) == ( bv_8_244_n49 )  ;
assign n1054 = in[15:8] ;
assign n1055 =  ( n1054 ) == ( bv_8_243_n53 )  ;
assign n1056 = in[15:8] ;
assign n1057 =  ( n1056 ) == ( bv_8_242_n57 )  ;
assign n1058 = in[15:8] ;
assign n1059 =  ( n1058 ) == ( bv_8_241_n61 )  ;
assign n1060 = in[15:8] ;
assign n1061 =  ( n1060 ) == ( bv_8_240_n65 )  ;
assign n1062 = in[15:8] ;
assign n1063 =  ( n1062 ) == ( bv_8_239_n69 )  ;
assign n1064 = in[15:8] ;
assign n1065 =  ( n1064 ) == ( bv_8_238_n73 )  ;
assign n1066 = in[15:8] ;
assign n1067 =  ( n1066 ) == ( bv_8_237_n77 )  ;
assign n1068 = in[15:8] ;
assign n1069 =  ( n1068 ) == ( bv_8_236_n81 )  ;
assign n1070 = in[15:8] ;
assign n1071 =  ( n1070 ) == ( bv_8_235_n85 )  ;
assign n1072 = in[15:8] ;
assign n1073 =  ( n1072 ) == ( bv_8_234_n89 )  ;
assign n1074 = in[15:8] ;
assign n1075 =  ( n1074 ) == ( bv_8_233_n87 )  ;
assign n1076 = in[15:8] ;
assign n1077 =  ( n1076 ) == ( bv_8_232_n96 )  ;
assign n1078 = in[15:8] ;
assign n1079 =  ( n1078 ) == ( bv_8_231_n100 )  ;
assign n1080 = in[15:8] ;
assign n1081 =  ( n1080 ) == ( bv_8_230_n47 )  ;
assign n1082 = in[15:8] ;
assign n1083 =  ( n1082 ) == ( bv_8_229_n107 )  ;
assign n1084 = in[15:8] ;
assign n1085 =  ( n1084 ) == ( bv_8_228_n111 )  ;
assign n1086 = in[15:8] ;
assign n1087 =  ( n1086 ) == ( bv_8_227_n115 )  ;
assign n1088 = in[15:8] ;
assign n1089 =  ( n1088 ) == ( bv_8_226_n119 )  ;
assign n1090 = in[15:8] ;
assign n1091 =  ( n1090 ) == ( bv_8_225_n123 )  ;
assign n1092 = in[15:8] ;
assign n1093 =  ( n1092 ) == ( bv_8_224_n126 )  ;
assign n1094 = in[15:8] ;
assign n1095 =  ( n1094 ) == ( bv_8_223_n71 )  ;
assign n1096 = in[15:8] ;
assign n1097 =  ( n1096 ) == ( bv_8_222_n132 )  ;
assign n1098 = in[15:8] ;
assign n1099 =  ( n1098 ) == ( bv_8_221_n136 )  ;
assign n1100 = in[15:8] ;
assign n1101 =  ( n1100 ) == ( bv_8_220_n140 )  ;
assign n1102 = in[15:8] ;
assign n1103 =  ( n1102 ) == ( bv_8_219_n144 )  ;
assign n1104 = in[15:8] ;
assign n1105 =  ( n1104 ) == ( bv_8_218_n148 )  ;
assign n1106 = in[15:8] ;
assign n1107 =  ( n1106 ) == ( bv_8_217_n109 )  ;
assign n1108 = in[15:8] ;
assign n1109 =  ( n1108 ) == ( bv_8_216_n155 )  ;
assign n1110 = in[15:8] ;
assign n1111 =  ( n1110 ) == ( bv_8_215_n159 )  ;
assign n1112 = in[15:8] ;
assign n1113 =  ( n1112 ) == ( bv_8_214_n163 )  ;
assign n1114 = in[15:8] ;
assign n1115 =  ( n1114 ) == ( bv_8_213_n166 )  ;
assign n1116 = in[15:8] ;
assign n1117 =  ( n1116 ) == ( bv_8_212_n170 )  ;
assign n1118 = in[15:8] ;
assign n1119 =  ( n1118 ) == ( bv_8_211_n174 )  ;
assign n1120 = in[15:8] ;
assign n1121 =  ( n1120 ) == ( bv_8_210_n178 )  ;
assign n1122 = in[15:8] ;
assign n1123 =  ( n1122 ) == ( bv_8_209_n182 )  ;
assign n1124 = in[15:8] ;
assign n1125 =  ( n1124 ) == ( bv_8_208_n186 )  ;
assign n1126 = in[15:8] ;
assign n1127 =  ( n1126 ) == ( bv_8_207_n190 )  ;
assign n1128 = in[15:8] ;
assign n1129 =  ( n1128 ) == ( bv_8_206_n83 )  ;
assign n1130 = in[15:8] ;
assign n1131 =  ( n1130 ) == ( bv_8_205_n197 )  ;
assign n1132 = in[15:8] ;
assign n1133 =  ( n1132 ) == ( bv_8_204_n201 )  ;
assign n1134 = in[15:8] ;
assign n1135 =  ( n1134 ) == ( bv_8_203_n205 )  ;
assign n1136 = in[15:8] ;
assign n1137 =  ( n1136 ) == ( bv_8_202_n209 )  ;
assign n1138 = in[15:8] ;
assign n1139 =  ( n1138 ) == ( bv_8_201_n213 )  ;
assign n1140 = in[15:8] ;
assign n1141 =  ( n1140 ) == ( bv_8_200_n216 )  ;
assign n1142 = in[15:8] ;
assign n1143 =  ( n1142 ) == ( bv_8_199_n219 )  ;
assign n1144 = in[15:8] ;
assign n1145 =  ( n1144 ) == ( bv_8_198_n221 )  ;
assign n1146 = in[15:8] ;
assign n1147 =  ( n1146 ) == ( bv_8_197_n226 )  ;
assign n1148 = in[15:8] ;
assign n1149 =  ( n1148 ) == ( bv_8_196_n230 )  ;
assign n1150 = in[15:8] ;
assign n1151 =  ( n1150 ) == ( bv_8_195_n234 )  ;
assign n1152 = in[15:8] ;
assign n1153 =  ( n1152 ) == ( bv_8_194_n238 )  ;
assign n1154 = in[15:8] ;
assign n1155 =  ( n1154 ) == ( bv_8_193_n138 )  ;
assign n1156 = in[15:8] ;
assign n1157 =  ( n1156 ) == ( bv_8_192_n245 )  ;
assign n1158 = in[15:8] ;
assign n1159 =  ( n1158 ) == ( bv_8_191_n51 )  ;
assign n1160 = in[15:8] ;
assign n1161 =  ( n1160 ) == ( bv_8_190_n252 )  ;
assign n1162 = in[15:8] ;
assign n1163 =  ( n1162 ) == ( bv_8_189_n199 )  ;
assign n1164 = in[15:8] ;
assign n1165 =  ( n1164 ) == ( bv_8_188_n259 )  ;
assign n1166 = in[15:8] ;
assign n1167 =  ( n1166 ) == ( bv_8_187_n11 )  ;
assign n1168 = in[15:8] ;
assign n1169 =  ( n1168 ) == ( bv_8_186_n247 )  ;
assign n1170 = in[15:8] ;
assign n1171 =  ( n1170 ) == ( bv_8_185_n146 )  ;
assign n1172 = in[15:8] ;
assign n1173 =  ( n1172 ) == ( bv_8_184_n270 )  ;
assign n1174 = in[15:8] ;
assign n1175 =  ( n1174 ) == ( bv_8_183_n274 )  ;
assign n1176 = in[15:8] ;
assign n1177 =  ( n1176 ) == ( bv_8_182_n278 )  ;
assign n1178 = in[15:8] ;
assign n1179 =  ( n1178 ) == ( bv_8_181_n180 )  ;
assign n1180 = in[15:8] ;
assign n1181 =  ( n1180 ) == ( bv_8_180_n224 )  ;
assign n1182 = in[15:8] ;
assign n1183 =  ( n1182 ) == ( bv_8_179_n287 )  ;
assign n1184 = in[15:8] ;
assign n1185 =  ( n1184 ) == ( bv_8_178_n291 )  ;
assign n1186 = in[15:8] ;
assign n1187 =  ( n1186 ) == ( bv_8_177_n295 )  ;
assign n1188 = in[15:8] ;
assign n1189 =  ( n1188 ) == ( bv_8_176_n19 )  ;
assign n1190 = in[15:8] ;
assign n1191 =  ( n1190 ) == ( bv_8_175_n300 )  ;
assign n1192 = in[15:8] ;
assign n1193 =  ( n1192 ) == ( bv_8_174_n254 )  ;
assign n1194 = in[15:8] ;
assign n1195 =  ( n1194 ) == ( bv_8_173_n306 )  ;
assign n1196 = in[15:8] ;
assign n1197 =  ( n1196 ) == ( bv_8_172_n310 )  ;
assign n1198 = in[15:8] ;
assign n1199 =  ( n1198 ) == ( bv_8_171_n314 )  ;
assign n1200 = in[15:8] ;
assign n1201 =  ( n1200 ) == ( bv_8_170_n318 )  ;
assign n1202 = in[15:8] ;
assign n1203 =  ( n1202 ) == ( bv_8_169_n276 )  ;
assign n1204 = in[15:8] ;
assign n1205 =  ( n1204 ) == ( bv_8_168_n323 )  ;
assign n1206 = in[15:8] ;
assign n1207 =  ( n1206 ) == ( bv_8_167_n326 )  ;
assign n1208 = in[15:8] ;
assign n1209 =  ( n1208 ) == ( bv_8_166_n228 )  ;
assign n1210 = in[15:8] ;
assign n1211 =  ( n1210 ) == ( bv_8_165_n333 )  ;
assign n1212 = in[15:8] ;
assign n1213 =  ( n1212 ) == ( bv_8_164_n337 )  ;
assign n1214 = in[15:8] ;
assign n1215 =  ( n1214 ) == ( bv_8_163_n341 )  ;
assign n1216 = in[15:8] ;
assign n1217 =  ( n1216 ) == ( bv_8_162_n345 )  ;
assign n1218 = in[15:8] ;
assign n1219 =  ( n1218 ) == ( bv_8_161_n63 )  ;
assign n1220 = in[15:8] ;
assign n1221 =  ( n1220 ) == ( bv_8_160_n352 )  ;
assign n1222 = in[15:8] ;
assign n1223 =  ( n1222 ) == ( bv_8_159_n355 )  ;
assign n1224 = in[15:8] ;
assign n1225 =  ( n1224 ) == ( bv_8_158_n130 )  ;
assign n1226 = in[15:8] ;
assign n1227 =  ( n1226 ) == ( bv_8_157_n361 )  ;
assign n1228 = in[15:8] ;
assign n1229 =  ( n1228 ) == ( bv_8_156_n365 )  ;
assign n1230 = in[15:8] ;
assign n1231 =  ( n1230 ) == ( bv_8_155_n98 )  ;
assign n1232 = in[15:8] ;
assign n1233 =  ( n1232 ) == ( bv_8_154_n371 )  ;
assign n1234 = in[15:8] ;
assign n1235 =  ( n1234 ) == ( bv_8_153_n31 )  ;
assign n1236 = in[15:8] ;
assign n1237 =  ( n1236 ) == ( bv_8_152_n121 )  ;
assign n1238 = in[15:8] ;
assign n1239 =  ( n1238 ) == ( bv_8_151_n379 )  ;
assign n1240 = in[15:8] ;
assign n1241 =  ( n1240 ) == ( bv_8_150_n383 )  ;
assign n1242 = in[15:8] ;
assign n1243 =  ( n1242 ) == ( bv_8_149_n308 )  ;
assign n1244 = in[15:8] ;
assign n1245 =  ( n1244 ) == ( bv_8_148_n102 )  ;
assign n1246 = in[15:8] ;
assign n1247 =  ( n1246 ) == ( bv_8_147_n393 )  ;
assign n1248 = in[15:8] ;
assign n1249 =  ( n1248 ) == ( bv_8_146_n396 )  ;
assign n1250 = in[15:8] ;
assign n1251 =  ( n1250 ) == ( bv_8_145_n312 )  ;
assign n1252 = in[15:8] ;
assign n1253 =  ( n1252 ) == ( bv_8_144_n385 )  ;
assign n1254 = in[15:8] ;
assign n1255 =  ( n1254 ) == ( bv_8_143_n406 )  ;
assign n1256 = in[15:8] ;
assign n1257 =  ( n1256 ) == ( bv_8_142_n105 )  ;
assign n1258 = in[15:8] ;
assign n1259 =  ( n1258 ) == ( bv_8_141_n285 )  ;
assign n1260 = in[15:8] ;
assign n1261 =  ( n1260 ) == ( bv_8_140_n67 )  ;
assign n1262 = in[15:8] ;
assign n1263 =  ( n1262 ) == ( bv_8_139_n195 )  ;
assign n1264 = in[15:8] ;
assign n1265 =  ( n1264 ) == ( bv_8_138_n192 )  ;
assign n1266 = in[15:8] ;
assign n1267 =  ( n1266 ) == ( bv_8_137_n59 )  ;
assign n1268 = in[15:8] ;
assign n1269 =  ( n1268 ) == ( bv_8_136_n381 )  ;
assign n1270 = in[15:8] ;
assign n1271 =  ( n1270 ) == ( bv_8_135_n91 )  ;
assign n1272 = in[15:8] ;
assign n1273 =  ( n1272 ) == ( bv_8_134_n142 )  ;
assign n1274 = in[15:8] ;
assign n1275 =  ( n1274 ) == ( bv_8_133_n435 )  ;
assign n1276 = in[15:8] ;
assign n1277 =  ( n1276 ) == ( bv_8_132_n438 )  ;
assign n1278 = in[15:8] ;
assign n1279 =  ( n1278 ) == ( bv_8_131_n442 )  ;
assign n1280 = in[15:8] ;
assign n1281 =  ( n1280 ) == ( bv_8_130_n445 )  ;
assign n1282 = in[15:8] ;
assign n1283 =  ( n1282 ) == ( bv_8_129_n401 )  ;
assign n1284 = in[15:8] ;
assign n1285 =  ( n1284 ) == ( bv_8_128_n452 )  ;
assign n1286 = in[15:8] ;
assign n1287 =  ( n1286 ) == ( bv_8_127_n455 )  ;
assign n1288 = in[15:8] ;
assign n1289 =  ( n1288 ) == ( bv_8_126_n423 )  ;
assign n1290 = in[15:8] ;
assign n1291 =  ( n1290 ) == ( bv_8_125_n460 )  ;
assign n1292 = in[15:8] ;
assign n1293 =  ( n1292 ) == ( bv_8_124_n463 )  ;
assign n1294 = in[15:8] ;
assign n1295 =  ( n1294 ) == ( bv_8_123_n467 )  ;
assign n1296 = in[15:8] ;
assign n1297 =  ( n1296 ) == ( bv_8_122_n257 )  ;
assign n1298 = in[15:8] ;
assign n1299 =  ( n1298 ) == ( bv_8_121_n302 )  ;
assign n1300 = in[15:8] ;
assign n1301 =  ( n1300 ) == ( bv_8_120_n243 )  ;
assign n1302 = in[15:8] ;
assign n1303 =  ( n1302 ) == ( bv_8_119_n477 )  ;
assign n1304 = in[15:8] ;
assign n1305 =  ( n1304 ) == ( bv_8_118_n480 )  ;
assign n1306 = in[15:8] ;
assign n1307 =  ( n1306 ) == ( bv_8_117_n484 )  ;
assign n1308 = in[15:8] ;
assign n1309 =  ( n1308 ) == ( bv_8_116_n211 )  ;
assign n1310 = in[15:8] ;
assign n1311 =  ( n1310 ) == ( bv_8_115_n408 )  ;
assign n1312 = in[15:8] ;
assign n1313 =  ( n1312 ) == ( bv_8_114_n491 )  ;
assign n1314 = in[15:8] ;
assign n1315 =  ( n1314 ) == ( bv_8_113_n495 )  ;
assign n1316 = in[15:8] ;
assign n1317 =  ( n1316 ) == ( bv_8_112_n188 )  ;
assign n1318 = in[15:8] ;
assign n1319 =  ( n1318 ) == ( bv_8_111_n501 )  ;
assign n1320 = in[15:8] ;
assign n1321 =  ( n1320 ) == ( bv_8_110_n504 )  ;
assign n1322 = in[15:8] ;
assign n1323 =  ( n1322 ) == ( bv_8_109_n289 )  ;
assign n1324 = in[15:8] ;
assign n1325 =  ( n1324 ) == ( bv_8_108_n272 )  ;
assign n1326 = in[15:8] ;
assign n1327 =  ( n1326 ) == ( bv_8_107_n513 )  ;
assign n1328 = in[15:8] ;
assign n1329 =  ( n1328 ) == ( bv_8_106_n516 )  ;
assign n1330 = in[15:8] ;
assign n1331 =  ( n1330 ) == ( bv_8_105_n113 )  ;
assign n1332 = in[15:8] ;
assign n1333 =  ( n1332 ) == ( bv_8_104_n39 )  ;
assign n1334 = in[15:8] ;
assign n1335 =  ( n1334 ) == ( bv_8_103_n525 )  ;
assign n1336 = in[15:8] ;
assign n1337 =  ( n1336 ) == ( bv_8_102_n176 )  ;
assign n1338 = in[15:8] ;
assign n1339 =  ( n1338 ) == ( bv_8_101_n261 )  ;
assign n1340 = in[15:8] ;
assign n1341 =  ( n1340 ) == ( bv_8_100_n417 )  ;
assign n1342 = in[15:8] ;
assign n1343 =  ( n1342 ) == ( bv_8_99_n537 )  ;
assign n1344 = in[15:8] ;
assign n1345 =  ( n1344 ) == ( bv_8_98_n316 )  ;
assign n1346 = in[15:8] ;
assign n1347 =  ( n1346 ) == ( bv_8_97_n157 )  ;
assign n1348 = in[15:8] ;
assign n1349 =  ( n1348 ) == ( bv_8_96_n404 )  ;
assign n1350 = in[15:8] ;
assign n1351 =  ( n1350 ) == ( bv_8_95_n440 )  ;
assign n1352 = in[15:8] ;
assign n1353 =  ( n1352 ) == ( bv_8_94_n363 )  ;
assign n1354 = in[15:8] ;
assign n1355 =  ( n1354 ) == ( bv_8_93_n414 )  ;
assign n1356 = in[15:8] ;
assign n1357 =  ( n1356 ) == ( bv_8_92_n328 )  ;
assign n1358 = in[15:8] ;
assign n1359 =  ( n1358 ) == ( bv_8_91_n557 )  ;
assign n1360 = in[15:8] ;
assign n1361 =  ( n1360 ) == ( bv_8_90_n561 )  ;
assign n1362 = in[15:8] ;
assign n1363 =  ( n1362 ) == ( bv_8_89_n564 )  ;
assign n1364 = in[15:8] ;
assign n1365 =  ( n1364 ) == ( bv_8_88_n549 )  ;
assign n1366 = in[15:8] ;
assign n1367 =  ( n1366 ) == ( bv_8_87_n150 )  ;
assign n1368 = in[15:8] ;
assign n1369 =  ( n1368 ) == ( bv_8_86_n268 )  ;
assign n1370 = in[15:8] ;
assign n1371 =  ( n1370 ) == ( bv_8_85_n79 )  ;
assign n1372 = in[15:8] ;
assign n1373 =  ( n1372 ) == ( bv_8_84_n15 )  ;
assign n1374 = in[15:8] ;
assign n1375 =  ( n1374 ) == ( bv_8_83_n578 )  ;
assign n1376 = in[15:8] ;
assign n1377 =  ( n1376 ) == ( bv_8_82_n581 )  ;
assign n1378 = in[15:8] ;
assign n1379 =  ( n1378 ) == ( bv_8_81_n499 )  ;
assign n1380 = in[15:8] ;
assign n1381 =  ( n1380 ) == ( bv_8_80_n511 )  ;
assign n1382 = in[15:8] ;
assign n1383 =  ( n1382 ) == ( bv_8_79_n398 )  ;
assign n1384 = in[15:8] ;
assign n1385 =  ( n1384 ) == ( bv_8_78_n280 )  ;
assign n1386 = in[15:8] ;
assign n1387 =  ( n1386 ) == ( bv_8_77_n532 )  ;
assign n1388 = in[15:8] ;
assign n1389 =  ( n1388 ) == ( bv_8_76_n552 )  ;
assign n1390 = in[15:8] ;
assign n1391 =  ( n1390 ) == ( bv_8_75_n203 )  ;
assign n1392 = in[15:8] ;
assign n1393 =  ( n1392 ) == ( bv_8_74_n555 )  ;
assign n1394 = in[15:8] ;
assign n1395 =  ( n1394 ) == ( bv_8_73_n339 )  ;
assign n1396 = in[15:8] ;
assign n1397 =  ( n1396 ) == ( bv_8_72_n172 )  ;
assign n1398 = in[15:8] ;
assign n1399 =  ( n1398 ) == ( bv_8_71_n608 )  ;
assign n1400 = in[15:8] ;
assign n1401 =  ( n1400 ) == ( bv_8_70_n377 )  ;
assign n1402 = in[15:8] ;
assign n1403 =  ( n1402 ) == ( bv_8_69_n523 )  ;
assign n1404 = in[15:8] ;
assign n1405 =  ( n1404 ) == ( bv_8_68_n433 )  ;
assign n1406 = in[15:8] ;
assign n1407 =  ( n1406 ) == ( bv_8_67_n535 )  ;
assign n1408 = in[15:8] ;
assign n1409 =  ( n1408 ) == ( bv_8_66_n43 )  ;
assign n1410 = in[15:8] ;
assign n1411 =  ( n1410 ) == ( bv_8_65_n35 )  ;
assign n1412 = in[15:8] ;
assign n1413 =  ( n1412 ) == ( bv_8_64_n493 )  ;
assign n1414 = in[15:8] ;
assign n1415 =  ( n1414 ) == ( bv_8_63_n629 )  ;
assign n1416 = in[15:8] ;
assign n1417 =  ( n1416 ) == ( bv_8_62_n184 )  ;
assign n1418 = in[15:8] ;
assign n1419 =  ( n1418 ) == ( bv_8_61_n420 )  ;
assign n1420 = in[15:8] ;
assign n1421 =  ( n1420 ) == ( bv_8_60_n508 )  ;
assign n1422 = in[15:8] ;
assign n1423 =  ( n1422 ) == ( bv_8_59_n604 )  ;
assign n1424 = in[15:8] ;
assign n1425 =  ( n1424 ) == ( bv_8_58_n347 )  ;
assign n1426 = in[15:8] ;
assign n1427 =  ( n1426 ) == ( bv_8_57_n559 )  ;
assign n1428 = in[15:8] ;
assign n1429 =  ( n1428 ) == ( bv_8_56_n482 )  ;
assign n1430 = in[15:8] ;
assign n1431 =  ( n1430 ) == ( bv_8_55_n293 )  ;
assign n1432 = in[15:8] ;
assign n1433 =  ( n1432 ) == ( bv_8_54_n651 )  ;
assign n1434 = in[15:8] ;
assign n1435 =  ( n1434 ) == ( bv_8_53_n153 )  ;
assign n1436 = in[15:8] ;
assign n1437 =  ( n1436 ) == ( bv_8_52_n657 )  ;
assign n1438 = in[15:8] ;
assign n1439 =  ( n1438 ) == ( bv_8_51_n529 )  ;
assign n1440 = in[15:8] ;
assign n1441 =  ( n1440 ) == ( bv_8_50_n350 )  ;
assign n1442 = in[15:8] ;
assign n1443 =  ( n1442 ) == ( bv_8_49_n666 )  ;
assign n1444 = in[15:8] ;
assign n1445 =  ( n1444 ) == ( bv_8_48_n669 )  ;
assign n1446 = in[15:8] ;
assign n1447 =  ( n1446 ) == ( bv_8_47_n592 )  ;
assign n1448 = in[15:8] ;
assign n1449 =  ( n1448 ) == ( bv_8_46_n236 )  ;
assign n1450 = in[15:8] ;
assign n1451 =  ( n1450 ) == ( bv_8_45_n27 )  ;
assign n1452 = in[15:8] ;
assign n1453 =  ( n1452 ) == ( bv_8_44_n622 )  ;
assign n1454 = in[15:8] ;
assign n1455 =  ( n1454 ) == ( bv_8_43_n682 )  ;
assign n1456 = in[15:8] ;
assign n1457 =  ( n1456 ) == ( bv_8_42_n388 )  ;
assign n1458 = in[15:8] ;
assign n1459 =  ( n1458 ) == ( bv_8_41_n597 )  ;
assign n1460 = in[15:8] ;
assign n1461 =  ( n1460 ) == ( bv_8_40_n75 )  ;
assign n1462 = in[15:8] ;
assign n1463 =  ( n1462 ) == ( bv_8_39_n635 )  ;
assign n1464 = in[15:8] ;
assign n1465 =  ( n1464 ) == ( bv_8_38_n693 )  ;
assign n1466 = in[15:8] ;
assign n1467 =  ( n1466 ) == ( bv_8_37_n240 )  ;
assign n1468 = in[15:8] ;
assign n1469 =  ( n1468 ) == ( bv_8_36_n331 )  ;
assign n1470 = in[15:8] ;
assign n1471 =  ( n1470 ) == ( bv_8_35_n664 )  ;
assign n1472 = in[15:8] ;
assign n1473 =  ( n1472 ) == ( bv_8_34_n391 )  ;
assign n1474 = in[15:8] ;
assign n1475 =  ( n1474 ) == ( bv_8_33_n469 )  ;
assign n1476 = in[15:8] ;
assign n1477 =  ( n1476 ) == ( bv_8_32_n576 )  ;
assign n1478 = in[15:8] ;
assign n1479 =  ( n1478 ) == ( bv_8_31_n207 )  ;
assign n1480 = in[15:8] ;
assign n1481 =  ( n1480 ) == ( bv_8_30_n94 )  ;
assign n1482 = in[15:8] ;
assign n1483 =  ( n1482 ) == ( bv_8_29_n134 )  ;
assign n1484 = in[15:8] ;
assign n1485 =  ( n1484 ) == ( bv_8_28_n232 )  ;
assign n1486 = in[15:8] ;
assign n1487 =  ( n1486 ) == ( bv_8_27_n616 )  ;
assign n1488 = in[15:8] ;
assign n1489 =  ( n1488 ) == ( bv_8_26_n619 )  ;
assign n1490 = in[15:8] ;
assign n1491 =  ( n1490 ) == ( bv_8_25_n411 )  ;
assign n1492 = in[15:8] ;
assign n1493 =  ( n1492 ) == ( bv_8_24_n659 )  ;
assign n1494 = in[15:8] ;
assign n1495 =  ( n1494 ) == ( bv_8_23_n430 )  ;
assign n1496 = in[15:8] ;
assign n1497 =  ( n1496 ) == ( bv_8_22_n7 )  ;
assign n1498 = in[15:8] ;
assign n1499 =  ( n1498 ) == ( bv_8_21_n674 )  ;
assign n1500 = in[15:8] ;
assign n1501 =  ( n1500 ) == ( bv_8_20_n369 )  ;
assign n1502 = in[15:8] ;
assign n1503 =  ( n1502 ) == ( bv_8_19_n447 )  ;
assign n1504 = in[15:8] ;
assign n1505 =  ( n1504 ) == ( bv_8_18_n644 )  ;
assign n1506 = in[15:8] ;
assign n1507 =  ( n1506 ) == ( bv_8_17_n117 )  ;
assign n1508 = in[15:8] ;
assign n1509 =  ( n1508 ) == ( bv_8_16_n465 )  ;
assign n1510 = in[15:8] ;
assign n1511 =  ( n1510 ) == ( bv_8_15_n23 )  ;
assign n1512 = in[15:8] ;
assign n1513 =  ( n1512 ) == ( bv_8_14_n161 )  ;
assign n1514 = in[15:8] ;
assign n1515 =  ( n1514 ) == ( bv_8_13_n55 )  ;
assign n1516 = in[15:8] ;
assign n1517 =  ( n1516 ) == ( bv_8_12_n450 )  ;
assign n1518 = in[15:8] ;
assign n1519 =  ( n1518 ) == ( bv_8_11_n359 )  ;
assign n1520 = in[15:8] ;
assign n1521 =  ( n1520 ) == ( bv_8_10_n343 )  ;
assign n1522 = in[15:8] ;
assign n1523 =  ( n1522 ) == ( bv_8_9_n627 )  ;
assign n1524 = in[15:8] ;
assign n1525 =  ( n1524 ) == ( bv_8_8_n250 )  ;
assign n1526 = in[15:8] ;
assign n1527 =  ( n1526 ) == ( bv_8_7_n647 )  ;
assign n1528 = in[15:8] ;
assign n1529 =  ( n1528 ) == ( bv_8_6_n335 )  ;
assign n1530 = in[15:8] ;
assign n1531 =  ( n1530 ) == ( bv_8_5_n653 )  ;
assign n1532 = in[15:8] ;
assign n1533 =  ( n1532 ) == ( bv_8_4_n671 )  ;
assign n1534 = in[15:8] ;
assign n1535 =  ( n1534 ) == ( bv_8_3_n168 )  ;
assign n1536 = in[15:8] ;
assign n1537 =  ( n1536 ) == ( bv_8_2_n518 )  ;
assign n1538 = in[15:8] ;
assign n1539 =  ( n1538 ) == ( bv_8_1_n753 )  ;
assign n1540 = in[15:8] ;
assign n1541 =  ( n1540 ) == ( bv_8_0_n583 )  ;
assign n1542 =  ( n1541 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n1543 =  ( n1539 ) ? ( bv_8_124_n463 ) : ( n1542 ) ;
assign n1544 =  ( n1537 ) ? ( bv_8_119_n477 ) : ( n1543 ) ;
assign n1545 =  ( n1535 ) ? ( bv_8_123_n467 ) : ( n1544 ) ;
assign n1546 =  ( n1533 ) ? ( bv_8_242_n57 ) : ( n1545 ) ;
assign n1547 =  ( n1531 ) ? ( bv_8_107_n513 ) : ( n1546 ) ;
assign n1548 =  ( n1529 ) ? ( bv_8_111_n501 ) : ( n1547 ) ;
assign n1549 =  ( n1527 ) ? ( bv_8_197_n226 ) : ( n1548 ) ;
assign n1550 =  ( n1525 ) ? ( bv_8_48_n669 ) : ( n1549 ) ;
assign n1551 =  ( n1523 ) ? ( bv_8_1_n753 ) : ( n1550 ) ;
assign n1552 =  ( n1521 ) ? ( bv_8_103_n525 ) : ( n1551 ) ;
assign n1553 =  ( n1519 ) ? ( bv_8_43_n682 ) : ( n1552 ) ;
assign n1554 =  ( n1517 ) ? ( bv_8_254_n9 ) : ( n1553 ) ;
assign n1555 =  ( n1515 ) ? ( bv_8_215_n159 ) : ( n1554 ) ;
assign n1556 =  ( n1513 ) ? ( bv_8_171_n314 ) : ( n1555 ) ;
assign n1557 =  ( n1511 ) ? ( bv_8_118_n480 ) : ( n1556 ) ;
assign n1558 =  ( n1509 ) ? ( bv_8_202_n209 ) : ( n1557 ) ;
assign n1559 =  ( n1507 ) ? ( bv_8_130_n445 ) : ( n1558 ) ;
assign n1560 =  ( n1505 ) ? ( bv_8_201_n213 ) : ( n1559 ) ;
assign n1561 =  ( n1503 ) ? ( bv_8_125_n460 ) : ( n1560 ) ;
assign n1562 =  ( n1501 ) ? ( bv_8_250_n25 ) : ( n1561 ) ;
assign n1563 =  ( n1499 ) ? ( bv_8_89_n564 ) : ( n1562 ) ;
assign n1564 =  ( n1497 ) ? ( bv_8_71_n608 ) : ( n1563 ) ;
assign n1565 =  ( n1495 ) ? ( bv_8_240_n65 ) : ( n1564 ) ;
assign n1566 =  ( n1493 ) ? ( bv_8_173_n306 ) : ( n1565 ) ;
assign n1567 =  ( n1491 ) ? ( bv_8_212_n170 ) : ( n1566 ) ;
assign n1568 =  ( n1489 ) ? ( bv_8_162_n345 ) : ( n1567 ) ;
assign n1569 =  ( n1487 ) ? ( bv_8_175_n300 ) : ( n1568 ) ;
assign n1570 =  ( n1485 ) ? ( bv_8_156_n365 ) : ( n1569 ) ;
assign n1571 =  ( n1483 ) ? ( bv_8_164_n337 ) : ( n1570 ) ;
assign n1572 =  ( n1481 ) ? ( bv_8_114_n491 ) : ( n1571 ) ;
assign n1573 =  ( n1479 ) ? ( bv_8_192_n245 ) : ( n1572 ) ;
assign n1574 =  ( n1477 ) ? ( bv_8_183_n274 ) : ( n1573 ) ;
assign n1575 =  ( n1475 ) ? ( bv_8_253_n13 ) : ( n1574 ) ;
assign n1576 =  ( n1473 ) ? ( bv_8_147_n393 ) : ( n1575 ) ;
assign n1577 =  ( n1471 ) ? ( bv_8_38_n693 ) : ( n1576 ) ;
assign n1578 =  ( n1469 ) ? ( bv_8_54_n651 ) : ( n1577 ) ;
assign n1579 =  ( n1467 ) ? ( bv_8_63_n629 ) : ( n1578 ) ;
assign n1580 =  ( n1465 ) ? ( bv_8_247_n37 ) : ( n1579 ) ;
assign n1581 =  ( n1463 ) ? ( bv_8_204_n201 ) : ( n1580 ) ;
assign n1582 =  ( n1461 ) ? ( bv_8_52_n657 ) : ( n1581 ) ;
assign n1583 =  ( n1459 ) ? ( bv_8_165_n333 ) : ( n1582 ) ;
assign n1584 =  ( n1457 ) ? ( bv_8_229_n107 ) : ( n1583 ) ;
assign n1585 =  ( n1455 ) ? ( bv_8_241_n61 ) : ( n1584 ) ;
assign n1586 =  ( n1453 ) ? ( bv_8_113_n495 ) : ( n1585 ) ;
assign n1587 =  ( n1451 ) ? ( bv_8_216_n155 ) : ( n1586 ) ;
assign n1588 =  ( n1449 ) ? ( bv_8_49_n666 ) : ( n1587 ) ;
assign n1589 =  ( n1447 ) ? ( bv_8_21_n674 ) : ( n1588 ) ;
assign n1590 =  ( n1445 ) ? ( bv_8_4_n671 ) : ( n1589 ) ;
assign n1591 =  ( n1443 ) ? ( bv_8_199_n219 ) : ( n1590 ) ;
assign n1592 =  ( n1441 ) ? ( bv_8_35_n664 ) : ( n1591 ) ;
assign n1593 =  ( n1439 ) ? ( bv_8_195_n234 ) : ( n1592 ) ;
assign n1594 =  ( n1437 ) ? ( bv_8_24_n659 ) : ( n1593 ) ;
assign n1595 =  ( n1435 ) ? ( bv_8_150_n383 ) : ( n1594 ) ;
assign n1596 =  ( n1433 ) ? ( bv_8_5_n653 ) : ( n1595 ) ;
assign n1597 =  ( n1431 ) ? ( bv_8_154_n371 ) : ( n1596 ) ;
assign n1598 =  ( n1429 ) ? ( bv_8_7_n647 ) : ( n1597 ) ;
assign n1599 =  ( n1427 ) ? ( bv_8_18_n644 ) : ( n1598 ) ;
assign n1600 =  ( n1425 ) ? ( bv_8_128_n452 ) : ( n1599 ) ;
assign n1601 =  ( n1423 ) ? ( bv_8_226_n119 ) : ( n1600 ) ;
assign n1602 =  ( n1421 ) ? ( bv_8_235_n85 ) : ( n1601 ) ;
assign n1603 =  ( n1419 ) ? ( bv_8_39_n635 ) : ( n1602 ) ;
assign n1604 =  ( n1417 ) ? ( bv_8_178_n291 ) : ( n1603 ) ;
assign n1605 =  ( n1415 ) ? ( bv_8_117_n484 ) : ( n1604 ) ;
assign n1606 =  ( n1413 ) ? ( bv_8_9_n627 ) : ( n1605 ) ;
assign n1607 =  ( n1411 ) ? ( bv_8_131_n442 ) : ( n1606 ) ;
assign n1608 =  ( n1409 ) ? ( bv_8_44_n622 ) : ( n1607 ) ;
assign n1609 =  ( n1407 ) ? ( bv_8_26_n619 ) : ( n1608 ) ;
assign n1610 =  ( n1405 ) ? ( bv_8_27_n616 ) : ( n1609 ) ;
assign n1611 =  ( n1403 ) ? ( bv_8_110_n504 ) : ( n1610 ) ;
assign n1612 =  ( n1401 ) ? ( bv_8_90_n561 ) : ( n1611 ) ;
assign n1613 =  ( n1399 ) ? ( bv_8_160_n352 ) : ( n1612 ) ;
assign n1614 =  ( n1397 ) ? ( bv_8_82_n581 ) : ( n1613 ) ;
assign n1615 =  ( n1395 ) ? ( bv_8_59_n604 ) : ( n1614 ) ;
assign n1616 =  ( n1393 ) ? ( bv_8_214_n163 ) : ( n1615 ) ;
assign n1617 =  ( n1391 ) ? ( bv_8_179_n287 ) : ( n1616 ) ;
assign n1618 =  ( n1389 ) ? ( bv_8_41_n597 ) : ( n1617 ) ;
assign n1619 =  ( n1387 ) ? ( bv_8_227_n115 ) : ( n1618 ) ;
assign n1620 =  ( n1385 ) ? ( bv_8_47_n592 ) : ( n1619 ) ;
assign n1621 =  ( n1383 ) ? ( bv_8_132_n438 ) : ( n1620 ) ;
assign n1622 =  ( n1381 ) ? ( bv_8_83_n578 ) : ( n1621 ) ;
assign n1623 =  ( n1379 ) ? ( bv_8_209_n182 ) : ( n1622 ) ;
assign n1624 =  ( n1377 ) ? ( bv_8_0_n583 ) : ( n1623 ) ;
assign n1625 =  ( n1375 ) ? ( bv_8_237_n77 ) : ( n1624 ) ;
assign n1626 =  ( n1373 ) ? ( bv_8_32_n576 ) : ( n1625 ) ;
assign n1627 =  ( n1371 ) ? ( bv_8_252_n17 ) : ( n1626 ) ;
assign n1628 =  ( n1369 ) ? ( bv_8_177_n295 ) : ( n1627 ) ;
assign n1629 =  ( n1367 ) ? ( bv_8_91_n557 ) : ( n1628 ) ;
assign n1630 =  ( n1365 ) ? ( bv_8_106_n516 ) : ( n1629 ) ;
assign n1631 =  ( n1363 ) ? ( bv_8_203_n205 ) : ( n1630 ) ;
assign n1632 =  ( n1361 ) ? ( bv_8_190_n252 ) : ( n1631 ) ;
assign n1633 =  ( n1359 ) ? ( bv_8_57_n559 ) : ( n1632 ) ;
assign n1634 =  ( n1357 ) ? ( bv_8_74_n555 ) : ( n1633 ) ;
assign n1635 =  ( n1355 ) ? ( bv_8_76_n552 ) : ( n1634 ) ;
assign n1636 =  ( n1353 ) ? ( bv_8_88_n549 ) : ( n1635 ) ;
assign n1637 =  ( n1351 ) ? ( bv_8_207_n190 ) : ( n1636 ) ;
assign n1638 =  ( n1349 ) ? ( bv_8_208_n186 ) : ( n1637 ) ;
assign n1639 =  ( n1347 ) ? ( bv_8_239_n69 ) : ( n1638 ) ;
assign n1640 =  ( n1345 ) ? ( bv_8_170_n318 ) : ( n1639 ) ;
assign n1641 =  ( n1343 ) ? ( bv_8_251_n21 ) : ( n1640 ) ;
assign n1642 =  ( n1341 ) ? ( bv_8_67_n535 ) : ( n1641 ) ;
assign n1643 =  ( n1339 ) ? ( bv_8_77_n532 ) : ( n1642 ) ;
assign n1644 =  ( n1337 ) ? ( bv_8_51_n529 ) : ( n1643 ) ;
assign n1645 =  ( n1335 ) ? ( bv_8_133_n435 ) : ( n1644 ) ;
assign n1646 =  ( n1333 ) ? ( bv_8_69_n523 ) : ( n1645 ) ;
assign n1647 =  ( n1331 ) ? ( bv_8_249_n29 ) : ( n1646 ) ;
assign n1648 =  ( n1329 ) ? ( bv_8_2_n518 ) : ( n1647 ) ;
assign n1649 =  ( n1327 ) ? ( bv_8_127_n455 ) : ( n1648 ) ;
assign n1650 =  ( n1325 ) ? ( bv_8_80_n511 ) : ( n1649 ) ;
assign n1651 =  ( n1323 ) ? ( bv_8_60_n508 ) : ( n1650 ) ;
assign n1652 =  ( n1321 ) ? ( bv_8_159_n355 ) : ( n1651 ) ;
assign n1653 =  ( n1319 ) ? ( bv_8_168_n323 ) : ( n1652 ) ;
assign n1654 =  ( n1317 ) ? ( bv_8_81_n499 ) : ( n1653 ) ;
assign n1655 =  ( n1315 ) ? ( bv_8_163_n341 ) : ( n1654 ) ;
assign n1656 =  ( n1313 ) ? ( bv_8_64_n493 ) : ( n1655 ) ;
assign n1657 =  ( n1311 ) ? ( bv_8_143_n406 ) : ( n1656 ) ;
assign n1658 =  ( n1309 ) ? ( bv_8_146_n396 ) : ( n1657 ) ;
assign n1659 =  ( n1307 ) ? ( bv_8_157_n361 ) : ( n1658 ) ;
assign n1660 =  ( n1305 ) ? ( bv_8_56_n482 ) : ( n1659 ) ;
assign n1661 =  ( n1303 ) ? ( bv_8_245_n45 ) : ( n1660 ) ;
assign n1662 =  ( n1301 ) ? ( bv_8_188_n259 ) : ( n1661 ) ;
assign n1663 =  ( n1299 ) ? ( bv_8_182_n278 ) : ( n1662 ) ;
assign n1664 =  ( n1297 ) ? ( bv_8_218_n148 ) : ( n1663 ) ;
assign n1665 =  ( n1295 ) ? ( bv_8_33_n469 ) : ( n1664 ) ;
assign n1666 =  ( n1293 ) ? ( bv_8_16_n465 ) : ( n1665 ) ;
assign n1667 =  ( n1291 ) ? ( bv_8_255_n5 ) : ( n1666 ) ;
assign n1668 =  ( n1289 ) ? ( bv_8_243_n53 ) : ( n1667 ) ;
assign n1669 =  ( n1287 ) ? ( bv_8_210_n178 ) : ( n1668 ) ;
assign n1670 =  ( n1285 ) ? ( bv_8_205_n197 ) : ( n1669 ) ;
assign n1671 =  ( n1283 ) ? ( bv_8_12_n450 ) : ( n1670 ) ;
assign n1672 =  ( n1281 ) ? ( bv_8_19_n447 ) : ( n1671 ) ;
assign n1673 =  ( n1279 ) ? ( bv_8_236_n81 ) : ( n1672 ) ;
assign n1674 =  ( n1277 ) ? ( bv_8_95_n440 ) : ( n1673 ) ;
assign n1675 =  ( n1275 ) ? ( bv_8_151_n379 ) : ( n1674 ) ;
assign n1676 =  ( n1273 ) ? ( bv_8_68_n433 ) : ( n1675 ) ;
assign n1677 =  ( n1271 ) ? ( bv_8_23_n430 ) : ( n1676 ) ;
assign n1678 =  ( n1269 ) ? ( bv_8_196_n230 ) : ( n1677 ) ;
assign n1679 =  ( n1267 ) ? ( bv_8_167_n326 ) : ( n1678 ) ;
assign n1680 =  ( n1265 ) ? ( bv_8_126_n423 ) : ( n1679 ) ;
assign n1681 =  ( n1263 ) ? ( bv_8_61_n420 ) : ( n1680 ) ;
assign n1682 =  ( n1261 ) ? ( bv_8_100_n417 ) : ( n1681 ) ;
assign n1683 =  ( n1259 ) ? ( bv_8_93_n414 ) : ( n1682 ) ;
assign n1684 =  ( n1257 ) ? ( bv_8_25_n411 ) : ( n1683 ) ;
assign n1685 =  ( n1255 ) ? ( bv_8_115_n408 ) : ( n1684 ) ;
assign n1686 =  ( n1253 ) ? ( bv_8_96_n404 ) : ( n1685 ) ;
assign n1687 =  ( n1251 ) ? ( bv_8_129_n401 ) : ( n1686 ) ;
assign n1688 =  ( n1249 ) ? ( bv_8_79_n398 ) : ( n1687 ) ;
assign n1689 =  ( n1247 ) ? ( bv_8_220_n140 ) : ( n1688 ) ;
assign n1690 =  ( n1245 ) ? ( bv_8_34_n391 ) : ( n1689 ) ;
assign n1691 =  ( n1243 ) ? ( bv_8_42_n388 ) : ( n1690 ) ;
assign n1692 =  ( n1241 ) ? ( bv_8_144_n385 ) : ( n1691 ) ;
assign n1693 =  ( n1239 ) ? ( bv_8_136_n381 ) : ( n1692 ) ;
assign n1694 =  ( n1237 ) ? ( bv_8_70_n377 ) : ( n1693 ) ;
assign n1695 =  ( n1235 ) ? ( bv_8_238_n73 ) : ( n1694 ) ;
assign n1696 =  ( n1233 ) ? ( bv_8_184_n270 ) : ( n1695 ) ;
assign n1697 =  ( n1231 ) ? ( bv_8_20_n369 ) : ( n1696 ) ;
assign n1698 =  ( n1229 ) ? ( bv_8_222_n132 ) : ( n1697 ) ;
assign n1699 =  ( n1227 ) ? ( bv_8_94_n363 ) : ( n1698 ) ;
assign n1700 =  ( n1225 ) ? ( bv_8_11_n359 ) : ( n1699 ) ;
assign n1701 =  ( n1223 ) ? ( bv_8_219_n144 ) : ( n1700 ) ;
assign n1702 =  ( n1221 ) ? ( bv_8_224_n126 ) : ( n1701 ) ;
assign n1703 =  ( n1219 ) ? ( bv_8_50_n350 ) : ( n1702 ) ;
assign n1704 =  ( n1217 ) ? ( bv_8_58_n347 ) : ( n1703 ) ;
assign n1705 =  ( n1215 ) ? ( bv_8_10_n343 ) : ( n1704 ) ;
assign n1706 =  ( n1213 ) ? ( bv_8_73_n339 ) : ( n1705 ) ;
assign n1707 =  ( n1211 ) ? ( bv_8_6_n335 ) : ( n1706 ) ;
assign n1708 =  ( n1209 ) ? ( bv_8_36_n331 ) : ( n1707 ) ;
assign n1709 =  ( n1207 ) ? ( bv_8_92_n328 ) : ( n1708 ) ;
assign n1710 =  ( n1205 ) ? ( bv_8_194_n238 ) : ( n1709 ) ;
assign n1711 =  ( n1203 ) ? ( bv_8_211_n174 ) : ( n1710 ) ;
assign n1712 =  ( n1201 ) ? ( bv_8_172_n310 ) : ( n1711 ) ;
assign n1713 =  ( n1199 ) ? ( bv_8_98_n316 ) : ( n1712 ) ;
assign n1714 =  ( n1197 ) ? ( bv_8_145_n312 ) : ( n1713 ) ;
assign n1715 =  ( n1195 ) ? ( bv_8_149_n308 ) : ( n1714 ) ;
assign n1716 =  ( n1193 ) ? ( bv_8_228_n111 ) : ( n1715 ) ;
assign n1717 =  ( n1191 ) ? ( bv_8_121_n302 ) : ( n1716 ) ;
assign n1718 =  ( n1189 ) ? ( bv_8_231_n100 ) : ( n1717 ) ;
assign n1719 =  ( n1187 ) ? ( bv_8_200_n216 ) : ( n1718 ) ;
assign n1720 =  ( n1185 ) ? ( bv_8_55_n293 ) : ( n1719 ) ;
assign n1721 =  ( n1183 ) ? ( bv_8_109_n289 ) : ( n1720 ) ;
assign n1722 =  ( n1181 ) ? ( bv_8_141_n285 ) : ( n1721 ) ;
assign n1723 =  ( n1179 ) ? ( bv_8_213_n166 ) : ( n1722 ) ;
assign n1724 =  ( n1177 ) ? ( bv_8_78_n280 ) : ( n1723 ) ;
assign n1725 =  ( n1175 ) ? ( bv_8_169_n276 ) : ( n1724 ) ;
assign n1726 =  ( n1173 ) ? ( bv_8_108_n272 ) : ( n1725 ) ;
assign n1727 =  ( n1171 ) ? ( bv_8_86_n268 ) : ( n1726 ) ;
assign n1728 =  ( n1169 ) ? ( bv_8_244_n49 ) : ( n1727 ) ;
assign n1729 =  ( n1167 ) ? ( bv_8_234_n89 ) : ( n1728 ) ;
assign n1730 =  ( n1165 ) ? ( bv_8_101_n261 ) : ( n1729 ) ;
assign n1731 =  ( n1163 ) ? ( bv_8_122_n257 ) : ( n1730 ) ;
assign n1732 =  ( n1161 ) ? ( bv_8_174_n254 ) : ( n1731 ) ;
assign n1733 =  ( n1159 ) ? ( bv_8_8_n250 ) : ( n1732 ) ;
assign n1734 =  ( n1157 ) ? ( bv_8_186_n247 ) : ( n1733 ) ;
assign n1735 =  ( n1155 ) ? ( bv_8_120_n243 ) : ( n1734 ) ;
assign n1736 =  ( n1153 ) ? ( bv_8_37_n240 ) : ( n1735 ) ;
assign n1737 =  ( n1151 ) ? ( bv_8_46_n236 ) : ( n1736 ) ;
assign n1738 =  ( n1149 ) ? ( bv_8_28_n232 ) : ( n1737 ) ;
assign n1739 =  ( n1147 ) ? ( bv_8_166_n228 ) : ( n1738 ) ;
assign n1740 =  ( n1145 ) ? ( bv_8_180_n224 ) : ( n1739 ) ;
assign n1741 =  ( n1143 ) ? ( bv_8_198_n221 ) : ( n1740 ) ;
assign n1742 =  ( n1141 ) ? ( bv_8_232_n96 ) : ( n1741 ) ;
assign n1743 =  ( n1139 ) ? ( bv_8_221_n136 ) : ( n1742 ) ;
assign n1744 =  ( n1137 ) ? ( bv_8_116_n211 ) : ( n1743 ) ;
assign n1745 =  ( n1135 ) ? ( bv_8_31_n207 ) : ( n1744 ) ;
assign n1746 =  ( n1133 ) ? ( bv_8_75_n203 ) : ( n1745 ) ;
assign n1747 =  ( n1131 ) ? ( bv_8_189_n199 ) : ( n1746 ) ;
assign n1748 =  ( n1129 ) ? ( bv_8_139_n195 ) : ( n1747 ) ;
assign n1749 =  ( n1127 ) ? ( bv_8_138_n192 ) : ( n1748 ) ;
assign n1750 =  ( n1125 ) ? ( bv_8_112_n188 ) : ( n1749 ) ;
assign n1751 =  ( n1123 ) ? ( bv_8_62_n184 ) : ( n1750 ) ;
assign n1752 =  ( n1121 ) ? ( bv_8_181_n180 ) : ( n1751 ) ;
assign n1753 =  ( n1119 ) ? ( bv_8_102_n176 ) : ( n1752 ) ;
assign n1754 =  ( n1117 ) ? ( bv_8_72_n172 ) : ( n1753 ) ;
assign n1755 =  ( n1115 ) ? ( bv_8_3_n168 ) : ( n1754 ) ;
assign n1756 =  ( n1113 ) ? ( bv_8_246_n41 ) : ( n1755 ) ;
assign n1757 =  ( n1111 ) ? ( bv_8_14_n161 ) : ( n1756 ) ;
assign n1758 =  ( n1109 ) ? ( bv_8_97_n157 ) : ( n1757 ) ;
assign n1759 =  ( n1107 ) ? ( bv_8_53_n153 ) : ( n1758 ) ;
assign n1760 =  ( n1105 ) ? ( bv_8_87_n150 ) : ( n1759 ) ;
assign n1761 =  ( n1103 ) ? ( bv_8_185_n146 ) : ( n1760 ) ;
assign n1762 =  ( n1101 ) ? ( bv_8_134_n142 ) : ( n1761 ) ;
assign n1763 =  ( n1099 ) ? ( bv_8_193_n138 ) : ( n1762 ) ;
assign n1764 =  ( n1097 ) ? ( bv_8_29_n134 ) : ( n1763 ) ;
assign n1765 =  ( n1095 ) ? ( bv_8_158_n130 ) : ( n1764 ) ;
assign n1766 =  ( n1093 ) ? ( bv_8_225_n123 ) : ( n1765 ) ;
assign n1767 =  ( n1091 ) ? ( bv_8_248_n33 ) : ( n1766 ) ;
assign n1768 =  ( n1089 ) ? ( bv_8_152_n121 ) : ( n1767 ) ;
assign n1769 =  ( n1087 ) ? ( bv_8_17_n117 ) : ( n1768 ) ;
assign n1770 =  ( n1085 ) ? ( bv_8_105_n113 ) : ( n1769 ) ;
assign n1771 =  ( n1083 ) ? ( bv_8_217_n109 ) : ( n1770 ) ;
assign n1772 =  ( n1081 ) ? ( bv_8_142_n105 ) : ( n1771 ) ;
assign n1773 =  ( n1079 ) ? ( bv_8_148_n102 ) : ( n1772 ) ;
assign n1774 =  ( n1077 ) ? ( bv_8_155_n98 ) : ( n1773 ) ;
assign n1775 =  ( n1075 ) ? ( bv_8_30_n94 ) : ( n1774 ) ;
assign n1776 =  ( n1073 ) ? ( bv_8_135_n91 ) : ( n1775 ) ;
assign n1777 =  ( n1071 ) ? ( bv_8_233_n87 ) : ( n1776 ) ;
assign n1778 =  ( n1069 ) ? ( bv_8_206_n83 ) : ( n1777 ) ;
assign n1779 =  ( n1067 ) ? ( bv_8_85_n79 ) : ( n1778 ) ;
assign n1780 =  ( n1065 ) ? ( bv_8_40_n75 ) : ( n1779 ) ;
assign n1781 =  ( n1063 ) ? ( bv_8_223_n71 ) : ( n1780 ) ;
assign n1782 =  ( n1061 ) ? ( bv_8_140_n67 ) : ( n1781 ) ;
assign n1783 =  ( n1059 ) ? ( bv_8_161_n63 ) : ( n1782 ) ;
assign n1784 =  ( n1057 ) ? ( bv_8_137_n59 ) : ( n1783 ) ;
assign n1785 =  ( n1055 ) ? ( bv_8_13_n55 ) : ( n1784 ) ;
assign n1786 =  ( n1053 ) ? ( bv_8_191_n51 ) : ( n1785 ) ;
assign n1787 =  ( n1051 ) ? ( bv_8_230_n47 ) : ( n1786 ) ;
assign n1788 =  ( n1049 ) ? ( bv_8_66_n43 ) : ( n1787 ) ;
assign n1789 =  ( n1047 ) ? ( bv_8_104_n39 ) : ( n1788 ) ;
assign n1790 =  ( n1045 ) ? ( bv_8_65_n35 ) : ( n1789 ) ;
assign n1791 =  ( n1043 ) ? ( bv_8_153_n31 ) : ( n1790 ) ;
assign n1792 =  ( n1041 ) ? ( bv_8_45_n27 ) : ( n1791 ) ;
assign n1793 =  ( n1039 ) ? ( bv_8_15_n23 ) : ( n1792 ) ;
assign n1794 =  ( n1037 ) ? ( bv_8_176_n19 ) : ( n1793 ) ;
assign n1795 =  ( n1035 ) ? ( bv_8_84_n15 ) : ( n1794 ) ;
assign n1796 =  ( n1033 ) ? ( bv_8_187_n11 ) : ( n1795 ) ;
assign n1797 =  ( n1031 ) ? ( bv_8_22_n7 ) : ( n1796 ) ;
assign n1798 =  ( n1029 ) ^ ( n1797 )  ;
assign n1799 =  { ( n1028 ) , ( n1798 ) }  ;
assign n1800 = in[111:104] ;
assign n1801 = in[7:0] ;
assign n1802 =  ( n1801 ) == ( bv_8_255_n5 )  ;
assign n1803 = in[7:0] ;
assign n1804 =  ( n1803 ) == ( bv_8_254_n9 )  ;
assign n1805 = in[7:0] ;
assign n1806 =  ( n1805 ) == ( bv_8_253_n13 )  ;
assign n1807 = in[7:0] ;
assign n1808 =  ( n1807 ) == ( bv_8_252_n17 )  ;
assign n1809 = in[7:0] ;
assign n1810 =  ( n1809 ) == ( bv_8_251_n21 )  ;
assign n1811 = in[7:0] ;
assign n1812 =  ( n1811 ) == ( bv_8_250_n25 )  ;
assign n1813 = in[7:0] ;
assign n1814 =  ( n1813 ) == ( bv_8_249_n29 )  ;
assign n1815 = in[7:0] ;
assign n1816 =  ( n1815 ) == ( bv_8_248_n33 )  ;
assign n1817 = in[7:0] ;
assign n1818 =  ( n1817 ) == ( bv_8_247_n37 )  ;
assign n1819 = in[7:0] ;
assign n1820 =  ( n1819 ) == ( bv_8_246_n41 )  ;
assign n1821 = in[7:0] ;
assign n1822 =  ( n1821 ) == ( bv_8_245_n45 )  ;
assign n1823 = in[7:0] ;
assign n1824 =  ( n1823 ) == ( bv_8_244_n49 )  ;
assign n1825 = in[7:0] ;
assign n1826 =  ( n1825 ) == ( bv_8_243_n53 )  ;
assign n1827 = in[7:0] ;
assign n1828 =  ( n1827 ) == ( bv_8_242_n57 )  ;
assign n1829 = in[7:0] ;
assign n1830 =  ( n1829 ) == ( bv_8_241_n61 )  ;
assign n1831 = in[7:0] ;
assign n1832 =  ( n1831 ) == ( bv_8_240_n65 )  ;
assign n1833 = in[7:0] ;
assign n1834 =  ( n1833 ) == ( bv_8_239_n69 )  ;
assign n1835 = in[7:0] ;
assign n1836 =  ( n1835 ) == ( bv_8_238_n73 )  ;
assign n1837 = in[7:0] ;
assign n1838 =  ( n1837 ) == ( bv_8_237_n77 )  ;
assign n1839 = in[7:0] ;
assign n1840 =  ( n1839 ) == ( bv_8_236_n81 )  ;
assign n1841 = in[7:0] ;
assign n1842 =  ( n1841 ) == ( bv_8_235_n85 )  ;
assign n1843 = in[7:0] ;
assign n1844 =  ( n1843 ) == ( bv_8_234_n89 )  ;
assign n1845 = in[7:0] ;
assign n1846 =  ( n1845 ) == ( bv_8_233_n87 )  ;
assign n1847 = in[7:0] ;
assign n1848 =  ( n1847 ) == ( bv_8_232_n96 )  ;
assign n1849 = in[7:0] ;
assign n1850 =  ( n1849 ) == ( bv_8_231_n100 )  ;
assign n1851 = in[7:0] ;
assign n1852 =  ( n1851 ) == ( bv_8_230_n47 )  ;
assign n1853 = in[7:0] ;
assign n1854 =  ( n1853 ) == ( bv_8_229_n107 )  ;
assign n1855 = in[7:0] ;
assign n1856 =  ( n1855 ) == ( bv_8_228_n111 )  ;
assign n1857 = in[7:0] ;
assign n1858 =  ( n1857 ) == ( bv_8_227_n115 )  ;
assign n1859 = in[7:0] ;
assign n1860 =  ( n1859 ) == ( bv_8_226_n119 )  ;
assign n1861 = in[7:0] ;
assign n1862 =  ( n1861 ) == ( bv_8_225_n123 )  ;
assign n1863 = in[7:0] ;
assign n1864 =  ( n1863 ) == ( bv_8_224_n126 )  ;
assign n1865 = in[7:0] ;
assign n1866 =  ( n1865 ) == ( bv_8_223_n71 )  ;
assign n1867 = in[7:0] ;
assign n1868 =  ( n1867 ) == ( bv_8_222_n132 )  ;
assign n1869 = in[7:0] ;
assign n1870 =  ( n1869 ) == ( bv_8_221_n136 )  ;
assign n1871 = in[7:0] ;
assign n1872 =  ( n1871 ) == ( bv_8_220_n140 )  ;
assign n1873 = in[7:0] ;
assign n1874 =  ( n1873 ) == ( bv_8_219_n144 )  ;
assign n1875 = in[7:0] ;
assign n1876 =  ( n1875 ) == ( bv_8_218_n148 )  ;
assign n1877 = in[7:0] ;
assign n1878 =  ( n1877 ) == ( bv_8_217_n109 )  ;
assign n1879 = in[7:0] ;
assign n1880 =  ( n1879 ) == ( bv_8_216_n155 )  ;
assign n1881 = in[7:0] ;
assign n1882 =  ( n1881 ) == ( bv_8_215_n159 )  ;
assign n1883 = in[7:0] ;
assign n1884 =  ( n1883 ) == ( bv_8_214_n163 )  ;
assign n1885 = in[7:0] ;
assign n1886 =  ( n1885 ) == ( bv_8_213_n166 )  ;
assign n1887 = in[7:0] ;
assign n1888 =  ( n1887 ) == ( bv_8_212_n170 )  ;
assign n1889 = in[7:0] ;
assign n1890 =  ( n1889 ) == ( bv_8_211_n174 )  ;
assign n1891 = in[7:0] ;
assign n1892 =  ( n1891 ) == ( bv_8_210_n178 )  ;
assign n1893 = in[7:0] ;
assign n1894 =  ( n1893 ) == ( bv_8_209_n182 )  ;
assign n1895 = in[7:0] ;
assign n1896 =  ( n1895 ) == ( bv_8_208_n186 )  ;
assign n1897 = in[7:0] ;
assign n1898 =  ( n1897 ) == ( bv_8_207_n190 )  ;
assign n1899 = in[7:0] ;
assign n1900 =  ( n1899 ) == ( bv_8_206_n83 )  ;
assign n1901 = in[7:0] ;
assign n1902 =  ( n1901 ) == ( bv_8_205_n197 )  ;
assign n1903 = in[7:0] ;
assign n1904 =  ( n1903 ) == ( bv_8_204_n201 )  ;
assign n1905 = in[7:0] ;
assign n1906 =  ( n1905 ) == ( bv_8_203_n205 )  ;
assign n1907 = in[7:0] ;
assign n1908 =  ( n1907 ) == ( bv_8_202_n209 )  ;
assign n1909 = in[7:0] ;
assign n1910 =  ( n1909 ) == ( bv_8_201_n213 )  ;
assign n1911 = in[7:0] ;
assign n1912 =  ( n1911 ) == ( bv_8_200_n216 )  ;
assign n1913 = in[7:0] ;
assign n1914 =  ( n1913 ) == ( bv_8_199_n219 )  ;
assign n1915 = in[7:0] ;
assign n1916 =  ( n1915 ) == ( bv_8_198_n221 )  ;
assign n1917 = in[7:0] ;
assign n1918 =  ( n1917 ) == ( bv_8_197_n226 )  ;
assign n1919 = in[7:0] ;
assign n1920 =  ( n1919 ) == ( bv_8_196_n230 )  ;
assign n1921 = in[7:0] ;
assign n1922 =  ( n1921 ) == ( bv_8_195_n234 )  ;
assign n1923 = in[7:0] ;
assign n1924 =  ( n1923 ) == ( bv_8_194_n238 )  ;
assign n1925 = in[7:0] ;
assign n1926 =  ( n1925 ) == ( bv_8_193_n138 )  ;
assign n1927 = in[7:0] ;
assign n1928 =  ( n1927 ) == ( bv_8_192_n245 )  ;
assign n1929 = in[7:0] ;
assign n1930 =  ( n1929 ) == ( bv_8_191_n51 )  ;
assign n1931 = in[7:0] ;
assign n1932 =  ( n1931 ) == ( bv_8_190_n252 )  ;
assign n1933 = in[7:0] ;
assign n1934 =  ( n1933 ) == ( bv_8_189_n199 )  ;
assign n1935 = in[7:0] ;
assign n1936 =  ( n1935 ) == ( bv_8_188_n259 )  ;
assign n1937 = in[7:0] ;
assign n1938 =  ( n1937 ) == ( bv_8_187_n11 )  ;
assign n1939 = in[7:0] ;
assign n1940 =  ( n1939 ) == ( bv_8_186_n247 )  ;
assign n1941 = in[7:0] ;
assign n1942 =  ( n1941 ) == ( bv_8_185_n146 )  ;
assign n1943 = in[7:0] ;
assign n1944 =  ( n1943 ) == ( bv_8_184_n270 )  ;
assign n1945 = in[7:0] ;
assign n1946 =  ( n1945 ) == ( bv_8_183_n274 )  ;
assign n1947 = in[7:0] ;
assign n1948 =  ( n1947 ) == ( bv_8_182_n278 )  ;
assign n1949 = in[7:0] ;
assign n1950 =  ( n1949 ) == ( bv_8_181_n180 )  ;
assign n1951 = in[7:0] ;
assign n1952 =  ( n1951 ) == ( bv_8_180_n224 )  ;
assign n1953 = in[7:0] ;
assign n1954 =  ( n1953 ) == ( bv_8_179_n287 )  ;
assign n1955 = in[7:0] ;
assign n1956 =  ( n1955 ) == ( bv_8_178_n291 )  ;
assign n1957 = in[7:0] ;
assign n1958 =  ( n1957 ) == ( bv_8_177_n295 )  ;
assign n1959 = in[7:0] ;
assign n1960 =  ( n1959 ) == ( bv_8_176_n19 )  ;
assign n1961 = in[7:0] ;
assign n1962 =  ( n1961 ) == ( bv_8_175_n300 )  ;
assign n1963 = in[7:0] ;
assign n1964 =  ( n1963 ) == ( bv_8_174_n254 )  ;
assign n1965 = in[7:0] ;
assign n1966 =  ( n1965 ) == ( bv_8_173_n306 )  ;
assign n1967 = in[7:0] ;
assign n1968 =  ( n1967 ) == ( bv_8_172_n310 )  ;
assign n1969 = in[7:0] ;
assign n1970 =  ( n1969 ) == ( bv_8_171_n314 )  ;
assign n1971 = in[7:0] ;
assign n1972 =  ( n1971 ) == ( bv_8_170_n318 )  ;
assign n1973 = in[7:0] ;
assign n1974 =  ( n1973 ) == ( bv_8_169_n276 )  ;
assign n1975 = in[7:0] ;
assign n1976 =  ( n1975 ) == ( bv_8_168_n323 )  ;
assign n1977 = in[7:0] ;
assign n1978 =  ( n1977 ) == ( bv_8_167_n326 )  ;
assign n1979 = in[7:0] ;
assign n1980 =  ( n1979 ) == ( bv_8_166_n228 )  ;
assign n1981 = in[7:0] ;
assign n1982 =  ( n1981 ) == ( bv_8_165_n333 )  ;
assign n1983 = in[7:0] ;
assign n1984 =  ( n1983 ) == ( bv_8_164_n337 )  ;
assign n1985 = in[7:0] ;
assign n1986 =  ( n1985 ) == ( bv_8_163_n341 )  ;
assign n1987 = in[7:0] ;
assign n1988 =  ( n1987 ) == ( bv_8_162_n345 )  ;
assign n1989 = in[7:0] ;
assign n1990 =  ( n1989 ) == ( bv_8_161_n63 )  ;
assign n1991 = in[7:0] ;
assign n1992 =  ( n1991 ) == ( bv_8_160_n352 )  ;
assign n1993 = in[7:0] ;
assign n1994 =  ( n1993 ) == ( bv_8_159_n355 )  ;
assign n1995 = in[7:0] ;
assign n1996 =  ( n1995 ) == ( bv_8_158_n130 )  ;
assign n1997 = in[7:0] ;
assign n1998 =  ( n1997 ) == ( bv_8_157_n361 )  ;
assign n1999 = in[7:0] ;
assign n2000 =  ( n1999 ) == ( bv_8_156_n365 )  ;
assign n2001 = in[7:0] ;
assign n2002 =  ( n2001 ) == ( bv_8_155_n98 )  ;
assign n2003 = in[7:0] ;
assign n2004 =  ( n2003 ) == ( bv_8_154_n371 )  ;
assign n2005 = in[7:0] ;
assign n2006 =  ( n2005 ) == ( bv_8_153_n31 )  ;
assign n2007 = in[7:0] ;
assign n2008 =  ( n2007 ) == ( bv_8_152_n121 )  ;
assign n2009 = in[7:0] ;
assign n2010 =  ( n2009 ) == ( bv_8_151_n379 )  ;
assign n2011 = in[7:0] ;
assign n2012 =  ( n2011 ) == ( bv_8_150_n383 )  ;
assign n2013 = in[7:0] ;
assign n2014 =  ( n2013 ) == ( bv_8_149_n308 )  ;
assign n2015 = in[7:0] ;
assign n2016 =  ( n2015 ) == ( bv_8_148_n102 )  ;
assign n2017 = in[7:0] ;
assign n2018 =  ( n2017 ) == ( bv_8_147_n393 )  ;
assign n2019 = in[7:0] ;
assign n2020 =  ( n2019 ) == ( bv_8_146_n396 )  ;
assign n2021 = in[7:0] ;
assign n2022 =  ( n2021 ) == ( bv_8_145_n312 )  ;
assign n2023 = in[7:0] ;
assign n2024 =  ( n2023 ) == ( bv_8_144_n385 )  ;
assign n2025 = in[7:0] ;
assign n2026 =  ( n2025 ) == ( bv_8_143_n406 )  ;
assign n2027 = in[7:0] ;
assign n2028 =  ( n2027 ) == ( bv_8_142_n105 )  ;
assign n2029 = in[7:0] ;
assign n2030 =  ( n2029 ) == ( bv_8_141_n285 )  ;
assign n2031 = in[7:0] ;
assign n2032 =  ( n2031 ) == ( bv_8_140_n67 )  ;
assign n2033 = in[7:0] ;
assign n2034 =  ( n2033 ) == ( bv_8_139_n195 )  ;
assign n2035 = in[7:0] ;
assign n2036 =  ( n2035 ) == ( bv_8_138_n192 )  ;
assign n2037 = in[7:0] ;
assign n2038 =  ( n2037 ) == ( bv_8_137_n59 )  ;
assign n2039 = in[7:0] ;
assign n2040 =  ( n2039 ) == ( bv_8_136_n381 )  ;
assign n2041 = in[7:0] ;
assign n2042 =  ( n2041 ) == ( bv_8_135_n91 )  ;
assign n2043 = in[7:0] ;
assign n2044 =  ( n2043 ) == ( bv_8_134_n142 )  ;
assign n2045 = in[7:0] ;
assign n2046 =  ( n2045 ) == ( bv_8_133_n435 )  ;
assign n2047 = in[7:0] ;
assign n2048 =  ( n2047 ) == ( bv_8_132_n438 )  ;
assign n2049 = in[7:0] ;
assign n2050 =  ( n2049 ) == ( bv_8_131_n442 )  ;
assign n2051 = in[7:0] ;
assign n2052 =  ( n2051 ) == ( bv_8_130_n445 )  ;
assign n2053 = in[7:0] ;
assign n2054 =  ( n2053 ) == ( bv_8_129_n401 )  ;
assign n2055 = in[7:0] ;
assign n2056 =  ( n2055 ) == ( bv_8_128_n452 )  ;
assign n2057 = in[7:0] ;
assign n2058 =  ( n2057 ) == ( bv_8_127_n455 )  ;
assign n2059 = in[7:0] ;
assign n2060 =  ( n2059 ) == ( bv_8_126_n423 )  ;
assign n2061 = in[7:0] ;
assign n2062 =  ( n2061 ) == ( bv_8_125_n460 )  ;
assign n2063 = in[7:0] ;
assign n2064 =  ( n2063 ) == ( bv_8_124_n463 )  ;
assign n2065 = in[7:0] ;
assign n2066 =  ( n2065 ) == ( bv_8_123_n467 )  ;
assign n2067 = in[7:0] ;
assign n2068 =  ( n2067 ) == ( bv_8_122_n257 )  ;
assign n2069 = in[7:0] ;
assign n2070 =  ( n2069 ) == ( bv_8_121_n302 )  ;
assign n2071 = in[7:0] ;
assign n2072 =  ( n2071 ) == ( bv_8_120_n243 )  ;
assign n2073 = in[7:0] ;
assign n2074 =  ( n2073 ) == ( bv_8_119_n477 )  ;
assign n2075 = in[7:0] ;
assign n2076 =  ( n2075 ) == ( bv_8_118_n480 )  ;
assign n2077 = in[7:0] ;
assign n2078 =  ( n2077 ) == ( bv_8_117_n484 )  ;
assign n2079 = in[7:0] ;
assign n2080 =  ( n2079 ) == ( bv_8_116_n211 )  ;
assign n2081 = in[7:0] ;
assign n2082 =  ( n2081 ) == ( bv_8_115_n408 )  ;
assign n2083 = in[7:0] ;
assign n2084 =  ( n2083 ) == ( bv_8_114_n491 )  ;
assign n2085 = in[7:0] ;
assign n2086 =  ( n2085 ) == ( bv_8_113_n495 )  ;
assign n2087 = in[7:0] ;
assign n2088 =  ( n2087 ) == ( bv_8_112_n188 )  ;
assign n2089 = in[7:0] ;
assign n2090 =  ( n2089 ) == ( bv_8_111_n501 )  ;
assign n2091 = in[7:0] ;
assign n2092 =  ( n2091 ) == ( bv_8_110_n504 )  ;
assign n2093 = in[7:0] ;
assign n2094 =  ( n2093 ) == ( bv_8_109_n289 )  ;
assign n2095 = in[7:0] ;
assign n2096 =  ( n2095 ) == ( bv_8_108_n272 )  ;
assign n2097 = in[7:0] ;
assign n2098 =  ( n2097 ) == ( bv_8_107_n513 )  ;
assign n2099 = in[7:0] ;
assign n2100 =  ( n2099 ) == ( bv_8_106_n516 )  ;
assign n2101 = in[7:0] ;
assign n2102 =  ( n2101 ) == ( bv_8_105_n113 )  ;
assign n2103 = in[7:0] ;
assign n2104 =  ( n2103 ) == ( bv_8_104_n39 )  ;
assign n2105 = in[7:0] ;
assign n2106 =  ( n2105 ) == ( bv_8_103_n525 )  ;
assign n2107 = in[7:0] ;
assign n2108 =  ( n2107 ) == ( bv_8_102_n176 )  ;
assign n2109 = in[7:0] ;
assign n2110 =  ( n2109 ) == ( bv_8_101_n261 )  ;
assign n2111 = in[7:0] ;
assign n2112 =  ( n2111 ) == ( bv_8_100_n417 )  ;
assign n2113 = in[7:0] ;
assign n2114 =  ( n2113 ) == ( bv_8_99_n537 )  ;
assign n2115 = in[7:0] ;
assign n2116 =  ( n2115 ) == ( bv_8_98_n316 )  ;
assign n2117 = in[7:0] ;
assign n2118 =  ( n2117 ) == ( bv_8_97_n157 )  ;
assign n2119 = in[7:0] ;
assign n2120 =  ( n2119 ) == ( bv_8_96_n404 )  ;
assign n2121 = in[7:0] ;
assign n2122 =  ( n2121 ) == ( bv_8_95_n440 )  ;
assign n2123 = in[7:0] ;
assign n2124 =  ( n2123 ) == ( bv_8_94_n363 )  ;
assign n2125 = in[7:0] ;
assign n2126 =  ( n2125 ) == ( bv_8_93_n414 )  ;
assign n2127 = in[7:0] ;
assign n2128 =  ( n2127 ) == ( bv_8_92_n328 )  ;
assign n2129 = in[7:0] ;
assign n2130 =  ( n2129 ) == ( bv_8_91_n557 )  ;
assign n2131 = in[7:0] ;
assign n2132 =  ( n2131 ) == ( bv_8_90_n561 )  ;
assign n2133 = in[7:0] ;
assign n2134 =  ( n2133 ) == ( bv_8_89_n564 )  ;
assign n2135 = in[7:0] ;
assign n2136 =  ( n2135 ) == ( bv_8_88_n549 )  ;
assign n2137 = in[7:0] ;
assign n2138 =  ( n2137 ) == ( bv_8_87_n150 )  ;
assign n2139 = in[7:0] ;
assign n2140 =  ( n2139 ) == ( bv_8_86_n268 )  ;
assign n2141 = in[7:0] ;
assign n2142 =  ( n2141 ) == ( bv_8_85_n79 )  ;
assign n2143 = in[7:0] ;
assign n2144 =  ( n2143 ) == ( bv_8_84_n15 )  ;
assign n2145 = in[7:0] ;
assign n2146 =  ( n2145 ) == ( bv_8_83_n578 )  ;
assign n2147 = in[7:0] ;
assign n2148 =  ( n2147 ) == ( bv_8_82_n581 )  ;
assign n2149 = in[7:0] ;
assign n2150 =  ( n2149 ) == ( bv_8_81_n499 )  ;
assign n2151 = in[7:0] ;
assign n2152 =  ( n2151 ) == ( bv_8_80_n511 )  ;
assign n2153 = in[7:0] ;
assign n2154 =  ( n2153 ) == ( bv_8_79_n398 )  ;
assign n2155 = in[7:0] ;
assign n2156 =  ( n2155 ) == ( bv_8_78_n280 )  ;
assign n2157 = in[7:0] ;
assign n2158 =  ( n2157 ) == ( bv_8_77_n532 )  ;
assign n2159 = in[7:0] ;
assign n2160 =  ( n2159 ) == ( bv_8_76_n552 )  ;
assign n2161 = in[7:0] ;
assign n2162 =  ( n2161 ) == ( bv_8_75_n203 )  ;
assign n2163 = in[7:0] ;
assign n2164 =  ( n2163 ) == ( bv_8_74_n555 )  ;
assign n2165 = in[7:0] ;
assign n2166 =  ( n2165 ) == ( bv_8_73_n339 )  ;
assign n2167 = in[7:0] ;
assign n2168 =  ( n2167 ) == ( bv_8_72_n172 )  ;
assign n2169 = in[7:0] ;
assign n2170 =  ( n2169 ) == ( bv_8_71_n608 )  ;
assign n2171 = in[7:0] ;
assign n2172 =  ( n2171 ) == ( bv_8_70_n377 )  ;
assign n2173 = in[7:0] ;
assign n2174 =  ( n2173 ) == ( bv_8_69_n523 )  ;
assign n2175 = in[7:0] ;
assign n2176 =  ( n2175 ) == ( bv_8_68_n433 )  ;
assign n2177 = in[7:0] ;
assign n2178 =  ( n2177 ) == ( bv_8_67_n535 )  ;
assign n2179 = in[7:0] ;
assign n2180 =  ( n2179 ) == ( bv_8_66_n43 )  ;
assign n2181 = in[7:0] ;
assign n2182 =  ( n2181 ) == ( bv_8_65_n35 )  ;
assign n2183 = in[7:0] ;
assign n2184 =  ( n2183 ) == ( bv_8_64_n493 )  ;
assign n2185 = in[7:0] ;
assign n2186 =  ( n2185 ) == ( bv_8_63_n629 )  ;
assign n2187 = in[7:0] ;
assign n2188 =  ( n2187 ) == ( bv_8_62_n184 )  ;
assign n2189 = in[7:0] ;
assign n2190 =  ( n2189 ) == ( bv_8_61_n420 )  ;
assign n2191 = in[7:0] ;
assign n2192 =  ( n2191 ) == ( bv_8_60_n508 )  ;
assign n2193 = in[7:0] ;
assign n2194 =  ( n2193 ) == ( bv_8_59_n604 )  ;
assign n2195 = in[7:0] ;
assign n2196 =  ( n2195 ) == ( bv_8_58_n347 )  ;
assign n2197 = in[7:0] ;
assign n2198 =  ( n2197 ) == ( bv_8_57_n559 )  ;
assign n2199 = in[7:0] ;
assign n2200 =  ( n2199 ) == ( bv_8_56_n482 )  ;
assign n2201 = in[7:0] ;
assign n2202 =  ( n2201 ) == ( bv_8_55_n293 )  ;
assign n2203 = in[7:0] ;
assign n2204 =  ( n2203 ) == ( bv_8_54_n651 )  ;
assign n2205 = in[7:0] ;
assign n2206 =  ( n2205 ) == ( bv_8_53_n153 )  ;
assign n2207 = in[7:0] ;
assign n2208 =  ( n2207 ) == ( bv_8_52_n657 )  ;
assign n2209 = in[7:0] ;
assign n2210 =  ( n2209 ) == ( bv_8_51_n529 )  ;
assign n2211 = in[7:0] ;
assign n2212 =  ( n2211 ) == ( bv_8_50_n350 )  ;
assign n2213 = in[7:0] ;
assign n2214 =  ( n2213 ) == ( bv_8_49_n666 )  ;
assign n2215 = in[7:0] ;
assign n2216 =  ( n2215 ) == ( bv_8_48_n669 )  ;
assign n2217 = in[7:0] ;
assign n2218 =  ( n2217 ) == ( bv_8_47_n592 )  ;
assign n2219 = in[7:0] ;
assign n2220 =  ( n2219 ) == ( bv_8_46_n236 )  ;
assign n2221 = in[7:0] ;
assign n2222 =  ( n2221 ) == ( bv_8_45_n27 )  ;
assign n2223 = in[7:0] ;
assign n2224 =  ( n2223 ) == ( bv_8_44_n622 )  ;
assign n2225 = in[7:0] ;
assign n2226 =  ( n2225 ) == ( bv_8_43_n682 )  ;
assign n2227 = in[7:0] ;
assign n2228 =  ( n2227 ) == ( bv_8_42_n388 )  ;
assign n2229 = in[7:0] ;
assign n2230 =  ( n2229 ) == ( bv_8_41_n597 )  ;
assign n2231 = in[7:0] ;
assign n2232 =  ( n2231 ) == ( bv_8_40_n75 )  ;
assign n2233 = in[7:0] ;
assign n2234 =  ( n2233 ) == ( bv_8_39_n635 )  ;
assign n2235 = in[7:0] ;
assign n2236 =  ( n2235 ) == ( bv_8_38_n693 )  ;
assign n2237 = in[7:0] ;
assign n2238 =  ( n2237 ) == ( bv_8_37_n240 )  ;
assign n2239 = in[7:0] ;
assign n2240 =  ( n2239 ) == ( bv_8_36_n331 )  ;
assign n2241 = in[7:0] ;
assign n2242 =  ( n2241 ) == ( bv_8_35_n664 )  ;
assign n2243 = in[7:0] ;
assign n2244 =  ( n2243 ) == ( bv_8_34_n391 )  ;
assign n2245 = in[7:0] ;
assign n2246 =  ( n2245 ) == ( bv_8_33_n469 )  ;
assign n2247 = in[7:0] ;
assign n2248 =  ( n2247 ) == ( bv_8_32_n576 )  ;
assign n2249 = in[7:0] ;
assign n2250 =  ( n2249 ) == ( bv_8_31_n207 )  ;
assign n2251 = in[7:0] ;
assign n2252 =  ( n2251 ) == ( bv_8_30_n94 )  ;
assign n2253 = in[7:0] ;
assign n2254 =  ( n2253 ) == ( bv_8_29_n134 )  ;
assign n2255 = in[7:0] ;
assign n2256 =  ( n2255 ) == ( bv_8_28_n232 )  ;
assign n2257 = in[7:0] ;
assign n2258 =  ( n2257 ) == ( bv_8_27_n616 )  ;
assign n2259 = in[7:0] ;
assign n2260 =  ( n2259 ) == ( bv_8_26_n619 )  ;
assign n2261 = in[7:0] ;
assign n2262 =  ( n2261 ) == ( bv_8_25_n411 )  ;
assign n2263 = in[7:0] ;
assign n2264 =  ( n2263 ) == ( bv_8_24_n659 )  ;
assign n2265 = in[7:0] ;
assign n2266 =  ( n2265 ) == ( bv_8_23_n430 )  ;
assign n2267 = in[7:0] ;
assign n2268 =  ( n2267 ) == ( bv_8_22_n7 )  ;
assign n2269 = in[7:0] ;
assign n2270 =  ( n2269 ) == ( bv_8_21_n674 )  ;
assign n2271 = in[7:0] ;
assign n2272 =  ( n2271 ) == ( bv_8_20_n369 )  ;
assign n2273 = in[7:0] ;
assign n2274 =  ( n2273 ) == ( bv_8_19_n447 )  ;
assign n2275 = in[7:0] ;
assign n2276 =  ( n2275 ) == ( bv_8_18_n644 )  ;
assign n2277 = in[7:0] ;
assign n2278 =  ( n2277 ) == ( bv_8_17_n117 )  ;
assign n2279 = in[7:0] ;
assign n2280 =  ( n2279 ) == ( bv_8_16_n465 )  ;
assign n2281 = in[7:0] ;
assign n2282 =  ( n2281 ) == ( bv_8_15_n23 )  ;
assign n2283 = in[7:0] ;
assign n2284 =  ( n2283 ) == ( bv_8_14_n161 )  ;
assign n2285 = in[7:0] ;
assign n2286 =  ( n2285 ) == ( bv_8_13_n55 )  ;
assign n2287 = in[7:0] ;
assign n2288 =  ( n2287 ) == ( bv_8_12_n450 )  ;
assign n2289 = in[7:0] ;
assign n2290 =  ( n2289 ) == ( bv_8_11_n359 )  ;
assign n2291 = in[7:0] ;
assign n2292 =  ( n2291 ) == ( bv_8_10_n343 )  ;
assign n2293 = in[7:0] ;
assign n2294 =  ( n2293 ) == ( bv_8_9_n627 )  ;
assign n2295 = in[7:0] ;
assign n2296 =  ( n2295 ) == ( bv_8_8_n250 )  ;
assign n2297 = in[7:0] ;
assign n2298 =  ( n2297 ) == ( bv_8_7_n647 )  ;
assign n2299 = in[7:0] ;
assign n2300 =  ( n2299 ) == ( bv_8_6_n335 )  ;
assign n2301 = in[7:0] ;
assign n2302 =  ( n2301 ) == ( bv_8_5_n653 )  ;
assign n2303 = in[7:0] ;
assign n2304 =  ( n2303 ) == ( bv_8_4_n671 )  ;
assign n2305 = in[7:0] ;
assign n2306 =  ( n2305 ) == ( bv_8_3_n168 )  ;
assign n2307 = in[7:0] ;
assign n2308 =  ( n2307 ) == ( bv_8_2_n518 )  ;
assign n2309 = in[7:0] ;
assign n2310 =  ( n2309 ) == ( bv_8_1_n753 )  ;
assign n2311 = in[7:0] ;
assign n2312 =  ( n2311 ) == ( bv_8_0_n583 )  ;
assign n2313 =  ( n2312 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n2314 =  ( n2310 ) ? ( bv_8_124_n463 ) : ( n2313 ) ;
assign n2315 =  ( n2308 ) ? ( bv_8_119_n477 ) : ( n2314 ) ;
assign n2316 =  ( n2306 ) ? ( bv_8_123_n467 ) : ( n2315 ) ;
assign n2317 =  ( n2304 ) ? ( bv_8_242_n57 ) : ( n2316 ) ;
assign n2318 =  ( n2302 ) ? ( bv_8_107_n513 ) : ( n2317 ) ;
assign n2319 =  ( n2300 ) ? ( bv_8_111_n501 ) : ( n2318 ) ;
assign n2320 =  ( n2298 ) ? ( bv_8_197_n226 ) : ( n2319 ) ;
assign n2321 =  ( n2296 ) ? ( bv_8_48_n669 ) : ( n2320 ) ;
assign n2322 =  ( n2294 ) ? ( bv_8_1_n753 ) : ( n2321 ) ;
assign n2323 =  ( n2292 ) ? ( bv_8_103_n525 ) : ( n2322 ) ;
assign n2324 =  ( n2290 ) ? ( bv_8_43_n682 ) : ( n2323 ) ;
assign n2325 =  ( n2288 ) ? ( bv_8_254_n9 ) : ( n2324 ) ;
assign n2326 =  ( n2286 ) ? ( bv_8_215_n159 ) : ( n2325 ) ;
assign n2327 =  ( n2284 ) ? ( bv_8_171_n314 ) : ( n2326 ) ;
assign n2328 =  ( n2282 ) ? ( bv_8_118_n480 ) : ( n2327 ) ;
assign n2329 =  ( n2280 ) ? ( bv_8_202_n209 ) : ( n2328 ) ;
assign n2330 =  ( n2278 ) ? ( bv_8_130_n445 ) : ( n2329 ) ;
assign n2331 =  ( n2276 ) ? ( bv_8_201_n213 ) : ( n2330 ) ;
assign n2332 =  ( n2274 ) ? ( bv_8_125_n460 ) : ( n2331 ) ;
assign n2333 =  ( n2272 ) ? ( bv_8_250_n25 ) : ( n2332 ) ;
assign n2334 =  ( n2270 ) ? ( bv_8_89_n564 ) : ( n2333 ) ;
assign n2335 =  ( n2268 ) ? ( bv_8_71_n608 ) : ( n2334 ) ;
assign n2336 =  ( n2266 ) ? ( bv_8_240_n65 ) : ( n2335 ) ;
assign n2337 =  ( n2264 ) ? ( bv_8_173_n306 ) : ( n2336 ) ;
assign n2338 =  ( n2262 ) ? ( bv_8_212_n170 ) : ( n2337 ) ;
assign n2339 =  ( n2260 ) ? ( bv_8_162_n345 ) : ( n2338 ) ;
assign n2340 =  ( n2258 ) ? ( bv_8_175_n300 ) : ( n2339 ) ;
assign n2341 =  ( n2256 ) ? ( bv_8_156_n365 ) : ( n2340 ) ;
assign n2342 =  ( n2254 ) ? ( bv_8_164_n337 ) : ( n2341 ) ;
assign n2343 =  ( n2252 ) ? ( bv_8_114_n491 ) : ( n2342 ) ;
assign n2344 =  ( n2250 ) ? ( bv_8_192_n245 ) : ( n2343 ) ;
assign n2345 =  ( n2248 ) ? ( bv_8_183_n274 ) : ( n2344 ) ;
assign n2346 =  ( n2246 ) ? ( bv_8_253_n13 ) : ( n2345 ) ;
assign n2347 =  ( n2244 ) ? ( bv_8_147_n393 ) : ( n2346 ) ;
assign n2348 =  ( n2242 ) ? ( bv_8_38_n693 ) : ( n2347 ) ;
assign n2349 =  ( n2240 ) ? ( bv_8_54_n651 ) : ( n2348 ) ;
assign n2350 =  ( n2238 ) ? ( bv_8_63_n629 ) : ( n2349 ) ;
assign n2351 =  ( n2236 ) ? ( bv_8_247_n37 ) : ( n2350 ) ;
assign n2352 =  ( n2234 ) ? ( bv_8_204_n201 ) : ( n2351 ) ;
assign n2353 =  ( n2232 ) ? ( bv_8_52_n657 ) : ( n2352 ) ;
assign n2354 =  ( n2230 ) ? ( bv_8_165_n333 ) : ( n2353 ) ;
assign n2355 =  ( n2228 ) ? ( bv_8_229_n107 ) : ( n2354 ) ;
assign n2356 =  ( n2226 ) ? ( bv_8_241_n61 ) : ( n2355 ) ;
assign n2357 =  ( n2224 ) ? ( bv_8_113_n495 ) : ( n2356 ) ;
assign n2358 =  ( n2222 ) ? ( bv_8_216_n155 ) : ( n2357 ) ;
assign n2359 =  ( n2220 ) ? ( bv_8_49_n666 ) : ( n2358 ) ;
assign n2360 =  ( n2218 ) ? ( bv_8_21_n674 ) : ( n2359 ) ;
assign n2361 =  ( n2216 ) ? ( bv_8_4_n671 ) : ( n2360 ) ;
assign n2362 =  ( n2214 ) ? ( bv_8_199_n219 ) : ( n2361 ) ;
assign n2363 =  ( n2212 ) ? ( bv_8_35_n664 ) : ( n2362 ) ;
assign n2364 =  ( n2210 ) ? ( bv_8_195_n234 ) : ( n2363 ) ;
assign n2365 =  ( n2208 ) ? ( bv_8_24_n659 ) : ( n2364 ) ;
assign n2366 =  ( n2206 ) ? ( bv_8_150_n383 ) : ( n2365 ) ;
assign n2367 =  ( n2204 ) ? ( bv_8_5_n653 ) : ( n2366 ) ;
assign n2368 =  ( n2202 ) ? ( bv_8_154_n371 ) : ( n2367 ) ;
assign n2369 =  ( n2200 ) ? ( bv_8_7_n647 ) : ( n2368 ) ;
assign n2370 =  ( n2198 ) ? ( bv_8_18_n644 ) : ( n2369 ) ;
assign n2371 =  ( n2196 ) ? ( bv_8_128_n452 ) : ( n2370 ) ;
assign n2372 =  ( n2194 ) ? ( bv_8_226_n119 ) : ( n2371 ) ;
assign n2373 =  ( n2192 ) ? ( bv_8_235_n85 ) : ( n2372 ) ;
assign n2374 =  ( n2190 ) ? ( bv_8_39_n635 ) : ( n2373 ) ;
assign n2375 =  ( n2188 ) ? ( bv_8_178_n291 ) : ( n2374 ) ;
assign n2376 =  ( n2186 ) ? ( bv_8_117_n484 ) : ( n2375 ) ;
assign n2377 =  ( n2184 ) ? ( bv_8_9_n627 ) : ( n2376 ) ;
assign n2378 =  ( n2182 ) ? ( bv_8_131_n442 ) : ( n2377 ) ;
assign n2379 =  ( n2180 ) ? ( bv_8_44_n622 ) : ( n2378 ) ;
assign n2380 =  ( n2178 ) ? ( bv_8_26_n619 ) : ( n2379 ) ;
assign n2381 =  ( n2176 ) ? ( bv_8_27_n616 ) : ( n2380 ) ;
assign n2382 =  ( n2174 ) ? ( bv_8_110_n504 ) : ( n2381 ) ;
assign n2383 =  ( n2172 ) ? ( bv_8_90_n561 ) : ( n2382 ) ;
assign n2384 =  ( n2170 ) ? ( bv_8_160_n352 ) : ( n2383 ) ;
assign n2385 =  ( n2168 ) ? ( bv_8_82_n581 ) : ( n2384 ) ;
assign n2386 =  ( n2166 ) ? ( bv_8_59_n604 ) : ( n2385 ) ;
assign n2387 =  ( n2164 ) ? ( bv_8_214_n163 ) : ( n2386 ) ;
assign n2388 =  ( n2162 ) ? ( bv_8_179_n287 ) : ( n2387 ) ;
assign n2389 =  ( n2160 ) ? ( bv_8_41_n597 ) : ( n2388 ) ;
assign n2390 =  ( n2158 ) ? ( bv_8_227_n115 ) : ( n2389 ) ;
assign n2391 =  ( n2156 ) ? ( bv_8_47_n592 ) : ( n2390 ) ;
assign n2392 =  ( n2154 ) ? ( bv_8_132_n438 ) : ( n2391 ) ;
assign n2393 =  ( n2152 ) ? ( bv_8_83_n578 ) : ( n2392 ) ;
assign n2394 =  ( n2150 ) ? ( bv_8_209_n182 ) : ( n2393 ) ;
assign n2395 =  ( n2148 ) ? ( bv_8_0_n583 ) : ( n2394 ) ;
assign n2396 =  ( n2146 ) ? ( bv_8_237_n77 ) : ( n2395 ) ;
assign n2397 =  ( n2144 ) ? ( bv_8_32_n576 ) : ( n2396 ) ;
assign n2398 =  ( n2142 ) ? ( bv_8_252_n17 ) : ( n2397 ) ;
assign n2399 =  ( n2140 ) ? ( bv_8_177_n295 ) : ( n2398 ) ;
assign n2400 =  ( n2138 ) ? ( bv_8_91_n557 ) : ( n2399 ) ;
assign n2401 =  ( n2136 ) ? ( bv_8_106_n516 ) : ( n2400 ) ;
assign n2402 =  ( n2134 ) ? ( bv_8_203_n205 ) : ( n2401 ) ;
assign n2403 =  ( n2132 ) ? ( bv_8_190_n252 ) : ( n2402 ) ;
assign n2404 =  ( n2130 ) ? ( bv_8_57_n559 ) : ( n2403 ) ;
assign n2405 =  ( n2128 ) ? ( bv_8_74_n555 ) : ( n2404 ) ;
assign n2406 =  ( n2126 ) ? ( bv_8_76_n552 ) : ( n2405 ) ;
assign n2407 =  ( n2124 ) ? ( bv_8_88_n549 ) : ( n2406 ) ;
assign n2408 =  ( n2122 ) ? ( bv_8_207_n190 ) : ( n2407 ) ;
assign n2409 =  ( n2120 ) ? ( bv_8_208_n186 ) : ( n2408 ) ;
assign n2410 =  ( n2118 ) ? ( bv_8_239_n69 ) : ( n2409 ) ;
assign n2411 =  ( n2116 ) ? ( bv_8_170_n318 ) : ( n2410 ) ;
assign n2412 =  ( n2114 ) ? ( bv_8_251_n21 ) : ( n2411 ) ;
assign n2413 =  ( n2112 ) ? ( bv_8_67_n535 ) : ( n2412 ) ;
assign n2414 =  ( n2110 ) ? ( bv_8_77_n532 ) : ( n2413 ) ;
assign n2415 =  ( n2108 ) ? ( bv_8_51_n529 ) : ( n2414 ) ;
assign n2416 =  ( n2106 ) ? ( bv_8_133_n435 ) : ( n2415 ) ;
assign n2417 =  ( n2104 ) ? ( bv_8_69_n523 ) : ( n2416 ) ;
assign n2418 =  ( n2102 ) ? ( bv_8_249_n29 ) : ( n2417 ) ;
assign n2419 =  ( n2100 ) ? ( bv_8_2_n518 ) : ( n2418 ) ;
assign n2420 =  ( n2098 ) ? ( bv_8_127_n455 ) : ( n2419 ) ;
assign n2421 =  ( n2096 ) ? ( bv_8_80_n511 ) : ( n2420 ) ;
assign n2422 =  ( n2094 ) ? ( bv_8_60_n508 ) : ( n2421 ) ;
assign n2423 =  ( n2092 ) ? ( bv_8_159_n355 ) : ( n2422 ) ;
assign n2424 =  ( n2090 ) ? ( bv_8_168_n323 ) : ( n2423 ) ;
assign n2425 =  ( n2088 ) ? ( bv_8_81_n499 ) : ( n2424 ) ;
assign n2426 =  ( n2086 ) ? ( bv_8_163_n341 ) : ( n2425 ) ;
assign n2427 =  ( n2084 ) ? ( bv_8_64_n493 ) : ( n2426 ) ;
assign n2428 =  ( n2082 ) ? ( bv_8_143_n406 ) : ( n2427 ) ;
assign n2429 =  ( n2080 ) ? ( bv_8_146_n396 ) : ( n2428 ) ;
assign n2430 =  ( n2078 ) ? ( bv_8_157_n361 ) : ( n2429 ) ;
assign n2431 =  ( n2076 ) ? ( bv_8_56_n482 ) : ( n2430 ) ;
assign n2432 =  ( n2074 ) ? ( bv_8_245_n45 ) : ( n2431 ) ;
assign n2433 =  ( n2072 ) ? ( bv_8_188_n259 ) : ( n2432 ) ;
assign n2434 =  ( n2070 ) ? ( bv_8_182_n278 ) : ( n2433 ) ;
assign n2435 =  ( n2068 ) ? ( bv_8_218_n148 ) : ( n2434 ) ;
assign n2436 =  ( n2066 ) ? ( bv_8_33_n469 ) : ( n2435 ) ;
assign n2437 =  ( n2064 ) ? ( bv_8_16_n465 ) : ( n2436 ) ;
assign n2438 =  ( n2062 ) ? ( bv_8_255_n5 ) : ( n2437 ) ;
assign n2439 =  ( n2060 ) ? ( bv_8_243_n53 ) : ( n2438 ) ;
assign n2440 =  ( n2058 ) ? ( bv_8_210_n178 ) : ( n2439 ) ;
assign n2441 =  ( n2056 ) ? ( bv_8_205_n197 ) : ( n2440 ) ;
assign n2442 =  ( n2054 ) ? ( bv_8_12_n450 ) : ( n2441 ) ;
assign n2443 =  ( n2052 ) ? ( bv_8_19_n447 ) : ( n2442 ) ;
assign n2444 =  ( n2050 ) ? ( bv_8_236_n81 ) : ( n2443 ) ;
assign n2445 =  ( n2048 ) ? ( bv_8_95_n440 ) : ( n2444 ) ;
assign n2446 =  ( n2046 ) ? ( bv_8_151_n379 ) : ( n2445 ) ;
assign n2447 =  ( n2044 ) ? ( bv_8_68_n433 ) : ( n2446 ) ;
assign n2448 =  ( n2042 ) ? ( bv_8_23_n430 ) : ( n2447 ) ;
assign n2449 =  ( n2040 ) ? ( bv_8_196_n230 ) : ( n2448 ) ;
assign n2450 =  ( n2038 ) ? ( bv_8_167_n326 ) : ( n2449 ) ;
assign n2451 =  ( n2036 ) ? ( bv_8_126_n423 ) : ( n2450 ) ;
assign n2452 =  ( n2034 ) ? ( bv_8_61_n420 ) : ( n2451 ) ;
assign n2453 =  ( n2032 ) ? ( bv_8_100_n417 ) : ( n2452 ) ;
assign n2454 =  ( n2030 ) ? ( bv_8_93_n414 ) : ( n2453 ) ;
assign n2455 =  ( n2028 ) ? ( bv_8_25_n411 ) : ( n2454 ) ;
assign n2456 =  ( n2026 ) ? ( bv_8_115_n408 ) : ( n2455 ) ;
assign n2457 =  ( n2024 ) ? ( bv_8_96_n404 ) : ( n2456 ) ;
assign n2458 =  ( n2022 ) ? ( bv_8_129_n401 ) : ( n2457 ) ;
assign n2459 =  ( n2020 ) ? ( bv_8_79_n398 ) : ( n2458 ) ;
assign n2460 =  ( n2018 ) ? ( bv_8_220_n140 ) : ( n2459 ) ;
assign n2461 =  ( n2016 ) ? ( bv_8_34_n391 ) : ( n2460 ) ;
assign n2462 =  ( n2014 ) ? ( bv_8_42_n388 ) : ( n2461 ) ;
assign n2463 =  ( n2012 ) ? ( bv_8_144_n385 ) : ( n2462 ) ;
assign n2464 =  ( n2010 ) ? ( bv_8_136_n381 ) : ( n2463 ) ;
assign n2465 =  ( n2008 ) ? ( bv_8_70_n377 ) : ( n2464 ) ;
assign n2466 =  ( n2006 ) ? ( bv_8_238_n73 ) : ( n2465 ) ;
assign n2467 =  ( n2004 ) ? ( bv_8_184_n270 ) : ( n2466 ) ;
assign n2468 =  ( n2002 ) ? ( bv_8_20_n369 ) : ( n2467 ) ;
assign n2469 =  ( n2000 ) ? ( bv_8_222_n132 ) : ( n2468 ) ;
assign n2470 =  ( n1998 ) ? ( bv_8_94_n363 ) : ( n2469 ) ;
assign n2471 =  ( n1996 ) ? ( bv_8_11_n359 ) : ( n2470 ) ;
assign n2472 =  ( n1994 ) ? ( bv_8_219_n144 ) : ( n2471 ) ;
assign n2473 =  ( n1992 ) ? ( bv_8_224_n126 ) : ( n2472 ) ;
assign n2474 =  ( n1990 ) ? ( bv_8_50_n350 ) : ( n2473 ) ;
assign n2475 =  ( n1988 ) ? ( bv_8_58_n347 ) : ( n2474 ) ;
assign n2476 =  ( n1986 ) ? ( bv_8_10_n343 ) : ( n2475 ) ;
assign n2477 =  ( n1984 ) ? ( bv_8_73_n339 ) : ( n2476 ) ;
assign n2478 =  ( n1982 ) ? ( bv_8_6_n335 ) : ( n2477 ) ;
assign n2479 =  ( n1980 ) ? ( bv_8_36_n331 ) : ( n2478 ) ;
assign n2480 =  ( n1978 ) ? ( bv_8_92_n328 ) : ( n2479 ) ;
assign n2481 =  ( n1976 ) ? ( bv_8_194_n238 ) : ( n2480 ) ;
assign n2482 =  ( n1974 ) ? ( bv_8_211_n174 ) : ( n2481 ) ;
assign n2483 =  ( n1972 ) ? ( bv_8_172_n310 ) : ( n2482 ) ;
assign n2484 =  ( n1970 ) ? ( bv_8_98_n316 ) : ( n2483 ) ;
assign n2485 =  ( n1968 ) ? ( bv_8_145_n312 ) : ( n2484 ) ;
assign n2486 =  ( n1966 ) ? ( bv_8_149_n308 ) : ( n2485 ) ;
assign n2487 =  ( n1964 ) ? ( bv_8_228_n111 ) : ( n2486 ) ;
assign n2488 =  ( n1962 ) ? ( bv_8_121_n302 ) : ( n2487 ) ;
assign n2489 =  ( n1960 ) ? ( bv_8_231_n100 ) : ( n2488 ) ;
assign n2490 =  ( n1958 ) ? ( bv_8_200_n216 ) : ( n2489 ) ;
assign n2491 =  ( n1956 ) ? ( bv_8_55_n293 ) : ( n2490 ) ;
assign n2492 =  ( n1954 ) ? ( bv_8_109_n289 ) : ( n2491 ) ;
assign n2493 =  ( n1952 ) ? ( bv_8_141_n285 ) : ( n2492 ) ;
assign n2494 =  ( n1950 ) ? ( bv_8_213_n166 ) : ( n2493 ) ;
assign n2495 =  ( n1948 ) ? ( bv_8_78_n280 ) : ( n2494 ) ;
assign n2496 =  ( n1946 ) ? ( bv_8_169_n276 ) : ( n2495 ) ;
assign n2497 =  ( n1944 ) ? ( bv_8_108_n272 ) : ( n2496 ) ;
assign n2498 =  ( n1942 ) ? ( bv_8_86_n268 ) : ( n2497 ) ;
assign n2499 =  ( n1940 ) ? ( bv_8_244_n49 ) : ( n2498 ) ;
assign n2500 =  ( n1938 ) ? ( bv_8_234_n89 ) : ( n2499 ) ;
assign n2501 =  ( n1936 ) ? ( bv_8_101_n261 ) : ( n2500 ) ;
assign n2502 =  ( n1934 ) ? ( bv_8_122_n257 ) : ( n2501 ) ;
assign n2503 =  ( n1932 ) ? ( bv_8_174_n254 ) : ( n2502 ) ;
assign n2504 =  ( n1930 ) ? ( bv_8_8_n250 ) : ( n2503 ) ;
assign n2505 =  ( n1928 ) ? ( bv_8_186_n247 ) : ( n2504 ) ;
assign n2506 =  ( n1926 ) ? ( bv_8_120_n243 ) : ( n2505 ) ;
assign n2507 =  ( n1924 ) ? ( bv_8_37_n240 ) : ( n2506 ) ;
assign n2508 =  ( n1922 ) ? ( bv_8_46_n236 ) : ( n2507 ) ;
assign n2509 =  ( n1920 ) ? ( bv_8_28_n232 ) : ( n2508 ) ;
assign n2510 =  ( n1918 ) ? ( bv_8_166_n228 ) : ( n2509 ) ;
assign n2511 =  ( n1916 ) ? ( bv_8_180_n224 ) : ( n2510 ) ;
assign n2512 =  ( n1914 ) ? ( bv_8_198_n221 ) : ( n2511 ) ;
assign n2513 =  ( n1912 ) ? ( bv_8_232_n96 ) : ( n2512 ) ;
assign n2514 =  ( n1910 ) ? ( bv_8_221_n136 ) : ( n2513 ) ;
assign n2515 =  ( n1908 ) ? ( bv_8_116_n211 ) : ( n2514 ) ;
assign n2516 =  ( n1906 ) ? ( bv_8_31_n207 ) : ( n2515 ) ;
assign n2517 =  ( n1904 ) ? ( bv_8_75_n203 ) : ( n2516 ) ;
assign n2518 =  ( n1902 ) ? ( bv_8_189_n199 ) : ( n2517 ) ;
assign n2519 =  ( n1900 ) ? ( bv_8_139_n195 ) : ( n2518 ) ;
assign n2520 =  ( n1898 ) ? ( bv_8_138_n192 ) : ( n2519 ) ;
assign n2521 =  ( n1896 ) ? ( bv_8_112_n188 ) : ( n2520 ) ;
assign n2522 =  ( n1894 ) ? ( bv_8_62_n184 ) : ( n2521 ) ;
assign n2523 =  ( n1892 ) ? ( bv_8_181_n180 ) : ( n2522 ) ;
assign n2524 =  ( n1890 ) ? ( bv_8_102_n176 ) : ( n2523 ) ;
assign n2525 =  ( n1888 ) ? ( bv_8_72_n172 ) : ( n2524 ) ;
assign n2526 =  ( n1886 ) ? ( bv_8_3_n168 ) : ( n2525 ) ;
assign n2527 =  ( n1884 ) ? ( bv_8_246_n41 ) : ( n2526 ) ;
assign n2528 =  ( n1882 ) ? ( bv_8_14_n161 ) : ( n2527 ) ;
assign n2529 =  ( n1880 ) ? ( bv_8_97_n157 ) : ( n2528 ) ;
assign n2530 =  ( n1878 ) ? ( bv_8_53_n153 ) : ( n2529 ) ;
assign n2531 =  ( n1876 ) ? ( bv_8_87_n150 ) : ( n2530 ) ;
assign n2532 =  ( n1874 ) ? ( bv_8_185_n146 ) : ( n2531 ) ;
assign n2533 =  ( n1872 ) ? ( bv_8_134_n142 ) : ( n2532 ) ;
assign n2534 =  ( n1870 ) ? ( bv_8_193_n138 ) : ( n2533 ) ;
assign n2535 =  ( n1868 ) ? ( bv_8_29_n134 ) : ( n2534 ) ;
assign n2536 =  ( n1866 ) ? ( bv_8_158_n130 ) : ( n2535 ) ;
assign n2537 =  ( n1864 ) ? ( bv_8_225_n123 ) : ( n2536 ) ;
assign n2538 =  ( n1862 ) ? ( bv_8_248_n33 ) : ( n2537 ) ;
assign n2539 =  ( n1860 ) ? ( bv_8_152_n121 ) : ( n2538 ) ;
assign n2540 =  ( n1858 ) ? ( bv_8_17_n117 ) : ( n2539 ) ;
assign n2541 =  ( n1856 ) ? ( bv_8_105_n113 ) : ( n2540 ) ;
assign n2542 =  ( n1854 ) ? ( bv_8_217_n109 ) : ( n2541 ) ;
assign n2543 =  ( n1852 ) ? ( bv_8_142_n105 ) : ( n2542 ) ;
assign n2544 =  ( n1850 ) ? ( bv_8_148_n102 ) : ( n2543 ) ;
assign n2545 =  ( n1848 ) ? ( bv_8_155_n98 ) : ( n2544 ) ;
assign n2546 =  ( n1846 ) ? ( bv_8_30_n94 ) : ( n2545 ) ;
assign n2547 =  ( n1844 ) ? ( bv_8_135_n91 ) : ( n2546 ) ;
assign n2548 =  ( n1842 ) ? ( bv_8_233_n87 ) : ( n2547 ) ;
assign n2549 =  ( n1840 ) ? ( bv_8_206_n83 ) : ( n2548 ) ;
assign n2550 =  ( n1838 ) ? ( bv_8_85_n79 ) : ( n2549 ) ;
assign n2551 =  ( n1836 ) ? ( bv_8_40_n75 ) : ( n2550 ) ;
assign n2552 =  ( n1834 ) ? ( bv_8_223_n71 ) : ( n2551 ) ;
assign n2553 =  ( n1832 ) ? ( bv_8_140_n67 ) : ( n2552 ) ;
assign n2554 =  ( n1830 ) ? ( bv_8_161_n63 ) : ( n2553 ) ;
assign n2555 =  ( n1828 ) ? ( bv_8_137_n59 ) : ( n2554 ) ;
assign n2556 =  ( n1826 ) ? ( bv_8_13_n55 ) : ( n2555 ) ;
assign n2557 =  ( n1824 ) ? ( bv_8_191_n51 ) : ( n2556 ) ;
assign n2558 =  ( n1822 ) ? ( bv_8_230_n47 ) : ( n2557 ) ;
assign n2559 =  ( n1820 ) ? ( bv_8_66_n43 ) : ( n2558 ) ;
assign n2560 =  ( n1818 ) ? ( bv_8_104_n39 ) : ( n2559 ) ;
assign n2561 =  ( n1816 ) ? ( bv_8_65_n35 ) : ( n2560 ) ;
assign n2562 =  ( n1814 ) ? ( bv_8_153_n31 ) : ( n2561 ) ;
assign n2563 =  ( n1812 ) ? ( bv_8_45_n27 ) : ( n2562 ) ;
assign n2564 =  ( n1810 ) ? ( bv_8_15_n23 ) : ( n2563 ) ;
assign n2565 =  ( n1808 ) ? ( bv_8_176_n19 ) : ( n2564 ) ;
assign n2566 =  ( n1806 ) ? ( bv_8_84_n15 ) : ( n2565 ) ;
assign n2567 =  ( n1804 ) ? ( bv_8_187_n11 ) : ( n2566 ) ;
assign n2568 =  ( n1802 ) ? ( bv_8_22_n7 ) : ( n2567 ) ;
assign n2569 =  ( n1800 ) ^ ( n2568 )  ;
assign n2570 =  { ( n1799 ) , ( n2569 ) }  ;
assign n2571 = in[103:96] ;
assign n2572 = in[31:24] ;
assign n2573 =  ( n2572 ) == ( bv_8_255_n5 )  ;
assign n2574 = in[31:24] ;
assign n2575 =  ( n2574 ) == ( bv_8_254_n9 )  ;
assign n2576 = in[31:24] ;
assign n2577 =  ( n2576 ) == ( bv_8_253_n13 )  ;
assign n2578 = in[31:24] ;
assign n2579 =  ( n2578 ) == ( bv_8_252_n17 )  ;
assign n2580 = in[31:24] ;
assign n2581 =  ( n2580 ) == ( bv_8_251_n21 )  ;
assign n2582 = in[31:24] ;
assign n2583 =  ( n2582 ) == ( bv_8_250_n25 )  ;
assign n2584 = in[31:24] ;
assign n2585 =  ( n2584 ) == ( bv_8_249_n29 )  ;
assign n2586 = in[31:24] ;
assign n2587 =  ( n2586 ) == ( bv_8_248_n33 )  ;
assign n2588 = in[31:24] ;
assign n2589 =  ( n2588 ) == ( bv_8_247_n37 )  ;
assign n2590 = in[31:24] ;
assign n2591 =  ( n2590 ) == ( bv_8_246_n41 )  ;
assign n2592 = in[31:24] ;
assign n2593 =  ( n2592 ) == ( bv_8_245_n45 )  ;
assign n2594 = in[31:24] ;
assign n2595 =  ( n2594 ) == ( bv_8_244_n49 )  ;
assign n2596 = in[31:24] ;
assign n2597 =  ( n2596 ) == ( bv_8_243_n53 )  ;
assign n2598 = in[31:24] ;
assign n2599 =  ( n2598 ) == ( bv_8_242_n57 )  ;
assign n2600 = in[31:24] ;
assign n2601 =  ( n2600 ) == ( bv_8_241_n61 )  ;
assign n2602 = in[31:24] ;
assign n2603 =  ( n2602 ) == ( bv_8_240_n65 )  ;
assign n2604 = in[31:24] ;
assign n2605 =  ( n2604 ) == ( bv_8_239_n69 )  ;
assign n2606 = in[31:24] ;
assign n2607 =  ( n2606 ) == ( bv_8_238_n73 )  ;
assign n2608 = in[31:24] ;
assign n2609 =  ( n2608 ) == ( bv_8_237_n77 )  ;
assign n2610 = in[31:24] ;
assign n2611 =  ( n2610 ) == ( bv_8_236_n81 )  ;
assign n2612 = in[31:24] ;
assign n2613 =  ( n2612 ) == ( bv_8_235_n85 )  ;
assign n2614 = in[31:24] ;
assign n2615 =  ( n2614 ) == ( bv_8_234_n89 )  ;
assign n2616 = in[31:24] ;
assign n2617 =  ( n2616 ) == ( bv_8_233_n87 )  ;
assign n2618 = in[31:24] ;
assign n2619 =  ( n2618 ) == ( bv_8_232_n96 )  ;
assign n2620 = in[31:24] ;
assign n2621 =  ( n2620 ) == ( bv_8_231_n100 )  ;
assign n2622 = in[31:24] ;
assign n2623 =  ( n2622 ) == ( bv_8_230_n47 )  ;
assign n2624 = in[31:24] ;
assign n2625 =  ( n2624 ) == ( bv_8_229_n107 )  ;
assign n2626 = in[31:24] ;
assign n2627 =  ( n2626 ) == ( bv_8_228_n111 )  ;
assign n2628 = in[31:24] ;
assign n2629 =  ( n2628 ) == ( bv_8_227_n115 )  ;
assign n2630 = in[31:24] ;
assign n2631 =  ( n2630 ) == ( bv_8_226_n119 )  ;
assign n2632 = in[31:24] ;
assign n2633 =  ( n2632 ) == ( bv_8_225_n123 )  ;
assign n2634 = in[31:24] ;
assign n2635 =  ( n2634 ) == ( bv_8_224_n126 )  ;
assign n2636 = in[31:24] ;
assign n2637 =  ( n2636 ) == ( bv_8_223_n71 )  ;
assign n2638 = in[31:24] ;
assign n2639 =  ( n2638 ) == ( bv_8_222_n132 )  ;
assign n2640 = in[31:24] ;
assign n2641 =  ( n2640 ) == ( bv_8_221_n136 )  ;
assign n2642 = in[31:24] ;
assign n2643 =  ( n2642 ) == ( bv_8_220_n140 )  ;
assign n2644 = in[31:24] ;
assign n2645 =  ( n2644 ) == ( bv_8_219_n144 )  ;
assign n2646 = in[31:24] ;
assign n2647 =  ( n2646 ) == ( bv_8_218_n148 )  ;
assign n2648 = in[31:24] ;
assign n2649 =  ( n2648 ) == ( bv_8_217_n109 )  ;
assign n2650 = in[31:24] ;
assign n2651 =  ( n2650 ) == ( bv_8_216_n155 )  ;
assign n2652 = in[31:24] ;
assign n2653 =  ( n2652 ) == ( bv_8_215_n159 )  ;
assign n2654 = in[31:24] ;
assign n2655 =  ( n2654 ) == ( bv_8_214_n163 )  ;
assign n2656 = in[31:24] ;
assign n2657 =  ( n2656 ) == ( bv_8_213_n166 )  ;
assign n2658 = in[31:24] ;
assign n2659 =  ( n2658 ) == ( bv_8_212_n170 )  ;
assign n2660 = in[31:24] ;
assign n2661 =  ( n2660 ) == ( bv_8_211_n174 )  ;
assign n2662 = in[31:24] ;
assign n2663 =  ( n2662 ) == ( bv_8_210_n178 )  ;
assign n2664 = in[31:24] ;
assign n2665 =  ( n2664 ) == ( bv_8_209_n182 )  ;
assign n2666 = in[31:24] ;
assign n2667 =  ( n2666 ) == ( bv_8_208_n186 )  ;
assign n2668 = in[31:24] ;
assign n2669 =  ( n2668 ) == ( bv_8_207_n190 )  ;
assign n2670 = in[31:24] ;
assign n2671 =  ( n2670 ) == ( bv_8_206_n83 )  ;
assign n2672 = in[31:24] ;
assign n2673 =  ( n2672 ) == ( bv_8_205_n197 )  ;
assign n2674 = in[31:24] ;
assign n2675 =  ( n2674 ) == ( bv_8_204_n201 )  ;
assign n2676 = in[31:24] ;
assign n2677 =  ( n2676 ) == ( bv_8_203_n205 )  ;
assign n2678 = in[31:24] ;
assign n2679 =  ( n2678 ) == ( bv_8_202_n209 )  ;
assign n2680 = in[31:24] ;
assign n2681 =  ( n2680 ) == ( bv_8_201_n213 )  ;
assign n2682 = in[31:24] ;
assign n2683 =  ( n2682 ) == ( bv_8_200_n216 )  ;
assign n2684 = in[31:24] ;
assign n2685 =  ( n2684 ) == ( bv_8_199_n219 )  ;
assign n2686 = in[31:24] ;
assign n2687 =  ( n2686 ) == ( bv_8_198_n221 )  ;
assign n2688 = in[31:24] ;
assign n2689 =  ( n2688 ) == ( bv_8_197_n226 )  ;
assign n2690 = in[31:24] ;
assign n2691 =  ( n2690 ) == ( bv_8_196_n230 )  ;
assign n2692 = in[31:24] ;
assign n2693 =  ( n2692 ) == ( bv_8_195_n234 )  ;
assign n2694 = in[31:24] ;
assign n2695 =  ( n2694 ) == ( bv_8_194_n238 )  ;
assign n2696 = in[31:24] ;
assign n2697 =  ( n2696 ) == ( bv_8_193_n138 )  ;
assign n2698 = in[31:24] ;
assign n2699 =  ( n2698 ) == ( bv_8_192_n245 )  ;
assign n2700 = in[31:24] ;
assign n2701 =  ( n2700 ) == ( bv_8_191_n51 )  ;
assign n2702 = in[31:24] ;
assign n2703 =  ( n2702 ) == ( bv_8_190_n252 )  ;
assign n2704 = in[31:24] ;
assign n2705 =  ( n2704 ) == ( bv_8_189_n199 )  ;
assign n2706 = in[31:24] ;
assign n2707 =  ( n2706 ) == ( bv_8_188_n259 )  ;
assign n2708 = in[31:24] ;
assign n2709 =  ( n2708 ) == ( bv_8_187_n11 )  ;
assign n2710 = in[31:24] ;
assign n2711 =  ( n2710 ) == ( bv_8_186_n247 )  ;
assign n2712 = in[31:24] ;
assign n2713 =  ( n2712 ) == ( bv_8_185_n146 )  ;
assign n2714 = in[31:24] ;
assign n2715 =  ( n2714 ) == ( bv_8_184_n270 )  ;
assign n2716 = in[31:24] ;
assign n2717 =  ( n2716 ) == ( bv_8_183_n274 )  ;
assign n2718 = in[31:24] ;
assign n2719 =  ( n2718 ) == ( bv_8_182_n278 )  ;
assign n2720 = in[31:24] ;
assign n2721 =  ( n2720 ) == ( bv_8_181_n180 )  ;
assign n2722 = in[31:24] ;
assign n2723 =  ( n2722 ) == ( bv_8_180_n224 )  ;
assign n2724 = in[31:24] ;
assign n2725 =  ( n2724 ) == ( bv_8_179_n287 )  ;
assign n2726 = in[31:24] ;
assign n2727 =  ( n2726 ) == ( bv_8_178_n291 )  ;
assign n2728 = in[31:24] ;
assign n2729 =  ( n2728 ) == ( bv_8_177_n295 )  ;
assign n2730 = in[31:24] ;
assign n2731 =  ( n2730 ) == ( bv_8_176_n19 )  ;
assign n2732 = in[31:24] ;
assign n2733 =  ( n2732 ) == ( bv_8_175_n300 )  ;
assign n2734 = in[31:24] ;
assign n2735 =  ( n2734 ) == ( bv_8_174_n254 )  ;
assign n2736 = in[31:24] ;
assign n2737 =  ( n2736 ) == ( bv_8_173_n306 )  ;
assign n2738 = in[31:24] ;
assign n2739 =  ( n2738 ) == ( bv_8_172_n310 )  ;
assign n2740 = in[31:24] ;
assign n2741 =  ( n2740 ) == ( bv_8_171_n314 )  ;
assign n2742 = in[31:24] ;
assign n2743 =  ( n2742 ) == ( bv_8_170_n318 )  ;
assign n2744 = in[31:24] ;
assign n2745 =  ( n2744 ) == ( bv_8_169_n276 )  ;
assign n2746 = in[31:24] ;
assign n2747 =  ( n2746 ) == ( bv_8_168_n323 )  ;
assign n2748 = in[31:24] ;
assign n2749 =  ( n2748 ) == ( bv_8_167_n326 )  ;
assign n2750 = in[31:24] ;
assign n2751 =  ( n2750 ) == ( bv_8_166_n228 )  ;
assign n2752 = in[31:24] ;
assign n2753 =  ( n2752 ) == ( bv_8_165_n333 )  ;
assign n2754 = in[31:24] ;
assign n2755 =  ( n2754 ) == ( bv_8_164_n337 )  ;
assign n2756 = in[31:24] ;
assign n2757 =  ( n2756 ) == ( bv_8_163_n341 )  ;
assign n2758 = in[31:24] ;
assign n2759 =  ( n2758 ) == ( bv_8_162_n345 )  ;
assign n2760 = in[31:24] ;
assign n2761 =  ( n2760 ) == ( bv_8_161_n63 )  ;
assign n2762 = in[31:24] ;
assign n2763 =  ( n2762 ) == ( bv_8_160_n352 )  ;
assign n2764 = in[31:24] ;
assign n2765 =  ( n2764 ) == ( bv_8_159_n355 )  ;
assign n2766 = in[31:24] ;
assign n2767 =  ( n2766 ) == ( bv_8_158_n130 )  ;
assign n2768 = in[31:24] ;
assign n2769 =  ( n2768 ) == ( bv_8_157_n361 )  ;
assign n2770 = in[31:24] ;
assign n2771 =  ( n2770 ) == ( bv_8_156_n365 )  ;
assign n2772 = in[31:24] ;
assign n2773 =  ( n2772 ) == ( bv_8_155_n98 )  ;
assign n2774 = in[31:24] ;
assign n2775 =  ( n2774 ) == ( bv_8_154_n371 )  ;
assign n2776 = in[31:24] ;
assign n2777 =  ( n2776 ) == ( bv_8_153_n31 )  ;
assign n2778 = in[31:24] ;
assign n2779 =  ( n2778 ) == ( bv_8_152_n121 )  ;
assign n2780 = in[31:24] ;
assign n2781 =  ( n2780 ) == ( bv_8_151_n379 )  ;
assign n2782 = in[31:24] ;
assign n2783 =  ( n2782 ) == ( bv_8_150_n383 )  ;
assign n2784 = in[31:24] ;
assign n2785 =  ( n2784 ) == ( bv_8_149_n308 )  ;
assign n2786 = in[31:24] ;
assign n2787 =  ( n2786 ) == ( bv_8_148_n102 )  ;
assign n2788 = in[31:24] ;
assign n2789 =  ( n2788 ) == ( bv_8_147_n393 )  ;
assign n2790 = in[31:24] ;
assign n2791 =  ( n2790 ) == ( bv_8_146_n396 )  ;
assign n2792 = in[31:24] ;
assign n2793 =  ( n2792 ) == ( bv_8_145_n312 )  ;
assign n2794 = in[31:24] ;
assign n2795 =  ( n2794 ) == ( bv_8_144_n385 )  ;
assign n2796 = in[31:24] ;
assign n2797 =  ( n2796 ) == ( bv_8_143_n406 )  ;
assign n2798 = in[31:24] ;
assign n2799 =  ( n2798 ) == ( bv_8_142_n105 )  ;
assign n2800 = in[31:24] ;
assign n2801 =  ( n2800 ) == ( bv_8_141_n285 )  ;
assign n2802 = in[31:24] ;
assign n2803 =  ( n2802 ) == ( bv_8_140_n67 )  ;
assign n2804 = in[31:24] ;
assign n2805 =  ( n2804 ) == ( bv_8_139_n195 )  ;
assign n2806 = in[31:24] ;
assign n2807 =  ( n2806 ) == ( bv_8_138_n192 )  ;
assign n2808 = in[31:24] ;
assign n2809 =  ( n2808 ) == ( bv_8_137_n59 )  ;
assign n2810 = in[31:24] ;
assign n2811 =  ( n2810 ) == ( bv_8_136_n381 )  ;
assign n2812 = in[31:24] ;
assign n2813 =  ( n2812 ) == ( bv_8_135_n91 )  ;
assign n2814 = in[31:24] ;
assign n2815 =  ( n2814 ) == ( bv_8_134_n142 )  ;
assign n2816 = in[31:24] ;
assign n2817 =  ( n2816 ) == ( bv_8_133_n435 )  ;
assign n2818 = in[31:24] ;
assign n2819 =  ( n2818 ) == ( bv_8_132_n438 )  ;
assign n2820 = in[31:24] ;
assign n2821 =  ( n2820 ) == ( bv_8_131_n442 )  ;
assign n2822 = in[31:24] ;
assign n2823 =  ( n2822 ) == ( bv_8_130_n445 )  ;
assign n2824 = in[31:24] ;
assign n2825 =  ( n2824 ) == ( bv_8_129_n401 )  ;
assign n2826 = in[31:24] ;
assign n2827 =  ( n2826 ) == ( bv_8_128_n452 )  ;
assign n2828 = in[31:24] ;
assign n2829 =  ( n2828 ) == ( bv_8_127_n455 )  ;
assign n2830 = in[31:24] ;
assign n2831 =  ( n2830 ) == ( bv_8_126_n423 )  ;
assign n2832 = in[31:24] ;
assign n2833 =  ( n2832 ) == ( bv_8_125_n460 )  ;
assign n2834 = in[31:24] ;
assign n2835 =  ( n2834 ) == ( bv_8_124_n463 )  ;
assign n2836 = in[31:24] ;
assign n2837 =  ( n2836 ) == ( bv_8_123_n467 )  ;
assign n2838 = in[31:24] ;
assign n2839 =  ( n2838 ) == ( bv_8_122_n257 )  ;
assign n2840 = in[31:24] ;
assign n2841 =  ( n2840 ) == ( bv_8_121_n302 )  ;
assign n2842 = in[31:24] ;
assign n2843 =  ( n2842 ) == ( bv_8_120_n243 )  ;
assign n2844 = in[31:24] ;
assign n2845 =  ( n2844 ) == ( bv_8_119_n477 )  ;
assign n2846 = in[31:24] ;
assign n2847 =  ( n2846 ) == ( bv_8_118_n480 )  ;
assign n2848 = in[31:24] ;
assign n2849 =  ( n2848 ) == ( bv_8_117_n484 )  ;
assign n2850 = in[31:24] ;
assign n2851 =  ( n2850 ) == ( bv_8_116_n211 )  ;
assign n2852 = in[31:24] ;
assign n2853 =  ( n2852 ) == ( bv_8_115_n408 )  ;
assign n2854 = in[31:24] ;
assign n2855 =  ( n2854 ) == ( bv_8_114_n491 )  ;
assign n2856 = in[31:24] ;
assign n2857 =  ( n2856 ) == ( bv_8_113_n495 )  ;
assign n2858 = in[31:24] ;
assign n2859 =  ( n2858 ) == ( bv_8_112_n188 )  ;
assign n2860 = in[31:24] ;
assign n2861 =  ( n2860 ) == ( bv_8_111_n501 )  ;
assign n2862 = in[31:24] ;
assign n2863 =  ( n2862 ) == ( bv_8_110_n504 )  ;
assign n2864 = in[31:24] ;
assign n2865 =  ( n2864 ) == ( bv_8_109_n289 )  ;
assign n2866 = in[31:24] ;
assign n2867 =  ( n2866 ) == ( bv_8_108_n272 )  ;
assign n2868 = in[31:24] ;
assign n2869 =  ( n2868 ) == ( bv_8_107_n513 )  ;
assign n2870 = in[31:24] ;
assign n2871 =  ( n2870 ) == ( bv_8_106_n516 )  ;
assign n2872 = in[31:24] ;
assign n2873 =  ( n2872 ) == ( bv_8_105_n113 )  ;
assign n2874 = in[31:24] ;
assign n2875 =  ( n2874 ) == ( bv_8_104_n39 )  ;
assign n2876 = in[31:24] ;
assign n2877 =  ( n2876 ) == ( bv_8_103_n525 )  ;
assign n2878 = in[31:24] ;
assign n2879 =  ( n2878 ) == ( bv_8_102_n176 )  ;
assign n2880 = in[31:24] ;
assign n2881 =  ( n2880 ) == ( bv_8_101_n261 )  ;
assign n2882 = in[31:24] ;
assign n2883 =  ( n2882 ) == ( bv_8_100_n417 )  ;
assign n2884 = in[31:24] ;
assign n2885 =  ( n2884 ) == ( bv_8_99_n537 )  ;
assign n2886 = in[31:24] ;
assign n2887 =  ( n2886 ) == ( bv_8_98_n316 )  ;
assign n2888 = in[31:24] ;
assign n2889 =  ( n2888 ) == ( bv_8_97_n157 )  ;
assign n2890 = in[31:24] ;
assign n2891 =  ( n2890 ) == ( bv_8_96_n404 )  ;
assign n2892 = in[31:24] ;
assign n2893 =  ( n2892 ) == ( bv_8_95_n440 )  ;
assign n2894 = in[31:24] ;
assign n2895 =  ( n2894 ) == ( bv_8_94_n363 )  ;
assign n2896 = in[31:24] ;
assign n2897 =  ( n2896 ) == ( bv_8_93_n414 )  ;
assign n2898 = in[31:24] ;
assign n2899 =  ( n2898 ) == ( bv_8_92_n328 )  ;
assign n2900 = in[31:24] ;
assign n2901 =  ( n2900 ) == ( bv_8_91_n557 )  ;
assign n2902 = in[31:24] ;
assign n2903 =  ( n2902 ) == ( bv_8_90_n561 )  ;
assign n2904 = in[31:24] ;
assign n2905 =  ( n2904 ) == ( bv_8_89_n564 )  ;
assign n2906 = in[31:24] ;
assign n2907 =  ( n2906 ) == ( bv_8_88_n549 )  ;
assign n2908 = in[31:24] ;
assign n2909 =  ( n2908 ) == ( bv_8_87_n150 )  ;
assign n2910 = in[31:24] ;
assign n2911 =  ( n2910 ) == ( bv_8_86_n268 )  ;
assign n2912 = in[31:24] ;
assign n2913 =  ( n2912 ) == ( bv_8_85_n79 )  ;
assign n2914 = in[31:24] ;
assign n2915 =  ( n2914 ) == ( bv_8_84_n15 )  ;
assign n2916 = in[31:24] ;
assign n2917 =  ( n2916 ) == ( bv_8_83_n578 )  ;
assign n2918 = in[31:24] ;
assign n2919 =  ( n2918 ) == ( bv_8_82_n581 )  ;
assign n2920 = in[31:24] ;
assign n2921 =  ( n2920 ) == ( bv_8_81_n499 )  ;
assign n2922 = in[31:24] ;
assign n2923 =  ( n2922 ) == ( bv_8_80_n511 )  ;
assign n2924 = in[31:24] ;
assign n2925 =  ( n2924 ) == ( bv_8_79_n398 )  ;
assign n2926 = in[31:24] ;
assign n2927 =  ( n2926 ) == ( bv_8_78_n280 )  ;
assign n2928 = in[31:24] ;
assign n2929 =  ( n2928 ) == ( bv_8_77_n532 )  ;
assign n2930 = in[31:24] ;
assign n2931 =  ( n2930 ) == ( bv_8_76_n552 )  ;
assign n2932 = in[31:24] ;
assign n2933 =  ( n2932 ) == ( bv_8_75_n203 )  ;
assign n2934 = in[31:24] ;
assign n2935 =  ( n2934 ) == ( bv_8_74_n555 )  ;
assign n2936 = in[31:24] ;
assign n2937 =  ( n2936 ) == ( bv_8_73_n339 )  ;
assign n2938 = in[31:24] ;
assign n2939 =  ( n2938 ) == ( bv_8_72_n172 )  ;
assign n2940 = in[31:24] ;
assign n2941 =  ( n2940 ) == ( bv_8_71_n608 )  ;
assign n2942 = in[31:24] ;
assign n2943 =  ( n2942 ) == ( bv_8_70_n377 )  ;
assign n2944 = in[31:24] ;
assign n2945 =  ( n2944 ) == ( bv_8_69_n523 )  ;
assign n2946 = in[31:24] ;
assign n2947 =  ( n2946 ) == ( bv_8_68_n433 )  ;
assign n2948 = in[31:24] ;
assign n2949 =  ( n2948 ) == ( bv_8_67_n535 )  ;
assign n2950 = in[31:24] ;
assign n2951 =  ( n2950 ) == ( bv_8_66_n43 )  ;
assign n2952 = in[31:24] ;
assign n2953 =  ( n2952 ) == ( bv_8_65_n35 )  ;
assign n2954 = in[31:24] ;
assign n2955 =  ( n2954 ) == ( bv_8_64_n493 )  ;
assign n2956 = in[31:24] ;
assign n2957 =  ( n2956 ) == ( bv_8_63_n629 )  ;
assign n2958 = in[31:24] ;
assign n2959 =  ( n2958 ) == ( bv_8_62_n184 )  ;
assign n2960 = in[31:24] ;
assign n2961 =  ( n2960 ) == ( bv_8_61_n420 )  ;
assign n2962 = in[31:24] ;
assign n2963 =  ( n2962 ) == ( bv_8_60_n508 )  ;
assign n2964 = in[31:24] ;
assign n2965 =  ( n2964 ) == ( bv_8_59_n604 )  ;
assign n2966 = in[31:24] ;
assign n2967 =  ( n2966 ) == ( bv_8_58_n347 )  ;
assign n2968 = in[31:24] ;
assign n2969 =  ( n2968 ) == ( bv_8_57_n559 )  ;
assign n2970 = in[31:24] ;
assign n2971 =  ( n2970 ) == ( bv_8_56_n482 )  ;
assign n2972 = in[31:24] ;
assign n2973 =  ( n2972 ) == ( bv_8_55_n293 )  ;
assign n2974 = in[31:24] ;
assign n2975 =  ( n2974 ) == ( bv_8_54_n651 )  ;
assign n2976 = in[31:24] ;
assign n2977 =  ( n2976 ) == ( bv_8_53_n153 )  ;
assign n2978 = in[31:24] ;
assign n2979 =  ( n2978 ) == ( bv_8_52_n657 )  ;
assign n2980 = in[31:24] ;
assign n2981 =  ( n2980 ) == ( bv_8_51_n529 )  ;
assign n2982 = in[31:24] ;
assign n2983 =  ( n2982 ) == ( bv_8_50_n350 )  ;
assign n2984 = in[31:24] ;
assign n2985 =  ( n2984 ) == ( bv_8_49_n666 )  ;
assign n2986 = in[31:24] ;
assign n2987 =  ( n2986 ) == ( bv_8_48_n669 )  ;
assign n2988 = in[31:24] ;
assign n2989 =  ( n2988 ) == ( bv_8_47_n592 )  ;
assign n2990 = in[31:24] ;
assign n2991 =  ( n2990 ) == ( bv_8_46_n236 )  ;
assign n2992 = in[31:24] ;
assign n2993 =  ( n2992 ) == ( bv_8_45_n27 )  ;
assign n2994 = in[31:24] ;
assign n2995 =  ( n2994 ) == ( bv_8_44_n622 )  ;
assign n2996 = in[31:24] ;
assign n2997 =  ( n2996 ) == ( bv_8_43_n682 )  ;
assign n2998 = in[31:24] ;
assign n2999 =  ( n2998 ) == ( bv_8_42_n388 )  ;
assign n3000 = in[31:24] ;
assign n3001 =  ( n3000 ) == ( bv_8_41_n597 )  ;
assign n3002 = in[31:24] ;
assign n3003 =  ( n3002 ) == ( bv_8_40_n75 )  ;
assign n3004 = in[31:24] ;
assign n3005 =  ( n3004 ) == ( bv_8_39_n635 )  ;
assign n3006 = in[31:24] ;
assign n3007 =  ( n3006 ) == ( bv_8_38_n693 )  ;
assign n3008 = in[31:24] ;
assign n3009 =  ( n3008 ) == ( bv_8_37_n240 )  ;
assign n3010 = in[31:24] ;
assign n3011 =  ( n3010 ) == ( bv_8_36_n331 )  ;
assign n3012 = in[31:24] ;
assign n3013 =  ( n3012 ) == ( bv_8_35_n664 )  ;
assign n3014 = in[31:24] ;
assign n3015 =  ( n3014 ) == ( bv_8_34_n391 )  ;
assign n3016 = in[31:24] ;
assign n3017 =  ( n3016 ) == ( bv_8_33_n469 )  ;
assign n3018 = in[31:24] ;
assign n3019 =  ( n3018 ) == ( bv_8_32_n576 )  ;
assign n3020 = in[31:24] ;
assign n3021 =  ( n3020 ) == ( bv_8_31_n207 )  ;
assign n3022 = in[31:24] ;
assign n3023 =  ( n3022 ) == ( bv_8_30_n94 )  ;
assign n3024 = in[31:24] ;
assign n3025 =  ( n3024 ) == ( bv_8_29_n134 )  ;
assign n3026 = in[31:24] ;
assign n3027 =  ( n3026 ) == ( bv_8_28_n232 )  ;
assign n3028 = in[31:24] ;
assign n3029 =  ( n3028 ) == ( bv_8_27_n616 )  ;
assign n3030 = in[31:24] ;
assign n3031 =  ( n3030 ) == ( bv_8_26_n619 )  ;
assign n3032 = in[31:24] ;
assign n3033 =  ( n3032 ) == ( bv_8_25_n411 )  ;
assign n3034 = in[31:24] ;
assign n3035 =  ( n3034 ) == ( bv_8_24_n659 )  ;
assign n3036 = in[31:24] ;
assign n3037 =  ( n3036 ) == ( bv_8_23_n430 )  ;
assign n3038 = in[31:24] ;
assign n3039 =  ( n3038 ) == ( bv_8_22_n7 )  ;
assign n3040 = in[31:24] ;
assign n3041 =  ( n3040 ) == ( bv_8_21_n674 )  ;
assign n3042 = in[31:24] ;
assign n3043 =  ( n3042 ) == ( bv_8_20_n369 )  ;
assign n3044 = in[31:24] ;
assign n3045 =  ( n3044 ) == ( bv_8_19_n447 )  ;
assign n3046 = in[31:24] ;
assign n3047 =  ( n3046 ) == ( bv_8_18_n644 )  ;
assign n3048 = in[31:24] ;
assign n3049 =  ( n3048 ) == ( bv_8_17_n117 )  ;
assign n3050 = in[31:24] ;
assign n3051 =  ( n3050 ) == ( bv_8_16_n465 )  ;
assign n3052 = in[31:24] ;
assign n3053 =  ( n3052 ) == ( bv_8_15_n23 )  ;
assign n3054 = in[31:24] ;
assign n3055 =  ( n3054 ) == ( bv_8_14_n161 )  ;
assign n3056 = in[31:24] ;
assign n3057 =  ( n3056 ) == ( bv_8_13_n55 )  ;
assign n3058 = in[31:24] ;
assign n3059 =  ( n3058 ) == ( bv_8_12_n450 )  ;
assign n3060 = in[31:24] ;
assign n3061 =  ( n3060 ) == ( bv_8_11_n359 )  ;
assign n3062 = in[31:24] ;
assign n3063 =  ( n3062 ) == ( bv_8_10_n343 )  ;
assign n3064 = in[31:24] ;
assign n3065 =  ( n3064 ) == ( bv_8_9_n627 )  ;
assign n3066 = in[31:24] ;
assign n3067 =  ( n3066 ) == ( bv_8_8_n250 )  ;
assign n3068 = in[31:24] ;
assign n3069 =  ( n3068 ) == ( bv_8_7_n647 )  ;
assign n3070 = in[31:24] ;
assign n3071 =  ( n3070 ) == ( bv_8_6_n335 )  ;
assign n3072 = in[31:24] ;
assign n3073 =  ( n3072 ) == ( bv_8_5_n653 )  ;
assign n3074 = in[31:24] ;
assign n3075 =  ( n3074 ) == ( bv_8_4_n671 )  ;
assign n3076 = in[31:24] ;
assign n3077 =  ( n3076 ) == ( bv_8_3_n168 )  ;
assign n3078 = in[31:24] ;
assign n3079 =  ( n3078 ) == ( bv_8_2_n518 )  ;
assign n3080 = in[31:24] ;
assign n3081 =  ( n3080 ) == ( bv_8_1_n753 )  ;
assign n3082 = in[31:24] ;
assign n3083 =  ( n3082 ) == ( bv_8_0_n583 )  ;
assign n3084 =  ( n3083 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n3085 =  ( n3081 ) ? ( bv_8_124_n463 ) : ( n3084 ) ;
assign n3086 =  ( n3079 ) ? ( bv_8_119_n477 ) : ( n3085 ) ;
assign n3087 =  ( n3077 ) ? ( bv_8_123_n467 ) : ( n3086 ) ;
assign n3088 =  ( n3075 ) ? ( bv_8_242_n57 ) : ( n3087 ) ;
assign n3089 =  ( n3073 ) ? ( bv_8_107_n513 ) : ( n3088 ) ;
assign n3090 =  ( n3071 ) ? ( bv_8_111_n501 ) : ( n3089 ) ;
assign n3091 =  ( n3069 ) ? ( bv_8_197_n226 ) : ( n3090 ) ;
assign n3092 =  ( n3067 ) ? ( bv_8_48_n669 ) : ( n3091 ) ;
assign n3093 =  ( n3065 ) ? ( bv_8_1_n753 ) : ( n3092 ) ;
assign n3094 =  ( n3063 ) ? ( bv_8_103_n525 ) : ( n3093 ) ;
assign n3095 =  ( n3061 ) ? ( bv_8_43_n682 ) : ( n3094 ) ;
assign n3096 =  ( n3059 ) ? ( bv_8_254_n9 ) : ( n3095 ) ;
assign n3097 =  ( n3057 ) ? ( bv_8_215_n159 ) : ( n3096 ) ;
assign n3098 =  ( n3055 ) ? ( bv_8_171_n314 ) : ( n3097 ) ;
assign n3099 =  ( n3053 ) ? ( bv_8_118_n480 ) : ( n3098 ) ;
assign n3100 =  ( n3051 ) ? ( bv_8_202_n209 ) : ( n3099 ) ;
assign n3101 =  ( n3049 ) ? ( bv_8_130_n445 ) : ( n3100 ) ;
assign n3102 =  ( n3047 ) ? ( bv_8_201_n213 ) : ( n3101 ) ;
assign n3103 =  ( n3045 ) ? ( bv_8_125_n460 ) : ( n3102 ) ;
assign n3104 =  ( n3043 ) ? ( bv_8_250_n25 ) : ( n3103 ) ;
assign n3105 =  ( n3041 ) ? ( bv_8_89_n564 ) : ( n3104 ) ;
assign n3106 =  ( n3039 ) ? ( bv_8_71_n608 ) : ( n3105 ) ;
assign n3107 =  ( n3037 ) ? ( bv_8_240_n65 ) : ( n3106 ) ;
assign n3108 =  ( n3035 ) ? ( bv_8_173_n306 ) : ( n3107 ) ;
assign n3109 =  ( n3033 ) ? ( bv_8_212_n170 ) : ( n3108 ) ;
assign n3110 =  ( n3031 ) ? ( bv_8_162_n345 ) : ( n3109 ) ;
assign n3111 =  ( n3029 ) ? ( bv_8_175_n300 ) : ( n3110 ) ;
assign n3112 =  ( n3027 ) ? ( bv_8_156_n365 ) : ( n3111 ) ;
assign n3113 =  ( n3025 ) ? ( bv_8_164_n337 ) : ( n3112 ) ;
assign n3114 =  ( n3023 ) ? ( bv_8_114_n491 ) : ( n3113 ) ;
assign n3115 =  ( n3021 ) ? ( bv_8_192_n245 ) : ( n3114 ) ;
assign n3116 =  ( n3019 ) ? ( bv_8_183_n274 ) : ( n3115 ) ;
assign n3117 =  ( n3017 ) ? ( bv_8_253_n13 ) : ( n3116 ) ;
assign n3118 =  ( n3015 ) ? ( bv_8_147_n393 ) : ( n3117 ) ;
assign n3119 =  ( n3013 ) ? ( bv_8_38_n693 ) : ( n3118 ) ;
assign n3120 =  ( n3011 ) ? ( bv_8_54_n651 ) : ( n3119 ) ;
assign n3121 =  ( n3009 ) ? ( bv_8_63_n629 ) : ( n3120 ) ;
assign n3122 =  ( n3007 ) ? ( bv_8_247_n37 ) : ( n3121 ) ;
assign n3123 =  ( n3005 ) ? ( bv_8_204_n201 ) : ( n3122 ) ;
assign n3124 =  ( n3003 ) ? ( bv_8_52_n657 ) : ( n3123 ) ;
assign n3125 =  ( n3001 ) ? ( bv_8_165_n333 ) : ( n3124 ) ;
assign n3126 =  ( n2999 ) ? ( bv_8_229_n107 ) : ( n3125 ) ;
assign n3127 =  ( n2997 ) ? ( bv_8_241_n61 ) : ( n3126 ) ;
assign n3128 =  ( n2995 ) ? ( bv_8_113_n495 ) : ( n3127 ) ;
assign n3129 =  ( n2993 ) ? ( bv_8_216_n155 ) : ( n3128 ) ;
assign n3130 =  ( n2991 ) ? ( bv_8_49_n666 ) : ( n3129 ) ;
assign n3131 =  ( n2989 ) ? ( bv_8_21_n674 ) : ( n3130 ) ;
assign n3132 =  ( n2987 ) ? ( bv_8_4_n671 ) : ( n3131 ) ;
assign n3133 =  ( n2985 ) ? ( bv_8_199_n219 ) : ( n3132 ) ;
assign n3134 =  ( n2983 ) ? ( bv_8_35_n664 ) : ( n3133 ) ;
assign n3135 =  ( n2981 ) ? ( bv_8_195_n234 ) : ( n3134 ) ;
assign n3136 =  ( n2979 ) ? ( bv_8_24_n659 ) : ( n3135 ) ;
assign n3137 =  ( n2977 ) ? ( bv_8_150_n383 ) : ( n3136 ) ;
assign n3138 =  ( n2975 ) ? ( bv_8_5_n653 ) : ( n3137 ) ;
assign n3139 =  ( n2973 ) ? ( bv_8_154_n371 ) : ( n3138 ) ;
assign n3140 =  ( n2971 ) ? ( bv_8_7_n647 ) : ( n3139 ) ;
assign n3141 =  ( n2969 ) ? ( bv_8_18_n644 ) : ( n3140 ) ;
assign n3142 =  ( n2967 ) ? ( bv_8_128_n452 ) : ( n3141 ) ;
assign n3143 =  ( n2965 ) ? ( bv_8_226_n119 ) : ( n3142 ) ;
assign n3144 =  ( n2963 ) ? ( bv_8_235_n85 ) : ( n3143 ) ;
assign n3145 =  ( n2961 ) ? ( bv_8_39_n635 ) : ( n3144 ) ;
assign n3146 =  ( n2959 ) ? ( bv_8_178_n291 ) : ( n3145 ) ;
assign n3147 =  ( n2957 ) ? ( bv_8_117_n484 ) : ( n3146 ) ;
assign n3148 =  ( n2955 ) ? ( bv_8_9_n627 ) : ( n3147 ) ;
assign n3149 =  ( n2953 ) ? ( bv_8_131_n442 ) : ( n3148 ) ;
assign n3150 =  ( n2951 ) ? ( bv_8_44_n622 ) : ( n3149 ) ;
assign n3151 =  ( n2949 ) ? ( bv_8_26_n619 ) : ( n3150 ) ;
assign n3152 =  ( n2947 ) ? ( bv_8_27_n616 ) : ( n3151 ) ;
assign n3153 =  ( n2945 ) ? ( bv_8_110_n504 ) : ( n3152 ) ;
assign n3154 =  ( n2943 ) ? ( bv_8_90_n561 ) : ( n3153 ) ;
assign n3155 =  ( n2941 ) ? ( bv_8_160_n352 ) : ( n3154 ) ;
assign n3156 =  ( n2939 ) ? ( bv_8_82_n581 ) : ( n3155 ) ;
assign n3157 =  ( n2937 ) ? ( bv_8_59_n604 ) : ( n3156 ) ;
assign n3158 =  ( n2935 ) ? ( bv_8_214_n163 ) : ( n3157 ) ;
assign n3159 =  ( n2933 ) ? ( bv_8_179_n287 ) : ( n3158 ) ;
assign n3160 =  ( n2931 ) ? ( bv_8_41_n597 ) : ( n3159 ) ;
assign n3161 =  ( n2929 ) ? ( bv_8_227_n115 ) : ( n3160 ) ;
assign n3162 =  ( n2927 ) ? ( bv_8_47_n592 ) : ( n3161 ) ;
assign n3163 =  ( n2925 ) ? ( bv_8_132_n438 ) : ( n3162 ) ;
assign n3164 =  ( n2923 ) ? ( bv_8_83_n578 ) : ( n3163 ) ;
assign n3165 =  ( n2921 ) ? ( bv_8_209_n182 ) : ( n3164 ) ;
assign n3166 =  ( n2919 ) ? ( bv_8_0_n583 ) : ( n3165 ) ;
assign n3167 =  ( n2917 ) ? ( bv_8_237_n77 ) : ( n3166 ) ;
assign n3168 =  ( n2915 ) ? ( bv_8_32_n576 ) : ( n3167 ) ;
assign n3169 =  ( n2913 ) ? ( bv_8_252_n17 ) : ( n3168 ) ;
assign n3170 =  ( n2911 ) ? ( bv_8_177_n295 ) : ( n3169 ) ;
assign n3171 =  ( n2909 ) ? ( bv_8_91_n557 ) : ( n3170 ) ;
assign n3172 =  ( n2907 ) ? ( bv_8_106_n516 ) : ( n3171 ) ;
assign n3173 =  ( n2905 ) ? ( bv_8_203_n205 ) : ( n3172 ) ;
assign n3174 =  ( n2903 ) ? ( bv_8_190_n252 ) : ( n3173 ) ;
assign n3175 =  ( n2901 ) ? ( bv_8_57_n559 ) : ( n3174 ) ;
assign n3176 =  ( n2899 ) ? ( bv_8_74_n555 ) : ( n3175 ) ;
assign n3177 =  ( n2897 ) ? ( bv_8_76_n552 ) : ( n3176 ) ;
assign n3178 =  ( n2895 ) ? ( bv_8_88_n549 ) : ( n3177 ) ;
assign n3179 =  ( n2893 ) ? ( bv_8_207_n190 ) : ( n3178 ) ;
assign n3180 =  ( n2891 ) ? ( bv_8_208_n186 ) : ( n3179 ) ;
assign n3181 =  ( n2889 ) ? ( bv_8_239_n69 ) : ( n3180 ) ;
assign n3182 =  ( n2887 ) ? ( bv_8_170_n318 ) : ( n3181 ) ;
assign n3183 =  ( n2885 ) ? ( bv_8_251_n21 ) : ( n3182 ) ;
assign n3184 =  ( n2883 ) ? ( bv_8_67_n535 ) : ( n3183 ) ;
assign n3185 =  ( n2881 ) ? ( bv_8_77_n532 ) : ( n3184 ) ;
assign n3186 =  ( n2879 ) ? ( bv_8_51_n529 ) : ( n3185 ) ;
assign n3187 =  ( n2877 ) ? ( bv_8_133_n435 ) : ( n3186 ) ;
assign n3188 =  ( n2875 ) ? ( bv_8_69_n523 ) : ( n3187 ) ;
assign n3189 =  ( n2873 ) ? ( bv_8_249_n29 ) : ( n3188 ) ;
assign n3190 =  ( n2871 ) ? ( bv_8_2_n518 ) : ( n3189 ) ;
assign n3191 =  ( n2869 ) ? ( bv_8_127_n455 ) : ( n3190 ) ;
assign n3192 =  ( n2867 ) ? ( bv_8_80_n511 ) : ( n3191 ) ;
assign n3193 =  ( n2865 ) ? ( bv_8_60_n508 ) : ( n3192 ) ;
assign n3194 =  ( n2863 ) ? ( bv_8_159_n355 ) : ( n3193 ) ;
assign n3195 =  ( n2861 ) ? ( bv_8_168_n323 ) : ( n3194 ) ;
assign n3196 =  ( n2859 ) ? ( bv_8_81_n499 ) : ( n3195 ) ;
assign n3197 =  ( n2857 ) ? ( bv_8_163_n341 ) : ( n3196 ) ;
assign n3198 =  ( n2855 ) ? ( bv_8_64_n493 ) : ( n3197 ) ;
assign n3199 =  ( n2853 ) ? ( bv_8_143_n406 ) : ( n3198 ) ;
assign n3200 =  ( n2851 ) ? ( bv_8_146_n396 ) : ( n3199 ) ;
assign n3201 =  ( n2849 ) ? ( bv_8_157_n361 ) : ( n3200 ) ;
assign n3202 =  ( n2847 ) ? ( bv_8_56_n482 ) : ( n3201 ) ;
assign n3203 =  ( n2845 ) ? ( bv_8_245_n45 ) : ( n3202 ) ;
assign n3204 =  ( n2843 ) ? ( bv_8_188_n259 ) : ( n3203 ) ;
assign n3205 =  ( n2841 ) ? ( bv_8_182_n278 ) : ( n3204 ) ;
assign n3206 =  ( n2839 ) ? ( bv_8_218_n148 ) : ( n3205 ) ;
assign n3207 =  ( n2837 ) ? ( bv_8_33_n469 ) : ( n3206 ) ;
assign n3208 =  ( n2835 ) ? ( bv_8_16_n465 ) : ( n3207 ) ;
assign n3209 =  ( n2833 ) ? ( bv_8_255_n5 ) : ( n3208 ) ;
assign n3210 =  ( n2831 ) ? ( bv_8_243_n53 ) : ( n3209 ) ;
assign n3211 =  ( n2829 ) ? ( bv_8_210_n178 ) : ( n3210 ) ;
assign n3212 =  ( n2827 ) ? ( bv_8_205_n197 ) : ( n3211 ) ;
assign n3213 =  ( n2825 ) ? ( bv_8_12_n450 ) : ( n3212 ) ;
assign n3214 =  ( n2823 ) ? ( bv_8_19_n447 ) : ( n3213 ) ;
assign n3215 =  ( n2821 ) ? ( bv_8_236_n81 ) : ( n3214 ) ;
assign n3216 =  ( n2819 ) ? ( bv_8_95_n440 ) : ( n3215 ) ;
assign n3217 =  ( n2817 ) ? ( bv_8_151_n379 ) : ( n3216 ) ;
assign n3218 =  ( n2815 ) ? ( bv_8_68_n433 ) : ( n3217 ) ;
assign n3219 =  ( n2813 ) ? ( bv_8_23_n430 ) : ( n3218 ) ;
assign n3220 =  ( n2811 ) ? ( bv_8_196_n230 ) : ( n3219 ) ;
assign n3221 =  ( n2809 ) ? ( bv_8_167_n326 ) : ( n3220 ) ;
assign n3222 =  ( n2807 ) ? ( bv_8_126_n423 ) : ( n3221 ) ;
assign n3223 =  ( n2805 ) ? ( bv_8_61_n420 ) : ( n3222 ) ;
assign n3224 =  ( n2803 ) ? ( bv_8_100_n417 ) : ( n3223 ) ;
assign n3225 =  ( n2801 ) ? ( bv_8_93_n414 ) : ( n3224 ) ;
assign n3226 =  ( n2799 ) ? ( bv_8_25_n411 ) : ( n3225 ) ;
assign n3227 =  ( n2797 ) ? ( bv_8_115_n408 ) : ( n3226 ) ;
assign n3228 =  ( n2795 ) ? ( bv_8_96_n404 ) : ( n3227 ) ;
assign n3229 =  ( n2793 ) ? ( bv_8_129_n401 ) : ( n3228 ) ;
assign n3230 =  ( n2791 ) ? ( bv_8_79_n398 ) : ( n3229 ) ;
assign n3231 =  ( n2789 ) ? ( bv_8_220_n140 ) : ( n3230 ) ;
assign n3232 =  ( n2787 ) ? ( bv_8_34_n391 ) : ( n3231 ) ;
assign n3233 =  ( n2785 ) ? ( bv_8_42_n388 ) : ( n3232 ) ;
assign n3234 =  ( n2783 ) ? ( bv_8_144_n385 ) : ( n3233 ) ;
assign n3235 =  ( n2781 ) ? ( bv_8_136_n381 ) : ( n3234 ) ;
assign n3236 =  ( n2779 ) ? ( bv_8_70_n377 ) : ( n3235 ) ;
assign n3237 =  ( n2777 ) ? ( bv_8_238_n73 ) : ( n3236 ) ;
assign n3238 =  ( n2775 ) ? ( bv_8_184_n270 ) : ( n3237 ) ;
assign n3239 =  ( n2773 ) ? ( bv_8_20_n369 ) : ( n3238 ) ;
assign n3240 =  ( n2771 ) ? ( bv_8_222_n132 ) : ( n3239 ) ;
assign n3241 =  ( n2769 ) ? ( bv_8_94_n363 ) : ( n3240 ) ;
assign n3242 =  ( n2767 ) ? ( bv_8_11_n359 ) : ( n3241 ) ;
assign n3243 =  ( n2765 ) ? ( bv_8_219_n144 ) : ( n3242 ) ;
assign n3244 =  ( n2763 ) ? ( bv_8_224_n126 ) : ( n3243 ) ;
assign n3245 =  ( n2761 ) ? ( bv_8_50_n350 ) : ( n3244 ) ;
assign n3246 =  ( n2759 ) ? ( bv_8_58_n347 ) : ( n3245 ) ;
assign n3247 =  ( n2757 ) ? ( bv_8_10_n343 ) : ( n3246 ) ;
assign n3248 =  ( n2755 ) ? ( bv_8_73_n339 ) : ( n3247 ) ;
assign n3249 =  ( n2753 ) ? ( bv_8_6_n335 ) : ( n3248 ) ;
assign n3250 =  ( n2751 ) ? ( bv_8_36_n331 ) : ( n3249 ) ;
assign n3251 =  ( n2749 ) ? ( bv_8_92_n328 ) : ( n3250 ) ;
assign n3252 =  ( n2747 ) ? ( bv_8_194_n238 ) : ( n3251 ) ;
assign n3253 =  ( n2745 ) ? ( bv_8_211_n174 ) : ( n3252 ) ;
assign n3254 =  ( n2743 ) ? ( bv_8_172_n310 ) : ( n3253 ) ;
assign n3255 =  ( n2741 ) ? ( bv_8_98_n316 ) : ( n3254 ) ;
assign n3256 =  ( n2739 ) ? ( bv_8_145_n312 ) : ( n3255 ) ;
assign n3257 =  ( n2737 ) ? ( bv_8_149_n308 ) : ( n3256 ) ;
assign n3258 =  ( n2735 ) ? ( bv_8_228_n111 ) : ( n3257 ) ;
assign n3259 =  ( n2733 ) ? ( bv_8_121_n302 ) : ( n3258 ) ;
assign n3260 =  ( n2731 ) ? ( bv_8_231_n100 ) : ( n3259 ) ;
assign n3261 =  ( n2729 ) ? ( bv_8_200_n216 ) : ( n3260 ) ;
assign n3262 =  ( n2727 ) ? ( bv_8_55_n293 ) : ( n3261 ) ;
assign n3263 =  ( n2725 ) ? ( bv_8_109_n289 ) : ( n3262 ) ;
assign n3264 =  ( n2723 ) ? ( bv_8_141_n285 ) : ( n3263 ) ;
assign n3265 =  ( n2721 ) ? ( bv_8_213_n166 ) : ( n3264 ) ;
assign n3266 =  ( n2719 ) ? ( bv_8_78_n280 ) : ( n3265 ) ;
assign n3267 =  ( n2717 ) ? ( bv_8_169_n276 ) : ( n3266 ) ;
assign n3268 =  ( n2715 ) ? ( bv_8_108_n272 ) : ( n3267 ) ;
assign n3269 =  ( n2713 ) ? ( bv_8_86_n268 ) : ( n3268 ) ;
assign n3270 =  ( n2711 ) ? ( bv_8_244_n49 ) : ( n3269 ) ;
assign n3271 =  ( n2709 ) ? ( bv_8_234_n89 ) : ( n3270 ) ;
assign n3272 =  ( n2707 ) ? ( bv_8_101_n261 ) : ( n3271 ) ;
assign n3273 =  ( n2705 ) ? ( bv_8_122_n257 ) : ( n3272 ) ;
assign n3274 =  ( n2703 ) ? ( bv_8_174_n254 ) : ( n3273 ) ;
assign n3275 =  ( n2701 ) ? ( bv_8_8_n250 ) : ( n3274 ) ;
assign n3276 =  ( n2699 ) ? ( bv_8_186_n247 ) : ( n3275 ) ;
assign n3277 =  ( n2697 ) ? ( bv_8_120_n243 ) : ( n3276 ) ;
assign n3278 =  ( n2695 ) ? ( bv_8_37_n240 ) : ( n3277 ) ;
assign n3279 =  ( n2693 ) ? ( bv_8_46_n236 ) : ( n3278 ) ;
assign n3280 =  ( n2691 ) ? ( bv_8_28_n232 ) : ( n3279 ) ;
assign n3281 =  ( n2689 ) ? ( bv_8_166_n228 ) : ( n3280 ) ;
assign n3282 =  ( n2687 ) ? ( bv_8_180_n224 ) : ( n3281 ) ;
assign n3283 =  ( n2685 ) ? ( bv_8_198_n221 ) : ( n3282 ) ;
assign n3284 =  ( n2683 ) ? ( bv_8_232_n96 ) : ( n3283 ) ;
assign n3285 =  ( n2681 ) ? ( bv_8_221_n136 ) : ( n3284 ) ;
assign n3286 =  ( n2679 ) ? ( bv_8_116_n211 ) : ( n3285 ) ;
assign n3287 =  ( n2677 ) ? ( bv_8_31_n207 ) : ( n3286 ) ;
assign n3288 =  ( n2675 ) ? ( bv_8_75_n203 ) : ( n3287 ) ;
assign n3289 =  ( n2673 ) ? ( bv_8_189_n199 ) : ( n3288 ) ;
assign n3290 =  ( n2671 ) ? ( bv_8_139_n195 ) : ( n3289 ) ;
assign n3291 =  ( n2669 ) ? ( bv_8_138_n192 ) : ( n3290 ) ;
assign n3292 =  ( n2667 ) ? ( bv_8_112_n188 ) : ( n3291 ) ;
assign n3293 =  ( n2665 ) ? ( bv_8_62_n184 ) : ( n3292 ) ;
assign n3294 =  ( n2663 ) ? ( bv_8_181_n180 ) : ( n3293 ) ;
assign n3295 =  ( n2661 ) ? ( bv_8_102_n176 ) : ( n3294 ) ;
assign n3296 =  ( n2659 ) ? ( bv_8_72_n172 ) : ( n3295 ) ;
assign n3297 =  ( n2657 ) ? ( bv_8_3_n168 ) : ( n3296 ) ;
assign n3298 =  ( n2655 ) ? ( bv_8_246_n41 ) : ( n3297 ) ;
assign n3299 =  ( n2653 ) ? ( bv_8_14_n161 ) : ( n3298 ) ;
assign n3300 =  ( n2651 ) ? ( bv_8_97_n157 ) : ( n3299 ) ;
assign n3301 =  ( n2649 ) ? ( bv_8_53_n153 ) : ( n3300 ) ;
assign n3302 =  ( n2647 ) ? ( bv_8_87_n150 ) : ( n3301 ) ;
assign n3303 =  ( n2645 ) ? ( bv_8_185_n146 ) : ( n3302 ) ;
assign n3304 =  ( n2643 ) ? ( bv_8_134_n142 ) : ( n3303 ) ;
assign n3305 =  ( n2641 ) ? ( bv_8_193_n138 ) : ( n3304 ) ;
assign n3306 =  ( n2639 ) ? ( bv_8_29_n134 ) : ( n3305 ) ;
assign n3307 =  ( n2637 ) ? ( bv_8_158_n130 ) : ( n3306 ) ;
assign n3308 =  ( n2635 ) ? ( bv_8_225_n123 ) : ( n3307 ) ;
assign n3309 =  ( n2633 ) ? ( bv_8_248_n33 ) : ( n3308 ) ;
assign n3310 =  ( n2631 ) ? ( bv_8_152_n121 ) : ( n3309 ) ;
assign n3311 =  ( n2629 ) ? ( bv_8_17_n117 ) : ( n3310 ) ;
assign n3312 =  ( n2627 ) ? ( bv_8_105_n113 ) : ( n3311 ) ;
assign n3313 =  ( n2625 ) ? ( bv_8_217_n109 ) : ( n3312 ) ;
assign n3314 =  ( n2623 ) ? ( bv_8_142_n105 ) : ( n3313 ) ;
assign n3315 =  ( n2621 ) ? ( bv_8_148_n102 ) : ( n3314 ) ;
assign n3316 =  ( n2619 ) ? ( bv_8_155_n98 ) : ( n3315 ) ;
assign n3317 =  ( n2617 ) ? ( bv_8_30_n94 ) : ( n3316 ) ;
assign n3318 =  ( n2615 ) ? ( bv_8_135_n91 ) : ( n3317 ) ;
assign n3319 =  ( n2613 ) ? ( bv_8_233_n87 ) : ( n3318 ) ;
assign n3320 =  ( n2611 ) ? ( bv_8_206_n83 ) : ( n3319 ) ;
assign n3321 =  ( n2609 ) ? ( bv_8_85_n79 ) : ( n3320 ) ;
assign n3322 =  ( n2607 ) ? ( bv_8_40_n75 ) : ( n3321 ) ;
assign n3323 =  ( n2605 ) ? ( bv_8_223_n71 ) : ( n3322 ) ;
assign n3324 =  ( n2603 ) ? ( bv_8_140_n67 ) : ( n3323 ) ;
assign n3325 =  ( n2601 ) ? ( bv_8_161_n63 ) : ( n3324 ) ;
assign n3326 =  ( n2599 ) ? ( bv_8_137_n59 ) : ( n3325 ) ;
assign n3327 =  ( n2597 ) ? ( bv_8_13_n55 ) : ( n3326 ) ;
assign n3328 =  ( n2595 ) ? ( bv_8_191_n51 ) : ( n3327 ) ;
assign n3329 =  ( n2593 ) ? ( bv_8_230_n47 ) : ( n3328 ) ;
assign n3330 =  ( n2591 ) ? ( bv_8_66_n43 ) : ( n3329 ) ;
assign n3331 =  ( n2589 ) ? ( bv_8_104_n39 ) : ( n3330 ) ;
assign n3332 =  ( n2587 ) ? ( bv_8_65_n35 ) : ( n3331 ) ;
assign n3333 =  ( n2585 ) ? ( bv_8_153_n31 ) : ( n3332 ) ;
assign n3334 =  ( n2583 ) ? ( bv_8_45_n27 ) : ( n3333 ) ;
assign n3335 =  ( n2581 ) ? ( bv_8_15_n23 ) : ( n3334 ) ;
assign n3336 =  ( n2579 ) ? ( bv_8_176_n19 ) : ( n3335 ) ;
assign n3337 =  ( n2577 ) ? ( bv_8_84_n15 ) : ( n3336 ) ;
assign n3338 =  ( n2575 ) ? ( bv_8_187_n11 ) : ( n3337 ) ;
assign n3339 =  ( n2573 ) ? ( bv_8_22_n7 ) : ( n3338 ) ;
assign n3340 =  ( n2571 ) ^ ( n3339 )  ;
assign n3341 =  { ( n2570 ) , ( n3340 ) }  ;
assign n3342 = in[127:120] ;
assign n3343 =  ( n3342 ) ^ ( rcon )  ;
assign n3344 = in[95:88] ;
assign n3345 =  ( n3343 ) ^ ( n3344 )  ;
assign n3346 =  ( n3345 ) ^ ( n1027 )  ;
assign n3347 =  { ( n3341 ) , ( n3346 ) }  ;
assign n3348 = in[119:112] ;
assign n3349 = in[87:80] ;
assign n3350 =  ( n3348 ) ^ ( n3349 )  ;
assign n3351 =  ( n3350 ) ^ ( n1797 )  ;
assign n3352 =  { ( n3347 ) , ( n3351 ) }  ;
assign n3353 = in[111:104] ;
assign n3354 = in[79:72] ;
assign n3355 =  ( n3353 ) ^ ( n3354 )  ;
assign n3356 =  ( n3355 ) ^ ( n2568 )  ;
assign n3357 =  { ( n3352 ) , ( n3356 ) }  ;
assign n3358 = in[103:96] ;
assign n3359 = in[71:64] ;
assign n3360 =  ( n3358 ) ^ ( n3359 )  ;
assign n3361 =  ( n3360 ) ^ ( n3339 )  ;
assign n3362 =  { ( n3357 ) , ( n3361 ) }  ;
assign n3363 = in[127:120] ;
assign n3364 =  ( n3363 ) ^ ( rcon )  ;
assign n3365 = in[95:88] ;
assign n3366 =  ( n3364 ) ^ ( n3365 )  ;
assign n3367 = in[63:56] ;
assign n3368 =  ( n3366 ) ^ ( n3367 )  ;
assign n3369 =  ( n3368 ) ^ ( n1027 )  ;
assign n3370 =  { ( n3362 ) , ( n3369 ) }  ;
assign n3371 = in[119:112] ;
assign n3372 = in[87:80] ;
assign n3373 =  ( n3371 ) ^ ( n3372 )  ;
assign n3374 = in[55:48] ;
assign n3375 =  ( n3373 ) ^ ( n3374 )  ;
assign n3376 =  ( n3375 ) ^ ( n1797 )  ;
assign n3377 =  { ( n3370 ) , ( n3376 ) }  ;
assign n3378 = in[111:104] ;
assign n3379 = in[79:72] ;
assign n3380 =  ( n3378 ) ^ ( n3379 )  ;
assign n3381 = in[47:40] ;
assign n3382 =  ( n3380 ) ^ ( n3381 )  ;
assign n3383 =  ( n3382 ) ^ ( n2568 )  ;
assign n3384 =  { ( n3377 ) , ( n3383 ) }  ;
assign n3385 = in[103:96] ;
assign n3386 = in[71:64] ;
assign n3387 =  ( n3385 ) ^ ( n3386 )  ;
assign n3388 = in[39:32] ;
assign n3389 =  ( n3387 ) ^ ( n3388 )  ;
assign n3390 =  ( n3389 ) ^ ( n3339 )  ;
assign n3391 =  { ( n3384 ) , ( n3390 ) }  ;
assign n3392 = in[127:120] ;
assign n3393 =  ( n3392 ) ^ ( rcon )  ;
assign n3394 = in[95:88] ;
assign n3395 =  ( n3393 ) ^ ( n3394 )  ;
assign n3396 = in[63:56] ;
assign n3397 =  ( n3395 ) ^ ( n3396 )  ;
assign n3398 = in[31:24] ;
assign n3399 =  ( n3397 ) ^ ( n3398 )  ;
assign n3400 =  ( n3399 ) ^ ( n1027 )  ;
assign n3401 =  { ( n3391 ) , ( n3400 ) }  ;
assign n3402 = in[119:112] ;
assign n3403 = in[87:80] ;
assign n3404 =  ( n3402 ) ^ ( n3403 )  ;
assign n3405 = in[55:48] ;
assign n3406 =  ( n3404 ) ^ ( n3405 )  ;
assign n3407 = in[23:16] ;
assign n3408 =  ( n3406 ) ^ ( n3407 )  ;
assign n3409 =  ( n3408 ) ^ ( n1797 )  ;
assign n3410 =  { ( n3401 ) , ( n3409 ) }  ;
assign n3411 = in[111:104] ;
assign n3412 = in[79:72] ;
assign n3413 =  ( n3411 ) ^ ( n3412 )  ;
assign n3414 = in[47:40] ;
assign n3415 =  ( n3413 ) ^ ( n3414 )  ;
assign n3416 = in[15:8] ;
assign n3417 =  ( n3415 ) ^ ( n3416 )  ;
assign n3418 =  ( n3417 ) ^ ( n2568 )  ;
assign n3419 =  { ( n3410 ) , ( n3418 ) }  ;
assign n3420 = in[103:96] ;
assign n3421 = in[71:64] ;
assign n3422 =  ( n3420 ) ^ ( n3421 )  ;
assign n3423 = in[39:32] ;
assign n3424 =  ( n3422 ) ^ ( n3423 )  ;
assign n3425 = in[7:0] ;
assign n3426 =  ( n3424 ) ^ ( n3425 )  ;
assign n3427 =  ( n3426 ) ^ ( n3339 )  ;
assign n3428 =  { ( n3419 ) , ( n3427 ) }  ;
assign n3429 =  ( bv_128_0_n1 ) + ( n3428 )  ;
assign n3430 = in[127:120] ;
assign n3431 =  ( n3430 ) ^ ( rcon )  ;
assign n3432 = in[23:16] ;
assign n3433 =  ( n3432 ) == ( bv_8_255_n5 )  ;
assign n3434 = in[23:16] ;
assign n3435 =  ( n3434 ) == ( bv_8_254_n9 )  ;
assign n3436 = in[23:16] ;
assign n3437 =  ( n3436 ) == ( bv_8_253_n13 )  ;
assign n3438 = in[23:16] ;
assign n3439 =  ( n3438 ) == ( bv_8_252_n17 )  ;
assign n3440 = in[23:16] ;
assign n3441 =  ( n3440 ) == ( bv_8_251_n21 )  ;
assign n3442 = in[23:16] ;
assign n3443 =  ( n3442 ) == ( bv_8_250_n25 )  ;
assign n3444 = in[23:16] ;
assign n3445 =  ( n3444 ) == ( bv_8_249_n29 )  ;
assign n3446 = in[23:16] ;
assign n3447 =  ( n3446 ) == ( bv_8_248_n33 )  ;
assign n3448 = in[23:16] ;
assign n3449 =  ( n3448 ) == ( bv_8_247_n37 )  ;
assign n3450 = in[23:16] ;
assign n3451 =  ( n3450 ) == ( bv_8_246_n41 )  ;
assign n3452 = in[23:16] ;
assign n3453 =  ( n3452 ) == ( bv_8_245_n45 )  ;
assign n3454 = in[23:16] ;
assign n3455 =  ( n3454 ) == ( bv_8_244_n49 )  ;
assign n3456 = in[23:16] ;
assign n3457 =  ( n3456 ) == ( bv_8_243_n53 )  ;
assign n3458 = in[23:16] ;
assign n3459 =  ( n3458 ) == ( bv_8_242_n57 )  ;
assign n3460 = in[23:16] ;
assign n3461 =  ( n3460 ) == ( bv_8_241_n61 )  ;
assign n3462 = in[23:16] ;
assign n3463 =  ( n3462 ) == ( bv_8_240_n65 )  ;
assign n3464 = in[23:16] ;
assign n3465 =  ( n3464 ) == ( bv_8_239_n69 )  ;
assign n3466 = in[23:16] ;
assign n3467 =  ( n3466 ) == ( bv_8_238_n73 )  ;
assign n3468 = in[23:16] ;
assign n3469 =  ( n3468 ) == ( bv_8_237_n77 )  ;
assign n3470 = in[23:16] ;
assign n3471 =  ( n3470 ) == ( bv_8_236_n81 )  ;
assign n3472 = in[23:16] ;
assign n3473 =  ( n3472 ) == ( bv_8_235_n85 )  ;
assign n3474 = in[23:16] ;
assign n3475 =  ( n3474 ) == ( bv_8_234_n89 )  ;
assign n3476 = in[23:16] ;
assign n3477 =  ( n3476 ) == ( bv_8_233_n87 )  ;
assign n3478 = in[23:16] ;
assign n3479 =  ( n3478 ) == ( bv_8_232_n96 )  ;
assign n3480 = in[23:16] ;
assign n3481 =  ( n3480 ) == ( bv_8_231_n100 )  ;
assign n3482 = in[23:16] ;
assign n3483 =  ( n3482 ) == ( bv_8_230_n47 )  ;
assign n3484 = in[23:16] ;
assign n3485 =  ( n3484 ) == ( bv_8_229_n107 )  ;
assign n3486 = in[23:16] ;
assign n3487 =  ( n3486 ) == ( bv_8_228_n111 )  ;
assign n3488 = in[23:16] ;
assign n3489 =  ( n3488 ) == ( bv_8_227_n115 )  ;
assign n3490 = in[23:16] ;
assign n3491 =  ( n3490 ) == ( bv_8_226_n119 )  ;
assign n3492 = in[23:16] ;
assign n3493 =  ( n3492 ) == ( bv_8_225_n123 )  ;
assign n3494 = in[23:16] ;
assign n3495 =  ( n3494 ) == ( bv_8_224_n126 )  ;
assign n3496 = in[23:16] ;
assign n3497 =  ( n3496 ) == ( bv_8_223_n71 )  ;
assign n3498 = in[23:16] ;
assign n3499 =  ( n3498 ) == ( bv_8_222_n132 )  ;
assign n3500 = in[23:16] ;
assign n3501 =  ( n3500 ) == ( bv_8_221_n136 )  ;
assign n3502 = in[23:16] ;
assign n3503 =  ( n3502 ) == ( bv_8_220_n140 )  ;
assign n3504 = in[23:16] ;
assign n3505 =  ( n3504 ) == ( bv_8_219_n144 )  ;
assign n3506 = in[23:16] ;
assign n3507 =  ( n3506 ) == ( bv_8_218_n148 )  ;
assign n3508 = in[23:16] ;
assign n3509 =  ( n3508 ) == ( bv_8_217_n109 )  ;
assign n3510 = in[23:16] ;
assign n3511 =  ( n3510 ) == ( bv_8_216_n155 )  ;
assign n3512 = in[23:16] ;
assign n3513 =  ( n3512 ) == ( bv_8_215_n159 )  ;
assign n3514 = in[23:16] ;
assign n3515 =  ( n3514 ) == ( bv_8_214_n163 )  ;
assign n3516 = in[23:16] ;
assign n3517 =  ( n3516 ) == ( bv_8_213_n166 )  ;
assign n3518 = in[23:16] ;
assign n3519 =  ( n3518 ) == ( bv_8_212_n170 )  ;
assign n3520 = in[23:16] ;
assign n3521 =  ( n3520 ) == ( bv_8_211_n174 )  ;
assign n3522 = in[23:16] ;
assign n3523 =  ( n3522 ) == ( bv_8_210_n178 )  ;
assign n3524 = in[23:16] ;
assign n3525 =  ( n3524 ) == ( bv_8_209_n182 )  ;
assign n3526 = in[23:16] ;
assign n3527 =  ( n3526 ) == ( bv_8_208_n186 )  ;
assign n3528 = in[23:16] ;
assign n3529 =  ( n3528 ) == ( bv_8_207_n190 )  ;
assign n3530 = in[23:16] ;
assign n3531 =  ( n3530 ) == ( bv_8_206_n83 )  ;
assign n3532 = in[23:16] ;
assign n3533 =  ( n3532 ) == ( bv_8_205_n197 )  ;
assign n3534 = in[23:16] ;
assign n3535 =  ( n3534 ) == ( bv_8_204_n201 )  ;
assign n3536 = in[23:16] ;
assign n3537 =  ( n3536 ) == ( bv_8_203_n205 )  ;
assign n3538 = in[23:16] ;
assign n3539 =  ( n3538 ) == ( bv_8_202_n209 )  ;
assign n3540 = in[23:16] ;
assign n3541 =  ( n3540 ) == ( bv_8_201_n213 )  ;
assign n3542 = in[23:16] ;
assign n3543 =  ( n3542 ) == ( bv_8_200_n216 )  ;
assign n3544 = in[23:16] ;
assign n3545 =  ( n3544 ) == ( bv_8_199_n219 )  ;
assign n3546 = in[23:16] ;
assign n3547 =  ( n3546 ) == ( bv_8_198_n221 )  ;
assign n3548 = in[23:16] ;
assign n3549 =  ( n3548 ) == ( bv_8_197_n226 )  ;
assign n3550 = in[23:16] ;
assign n3551 =  ( n3550 ) == ( bv_8_196_n230 )  ;
assign n3552 = in[23:16] ;
assign n3553 =  ( n3552 ) == ( bv_8_195_n234 )  ;
assign n3554 = in[23:16] ;
assign n3555 =  ( n3554 ) == ( bv_8_194_n238 )  ;
assign n3556 = in[23:16] ;
assign n3557 =  ( n3556 ) == ( bv_8_193_n138 )  ;
assign n3558 = in[23:16] ;
assign n3559 =  ( n3558 ) == ( bv_8_192_n245 )  ;
assign n3560 = in[23:16] ;
assign n3561 =  ( n3560 ) == ( bv_8_191_n51 )  ;
assign n3562 = in[23:16] ;
assign n3563 =  ( n3562 ) == ( bv_8_190_n252 )  ;
assign n3564 = in[23:16] ;
assign n3565 =  ( n3564 ) == ( bv_8_189_n199 )  ;
assign n3566 = in[23:16] ;
assign n3567 =  ( n3566 ) == ( bv_8_188_n259 )  ;
assign n3568 = in[23:16] ;
assign n3569 =  ( n3568 ) == ( bv_8_187_n11 )  ;
assign n3570 = in[23:16] ;
assign n3571 =  ( n3570 ) == ( bv_8_186_n247 )  ;
assign n3572 = in[23:16] ;
assign n3573 =  ( n3572 ) == ( bv_8_185_n146 )  ;
assign n3574 = in[23:16] ;
assign n3575 =  ( n3574 ) == ( bv_8_184_n270 )  ;
assign n3576 = in[23:16] ;
assign n3577 =  ( n3576 ) == ( bv_8_183_n274 )  ;
assign n3578 = in[23:16] ;
assign n3579 =  ( n3578 ) == ( bv_8_182_n278 )  ;
assign n3580 = in[23:16] ;
assign n3581 =  ( n3580 ) == ( bv_8_181_n180 )  ;
assign n3582 = in[23:16] ;
assign n3583 =  ( n3582 ) == ( bv_8_180_n224 )  ;
assign n3584 = in[23:16] ;
assign n3585 =  ( n3584 ) == ( bv_8_179_n287 )  ;
assign n3586 = in[23:16] ;
assign n3587 =  ( n3586 ) == ( bv_8_178_n291 )  ;
assign n3588 = in[23:16] ;
assign n3589 =  ( n3588 ) == ( bv_8_177_n295 )  ;
assign n3590 = in[23:16] ;
assign n3591 =  ( n3590 ) == ( bv_8_176_n19 )  ;
assign n3592 = in[23:16] ;
assign n3593 =  ( n3592 ) == ( bv_8_175_n300 )  ;
assign n3594 = in[23:16] ;
assign n3595 =  ( n3594 ) == ( bv_8_174_n254 )  ;
assign n3596 = in[23:16] ;
assign n3597 =  ( n3596 ) == ( bv_8_173_n306 )  ;
assign n3598 = in[23:16] ;
assign n3599 =  ( n3598 ) == ( bv_8_172_n310 )  ;
assign n3600 = in[23:16] ;
assign n3601 =  ( n3600 ) == ( bv_8_171_n314 )  ;
assign n3602 = in[23:16] ;
assign n3603 =  ( n3602 ) == ( bv_8_170_n318 )  ;
assign n3604 = in[23:16] ;
assign n3605 =  ( n3604 ) == ( bv_8_169_n276 )  ;
assign n3606 = in[23:16] ;
assign n3607 =  ( n3606 ) == ( bv_8_168_n323 )  ;
assign n3608 = in[23:16] ;
assign n3609 =  ( n3608 ) == ( bv_8_167_n326 )  ;
assign n3610 = in[23:16] ;
assign n3611 =  ( n3610 ) == ( bv_8_166_n228 )  ;
assign n3612 = in[23:16] ;
assign n3613 =  ( n3612 ) == ( bv_8_165_n333 )  ;
assign n3614 = in[23:16] ;
assign n3615 =  ( n3614 ) == ( bv_8_164_n337 )  ;
assign n3616 = in[23:16] ;
assign n3617 =  ( n3616 ) == ( bv_8_163_n341 )  ;
assign n3618 = in[23:16] ;
assign n3619 =  ( n3618 ) == ( bv_8_162_n345 )  ;
assign n3620 = in[23:16] ;
assign n3621 =  ( n3620 ) == ( bv_8_161_n63 )  ;
assign n3622 = in[23:16] ;
assign n3623 =  ( n3622 ) == ( bv_8_160_n352 )  ;
assign n3624 = in[23:16] ;
assign n3625 =  ( n3624 ) == ( bv_8_159_n355 )  ;
assign n3626 = in[23:16] ;
assign n3627 =  ( n3626 ) == ( bv_8_158_n130 )  ;
assign n3628 = in[23:16] ;
assign n3629 =  ( n3628 ) == ( bv_8_157_n361 )  ;
assign n3630 = in[23:16] ;
assign n3631 =  ( n3630 ) == ( bv_8_156_n365 )  ;
assign n3632 = in[23:16] ;
assign n3633 =  ( n3632 ) == ( bv_8_155_n98 )  ;
assign n3634 = in[23:16] ;
assign n3635 =  ( n3634 ) == ( bv_8_154_n371 )  ;
assign n3636 = in[23:16] ;
assign n3637 =  ( n3636 ) == ( bv_8_153_n31 )  ;
assign n3638 = in[23:16] ;
assign n3639 =  ( n3638 ) == ( bv_8_152_n121 )  ;
assign n3640 = in[23:16] ;
assign n3641 =  ( n3640 ) == ( bv_8_151_n379 )  ;
assign n3642 = in[23:16] ;
assign n3643 =  ( n3642 ) == ( bv_8_150_n383 )  ;
assign n3644 = in[23:16] ;
assign n3645 =  ( n3644 ) == ( bv_8_149_n308 )  ;
assign n3646 = in[23:16] ;
assign n3647 =  ( n3646 ) == ( bv_8_148_n102 )  ;
assign n3648 = in[23:16] ;
assign n3649 =  ( n3648 ) == ( bv_8_147_n393 )  ;
assign n3650 = in[23:16] ;
assign n3651 =  ( n3650 ) == ( bv_8_146_n396 )  ;
assign n3652 = in[23:16] ;
assign n3653 =  ( n3652 ) == ( bv_8_145_n312 )  ;
assign n3654 = in[23:16] ;
assign n3655 =  ( n3654 ) == ( bv_8_144_n385 )  ;
assign n3656 = in[23:16] ;
assign n3657 =  ( n3656 ) == ( bv_8_143_n406 )  ;
assign n3658 = in[23:16] ;
assign n3659 =  ( n3658 ) == ( bv_8_142_n105 )  ;
assign n3660 = in[23:16] ;
assign n3661 =  ( n3660 ) == ( bv_8_141_n285 )  ;
assign n3662 = in[23:16] ;
assign n3663 =  ( n3662 ) == ( bv_8_140_n67 )  ;
assign n3664 = in[23:16] ;
assign n3665 =  ( n3664 ) == ( bv_8_139_n195 )  ;
assign n3666 = in[23:16] ;
assign n3667 =  ( n3666 ) == ( bv_8_138_n192 )  ;
assign n3668 = in[23:16] ;
assign n3669 =  ( n3668 ) == ( bv_8_137_n59 )  ;
assign n3670 = in[23:16] ;
assign n3671 =  ( n3670 ) == ( bv_8_136_n381 )  ;
assign n3672 = in[23:16] ;
assign n3673 =  ( n3672 ) == ( bv_8_135_n91 )  ;
assign n3674 = in[23:16] ;
assign n3675 =  ( n3674 ) == ( bv_8_134_n142 )  ;
assign n3676 = in[23:16] ;
assign n3677 =  ( n3676 ) == ( bv_8_133_n435 )  ;
assign n3678 = in[23:16] ;
assign n3679 =  ( n3678 ) == ( bv_8_132_n438 )  ;
assign n3680 = in[23:16] ;
assign n3681 =  ( n3680 ) == ( bv_8_131_n442 )  ;
assign n3682 = in[23:16] ;
assign n3683 =  ( n3682 ) == ( bv_8_130_n445 )  ;
assign n3684 = in[23:16] ;
assign n3685 =  ( n3684 ) == ( bv_8_129_n401 )  ;
assign n3686 = in[23:16] ;
assign n3687 =  ( n3686 ) == ( bv_8_128_n452 )  ;
assign n3688 = in[23:16] ;
assign n3689 =  ( n3688 ) == ( bv_8_127_n455 )  ;
assign n3690 = in[23:16] ;
assign n3691 =  ( n3690 ) == ( bv_8_126_n423 )  ;
assign n3692 = in[23:16] ;
assign n3693 =  ( n3692 ) == ( bv_8_125_n460 )  ;
assign n3694 = in[23:16] ;
assign n3695 =  ( n3694 ) == ( bv_8_124_n463 )  ;
assign n3696 = in[23:16] ;
assign n3697 =  ( n3696 ) == ( bv_8_123_n467 )  ;
assign n3698 = in[23:16] ;
assign n3699 =  ( n3698 ) == ( bv_8_122_n257 )  ;
assign n3700 = in[23:16] ;
assign n3701 =  ( n3700 ) == ( bv_8_121_n302 )  ;
assign n3702 = in[23:16] ;
assign n3703 =  ( n3702 ) == ( bv_8_120_n243 )  ;
assign n3704 = in[23:16] ;
assign n3705 =  ( n3704 ) == ( bv_8_119_n477 )  ;
assign n3706 = in[23:16] ;
assign n3707 =  ( n3706 ) == ( bv_8_118_n480 )  ;
assign n3708 = in[23:16] ;
assign n3709 =  ( n3708 ) == ( bv_8_117_n484 )  ;
assign n3710 = in[23:16] ;
assign n3711 =  ( n3710 ) == ( bv_8_116_n211 )  ;
assign n3712 = in[23:16] ;
assign n3713 =  ( n3712 ) == ( bv_8_115_n408 )  ;
assign n3714 = in[23:16] ;
assign n3715 =  ( n3714 ) == ( bv_8_114_n491 )  ;
assign n3716 = in[23:16] ;
assign n3717 =  ( n3716 ) == ( bv_8_113_n495 )  ;
assign n3718 = in[23:16] ;
assign n3719 =  ( n3718 ) == ( bv_8_112_n188 )  ;
assign n3720 = in[23:16] ;
assign n3721 =  ( n3720 ) == ( bv_8_111_n501 )  ;
assign n3722 = in[23:16] ;
assign n3723 =  ( n3722 ) == ( bv_8_110_n504 )  ;
assign n3724 = in[23:16] ;
assign n3725 =  ( n3724 ) == ( bv_8_109_n289 )  ;
assign n3726 = in[23:16] ;
assign n3727 =  ( n3726 ) == ( bv_8_108_n272 )  ;
assign n3728 = in[23:16] ;
assign n3729 =  ( n3728 ) == ( bv_8_107_n513 )  ;
assign n3730 = in[23:16] ;
assign n3731 =  ( n3730 ) == ( bv_8_106_n516 )  ;
assign n3732 = in[23:16] ;
assign n3733 =  ( n3732 ) == ( bv_8_105_n113 )  ;
assign n3734 = in[23:16] ;
assign n3735 =  ( n3734 ) == ( bv_8_104_n39 )  ;
assign n3736 = in[23:16] ;
assign n3737 =  ( n3736 ) == ( bv_8_103_n525 )  ;
assign n3738 = in[23:16] ;
assign n3739 =  ( n3738 ) == ( bv_8_102_n176 )  ;
assign n3740 = in[23:16] ;
assign n3741 =  ( n3740 ) == ( bv_8_101_n261 )  ;
assign n3742 = in[23:16] ;
assign n3743 =  ( n3742 ) == ( bv_8_100_n417 )  ;
assign n3744 = in[23:16] ;
assign n3745 =  ( n3744 ) == ( bv_8_99_n537 )  ;
assign n3746 = in[23:16] ;
assign n3747 =  ( n3746 ) == ( bv_8_98_n316 )  ;
assign n3748 = in[23:16] ;
assign n3749 =  ( n3748 ) == ( bv_8_97_n157 )  ;
assign n3750 = in[23:16] ;
assign n3751 =  ( n3750 ) == ( bv_8_96_n404 )  ;
assign n3752 = in[23:16] ;
assign n3753 =  ( n3752 ) == ( bv_8_95_n440 )  ;
assign n3754 = in[23:16] ;
assign n3755 =  ( n3754 ) == ( bv_8_94_n363 )  ;
assign n3756 = in[23:16] ;
assign n3757 =  ( n3756 ) == ( bv_8_93_n414 )  ;
assign n3758 = in[23:16] ;
assign n3759 =  ( n3758 ) == ( bv_8_92_n328 )  ;
assign n3760 = in[23:16] ;
assign n3761 =  ( n3760 ) == ( bv_8_91_n557 )  ;
assign n3762 = in[23:16] ;
assign n3763 =  ( n3762 ) == ( bv_8_90_n561 )  ;
assign n3764 = in[23:16] ;
assign n3765 =  ( n3764 ) == ( bv_8_89_n564 )  ;
assign n3766 = in[23:16] ;
assign n3767 =  ( n3766 ) == ( bv_8_88_n549 )  ;
assign n3768 = in[23:16] ;
assign n3769 =  ( n3768 ) == ( bv_8_87_n150 )  ;
assign n3770 = in[23:16] ;
assign n3771 =  ( n3770 ) == ( bv_8_86_n268 )  ;
assign n3772 = in[23:16] ;
assign n3773 =  ( n3772 ) == ( bv_8_85_n79 )  ;
assign n3774 = in[23:16] ;
assign n3775 =  ( n3774 ) == ( bv_8_84_n15 )  ;
assign n3776 = in[23:16] ;
assign n3777 =  ( n3776 ) == ( bv_8_83_n578 )  ;
assign n3778 = in[23:16] ;
assign n3779 =  ( n3778 ) == ( bv_8_82_n581 )  ;
assign n3780 = in[23:16] ;
assign n3781 =  ( n3780 ) == ( bv_8_81_n499 )  ;
assign n3782 = in[23:16] ;
assign n3783 =  ( n3782 ) == ( bv_8_80_n511 )  ;
assign n3784 = in[23:16] ;
assign n3785 =  ( n3784 ) == ( bv_8_79_n398 )  ;
assign n3786 = in[23:16] ;
assign n3787 =  ( n3786 ) == ( bv_8_78_n280 )  ;
assign n3788 = in[23:16] ;
assign n3789 =  ( n3788 ) == ( bv_8_77_n532 )  ;
assign n3790 = in[23:16] ;
assign n3791 =  ( n3790 ) == ( bv_8_76_n552 )  ;
assign n3792 = in[23:16] ;
assign n3793 =  ( n3792 ) == ( bv_8_75_n203 )  ;
assign n3794 = in[23:16] ;
assign n3795 =  ( n3794 ) == ( bv_8_74_n555 )  ;
assign n3796 = in[23:16] ;
assign n3797 =  ( n3796 ) == ( bv_8_73_n339 )  ;
assign n3798 = in[23:16] ;
assign n3799 =  ( n3798 ) == ( bv_8_72_n172 )  ;
assign n3800 = in[23:16] ;
assign n3801 =  ( n3800 ) == ( bv_8_71_n608 )  ;
assign n3802 = in[23:16] ;
assign n3803 =  ( n3802 ) == ( bv_8_70_n377 )  ;
assign n3804 = in[23:16] ;
assign n3805 =  ( n3804 ) == ( bv_8_69_n523 )  ;
assign n3806 = in[23:16] ;
assign n3807 =  ( n3806 ) == ( bv_8_68_n433 )  ;
assign n3808 = in[23:16] ;
assign n3809 =  ( n3808 ) == ( bv_8_67_n535 )  ;
assign n3810 = in[23:16] ;
assign n3811 =  ( n3810 ) == ( bv_8_66_n43 )  ;
assign n3812 = in[23:16] ;
assign n3813 =  ( n3812 ) == ( bv_8_65_n35 )  ;
assign n3814 = in[23:16] ;
assign n3815 =  ( n3814 ) == ( bv_8_64_n493 )  ;
assign n3816 = in[23:16] ;
assign n3817 =  ( n3816 ) == ( bv_8_63_n629 )  ;
assign n3818 = in[23:16] ;
assign n3819 =  ( n3818 ) == ( bv_8_62_n184 )  ;
assign n3820 = in[23:16] ;
assign n3821 =  ( n3820 ) == ( bv_8_61_n420 )  ;
assign n3822 = in[23:16] ;
assign n3823 =  ( n3822 ) == ( bv_8_60_n508 )  ;
assign n3824 = in[23:16] ;
assign n3825 =  ( n3824 ) == ( bv_8_59_n604 )  ;
assign n3826 = in[23:16] ;
assign n3827 =  ( n3826 ) == ( bv_8_58_n347 )  ;
assign n3828 = in[23:16] ;
assign n3829 =  ( n3828 ) == ( bv_8_57_n559 )  ;
assign n3830 = in[23:16] ;
assign n3831 =  ( n3830 ) == ( bv_8_56_n482 )  ;
assign n3832 = in[23:16] ;
assign n3833 =  ( n3832 ) == ( bv_8_55_n293 )  ;
assign n3834 = in[23:16] ;
assign n3835 =  ( n3834 ) == ( bv_8_54_n651 )  ;
assign n3836 = in[23:16] ;
assign n3837 =  ( n3836 ) == ( bv_8_53_n153 )  ;
assign n3838 = in[23:16] ;
assign n3839 =  ( n3838 ) == ( bv_8_52_n657 )  ;
assign n3840 = in[23:16] ;
assign n3841 =  ( n3840 ) == ( bv_8_51_n529 )  ;
assign n3842 = in[23:16] ;
assign n3843 =  ( n3842 ) == ( bv_8_50_n350 )  ;
assign n3844 = in[23:16] ;
assign n3845 =  ( n3844 ) == ( bv_8_49_n666 )  ;
assign n3846 = in[23:16] ;
assign n3847 =  ( n3846 ) == ( bv_8_48_n669 )  ;
assign n3848 = in[23:16] ;
assign n3849 =  ( n3848 ) == ( bv_8_47_n592 )  ;
assign n3850 = in[23:16] ;
assign n3851 =  ( n3850 ) == ( bv_8_46_n236 )  ;
assign n3852 = in[23:16] ;
assign n3853 =  ( n3852 ) == ( bv_8_45_n27 )  ;
assign n3854 = in[23:16] ;
assign n3855 =  ( n3854 ) == ( bv_8_44_n622 )  ;
assign n3856 = in[23:16] ;
assign n3857 =  ( n3856 ) == ( bv_8_43_n682 )  ;
assign n3858 = in[23:16] ;
assign n3859 =  ( n3858 ) == ( bv_8_42_n388 )  ;
assign n3860 = in[23:16] ;
assign n3861 =  ( n3860 ) == ( bv_8_41_n597 )  ;
assign n3862 = in[23:16] ;
assign n3863 =  ( n3862 ) == ( bv_8_40_n75 )  ;
assign n3864 = in[23:16] ;
assign n3865 =  ( n3864 ) == ( bv_8_39_n635 )  ;
assign n3866 = in[23:16] ;
assign n3867 =  ( n3866 ) == ( bv_8_38_n693 )  ;
assign n3868 = in[23:16] ;
assign n3869 =  ( n3868 ) == ( bv_8_37_n240 )  ;
assign n3870 = in[23:16] ;
assign n3871 =  ( n3870 ) == ( bv_8_36_n331 )  ;
assign n3872 = in[23:16] ;
assign n3873 =  ( n3872 ) == ( bv_8_35_n664 )  ;
assign n3874 = in[23:16] ;
assign n3875 =  ( n3874 ) == ( bv_8_34_n391 )  ;
assign n3876 = in[23:16] ;
assign n3877 =  ( n3876 ) == ( bv_8_33_n469 )  ;
assign n3878 = in[23:16] ;
assign n3879 =  ( n3878 ) == ( bv_8_32_n576 )  ;
assign n3880 = in[23:16] ;
assign n3881 =  ( n3880 ) == ( bv_8_31_n207 )  ;
assign n3882 = in[23:16] ;
assign n3883 =  ( n3882 ) == ( bv_8_30_n94 )  ;
assign n3884 = in[23:16] ;
assign n3885 =  ( n3884 ) == ( bv_8_29_n134 )  ;
assign n3886 = in[23:16] ;
assign n3887 =  ( n3886 ) == ( bv_8_28_n232 )  ;
assign n3888 = in[23:16] ;
assign n3889 =  ( n3888 ) == ( bv_8_27_n616 )  ;
assign n3890 = in[23:16] ;
assign n3891 =  ( n3890 ) == ( bv_8_26_n619 )  ;
assign n3892 = in[23:16] ;
assign n3893 =  ( n3892 ) == ( bv_8_25_n411 )  ;
assign n3894 = in[23:16] ;
assign n3895 =  ( n3894 ) == ( bv_8_24_n659 )  ;
assign n3896 = in[23:16] ;
assign n3897 =  ( n3896 ) == ( bv_8_23_n430 )  ;
assign n3898 = in[23:16] ;
assign n3899 =  ( n3898 ) == ( bv_8_22_n7 )  ;
assign n3900 = in[23:16] ;
assign n3901 =  ( n3900 ) == ( bv_8_21_n674 )  ;
assign n3902 = in[23:16] ;
assign n3903 =  ( n3902 ) == ( bv_8_20_n369 )  ;
assign n3904 = in[23:16] ;
assign n3905 =  ( n3904 ) == ( bv_8_19_n447 )  ;
assign n3906 = in[23:16] ;
assign n3907 =  ( n3906 ) == ( bv_8_18_n644 )  ;
assign n3908 = in[23:16] ;
assign n3909 =  ( n3908 ) == ( bv_8_17_n117 )  ;
assign n3910 = in[23:16] ;
assign n3911 =  ( n3910 ) == ( bv_8_16_n465 )  ;
assign n3912 = in[23:16] ;
assign n3913 =  ( n3912 ) == ( bv_8_15_n23 )  ;
assign n3914 = in[23:16] ;
assign n3915 =  ( n3914 ) == ( bv_8_14_n161 )  ;
assign n3916 = in[23:16] ;
assign n3917 =  ( n3916 ) == ( bv_8_13_n55 )  ;
assign n3918 = in[23:16] ;
assign n3919 =  ( n3918 ) == ( bv_8_12_n450 )  ;
assign n3920 = in[23:16] ;
assign n3921 =  ( n3920 ) == ( bv_8_11_n359 )  ;
assign n3922 = in[23:16] ;
assign n3923 =  ( n3922 ) == ( bv_8_10_n343 )  ;
assign n3924 = in[23:16] ;
assign n3925 =  ( n3924 ) == ( bv_8_9_n627 )  ;
assign n3926 = in[23:16] ;
assign n3927 =  ( n3926 ) == ( bv_8_8_n250 )  ;
assign n3928 = in[23:16] ;
assign n3929 =  ( n3928 ) == ( bv_8_7_n647 )  ;
assign n3930 = in[23:16] ;
assign n3931 =  ( n3930 ) == ( bv_8_6_n335 )  ;
assign n3932 = in[23:16] ;
assign n3933 =  ( n3932 ) == ( bv_8_5_n653 )  ;
assign n3934 = in[23:16] ;
assign n3935 =  ( n3934 ) == ( bv_8_4_n671 )  ;
assign n3936 = in[23:16] ;
assign n3937 =  ( n3936 ) == ( bv_8_3_n168 )  ;
assign n3938 = in[23:16] ;
assign n3939 =  ( n3938 ) == ( bv_8_2_n518 )  ;
assign n3940 = in[23:16] ;
assign n3941 =  ( n3940 ) == ( bv_8_1_n753 )  ;
assign n3942 = in[23:16] ;
assign n3943 =  ( n3942 ) == ( bv_8_0_n583 )  ;
assign n3944 =  ( n3943 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n3945 =  ( n3941 ) ? ( bv_8_124_n463 ) : ( n3944 ) ;
assign n3946 =  ( n3939 ) ? ( bv_8_119_n477 ) : ( n3945 ) ;
assign n3947 =  ( n3937 ) ? ( bv_8_123_n467 ) : ( n3946 ) ;
assign n3948 =  ( n3935 ) ? ( bv_8_242_n57 ) : ( n3947 ) ;
assign n3949 =  ( n3933 ) ? ( bv_8_107_n513 ) : ( n3948 ) ;
assign n3950 =  ( n3931 ) ? ( bv_8_111_n501 ) : ( n3949 ) ;
assign n3951 =  ( n3929 ) ? ( bv_8_197_n226 ) : ( n3950 ) ;
assign n3952 =  ( n3927 ) ? ( bv_8_48_n669 ) : ( n3951 ) ;
assign n3953 =  ( n3925 ) ? ( bv_8_1_n753 ) : ( n3952 ) ;
assign n3954 =  ( n3923 ) ? ( bv_8_103_n525 ) : ( n3953 ) ;
assign n3955 =  ( n3921 ) ? ( bv_8_43_n682 ) : ( n3954 ) ;
assign n3956 =  ( n3919 ) ? ( bv_8_254_n9 ) : ( n3955 ) ;
assign n3957 =  ( n3917 ) ? ( bv_8_215_n159 ) : ( n3956 ) ;
assign n3958 =  ( n3915 ) ? ( bv_8_171_n314 ) : ( n3957 ) ;
assign n3959 =  ( n3913 ) ? ( bv_8_118_n480 ) : ( n3958 ) ;
assign n3960 =  ( n3911 ) ? ( bv_8_202_n209 ) : ( n3959 ) ;
assign n3961 =  ( n3909 ) ? ( bv_8_130_n445 ) : ( n3960 ) ;
assign n3962 =  ( n3907 ) ? ( bv_8_201_n213 ) : ( n3961 ) ;
assign n3963 =  ( n3905 ) ? ( bv_8_125_n460 ) : ( n3962 ) ;
assign n3964 =  ( n3903 ) ? ( bv_8_250_n25 ) : ( n3963 ) ;
assign n3965 =  ( n3901 ) ? ( bv_8_89_n564 ) : ( n3964 ) ;
assign n3966 =  ( n3899 ) ? ( bv_8_71_n608 ) : ( n3965 ) ;
assign n3967 =  ( n3897 ) ? ( bv_8_240_n65 ) : ( n3966 ) ;
assign n3968 =  ( n3895 ) ? ( bv_8_173_n306 ) : ( n3967 ) ;
assign n3969 =  ( n3893 ) ? ( bv_8_212_n170 ) : ( n3968 ) ;
assign n3970 =  ( n3891 ) ? ( bv_8_162_n345 ) : ( n3969 ) ;
assign n3971 =  ( n3889 ) ? ( bv_8_175_n300 ) : ( n3970 ) ;
assign n3972 =  ( n3887 ) ? ( bv_8_156_n365 ) : ( n3971 ) ;
assign n3973 =  ( n3885 ) ? ( bv_8_164_n337 ) : ( n3972 ) ;
assign n3974 =  ( n3883 ) ? ( bv_8_114_n491 ) : ( n3973 ) ;
assign n3975 =  ( n3881 ) ? ( bv_8_192_n245 ) : ( n3974 ) ;
assign n3976 =  ( n3879 ) ? ( bv_8_183_n274 ) : ( n3975 ) ;
assign n3977 =  ( n3877 ) ? ( bv_8_253_n13 ) : ( n3976 ) ;
assign n3978 =  ( n3875 ) ? ( bv_8_147_n393 ) : ( n3977 ) ;
assign n3979 =  ( n3873 ) ? ( bv_8_38_n693 ) : ( n3978 ) ;
assign n3980 =  ( n3871 ) ? ( bv_8_54_n651 ) : ( n3979 ) ;
assign n3981 =  ( n3869 ) ? ( bv_8_63_n629 ) : ( n3980 ) ;
assign n3982 =  ( n3867 ) ? ( bv_8_247_n37 ) : ( n3981 ) ;
assign n3983 =  ( n3865 ) ? ( bv_8_204_n201 ) : ( n3982 ) ;
assign n3984 =  ( n3863 ) ? ( bv_8_52_n657 ) : ( n3983 ) ;
assign n3985 =  ( n3861 ) ? ( bv_8_165_n333 ) : ( n3984 ) ;
assign n3986 =  ( n3859 ) ? ( bv_8_229_n107 ) : ( n3985 ) ;
assign n3987 =  ( n3857 ) ? ( bv_8_241_n61 ) : ( n3986 ) ;
assign n3988 =  ( n3855 ) ? ( bv_8_113_n495 ) : ( n3987 ) ;
assign n3989 =  ( n3853 ) ? ( bv_8_216_n155 ) : ( n3988 ) ;
assign n3990 =  ( n3851 ) ? ( bv_8_49_n666 ) : ( n3989 ) ;
assign n3991 =  ( n3849 ) ? ( bv_8_21_n674 ) : ( n3990 ) ;
assign n3992 =  ( n3847 ) ? ( bv_8_4_n671 ) : ( n3991 ) ;
assign n3993 =  ( n3845 ) ? ( bv_8_199_n219 ) : ( n3992 ) ;
assign n3994 =  ( n3843 ) ? ( bv_8_35_n664 ) : ( n3993 ) ;
assign n3995 =  ( n3841 ) ? ( bv_8_195_n234 ) : ( n3994 ) ;
assign n3996 =  ( n3839 ) ? ( bv_8_24_n659 ) : ( n3995 ) ;
assign n3997 =  ( n3837 ) ? ( bv_8_150_n383 ) : ( n3996 ) ;
assign n3998 =  ( n3835 ) ? ( bv_8_5_n653 ) : ( n3997 ) ;
assign n3999 =  ( n3833 ) ? ( bv_8_154_n371 ) : ( n3998 ) ;
assign n4000 =  ( n3831 ) ? ( bv_8_7_n647 ) : ( n3999 ) ;
assign n4001 =  ( n3829 ) ? ( bv_8_18_n644 ) : ( n4000 ) ;
assign n4002 =  ( n3827 ) ? ( bv_8_128_n452 ) : ( n4001 ) ;
assign n4003 =  ( n3825 ) ? ( bv_8_226_n119 ) : ( n4002 ) ;
assign n4004 =  ( n3823 ) ? ( bv_8_235_n85 ) : ( n4003 ) ;
assign n4005 =  ( n3821 ) ? ( bv_8_39_n635 ) : ( n4004 ) ;
assign n4006 =  ( n3819 ) ? ( bv_8_178_n291 ) : ( n4005 ) ;
assign n4007 =  ( n3817 ) ? ( bv_8_117_n484 ) : ( n4006 ) ;
assign n4008 =  ( n3815 ) ? ( bv_8_9_n627 ) : ( n4007 ) ;
assign n4009 =  ( n3813 ) ? ( bv_8_131_n442 ) : ( n4008 ) ;
assign n4010 =  ( n3811 ) ? ( bv_8_44_n622 ) : ( n4009 ) ;
assign n4011 =  ( n3809 ) ? ( bv_8_26_n619 ) : ( n4010 ) ;
assign n4012 =  ( n3807 ) ? ( bv_8_27_n616 ) : ( n4011 ) ;
assign n4013 =  ( n3805 ) ? ( bv_8_110_n504 ) : ( n4012 ) ;
assign n4014 =  ( n3803 ) ? ( bv_8_90_n561 ) : ( n4013 ) ;
assign n4015 =  ( n3801 ) ? ( bv_8_160_n352 ) : ( n4014 ) ;
assign n4016 =  ( n3799 ) ? ( bv_8_82_n581 ) : ( n4015 ) ;
assign n4017 =  ( n3797 ) ? ( bv_8_59_n604 ) : ( n4016 ) ;
assign n4018 =  ( n3795 ) ? ( bv_8_214_n163 ) : ( n4017 ) ;
assign n4019 =  ( n3793 ) ? ( bv_8_179_n287 ) : ( n4018 ) ;
assign n4020 =  ( n3791 ) ? ( bv_8_41_n597 ) : ( n4019 ) ;
assign n4021 =  ( n3789 ) ? ( bv_8_227_n115 ) : ( n4020 ) ;
assign n4022 =  ( n3787 ) ? ( bv_8_47_n592 ) : ( n4021 ) ;
assign n4023 =  ( n3785 ) ? ( bv_8_132_n438 ) : ( n4022 ) ;
assign n4024 =  ( n3783 ) ? ( bv_8_83_n578 ) : ( n4023 ) ;
assign n4025 =  ( n3781 ) ? ( bv_8_209_n182 ) : ( n4024 ) ;
assign n4026 =  ( n3779 ) ? ( bv_8_0_n583 ) : ( n4025 ) ;
assign n4027 =  ( n3777 ) ? ( bv_8_237_n77 ) : ( n4026 ) ;
assign n4028 =  ( n3775 ) ? ( bv_8_32_n576 ) : ( n4027 ) ;
assign n4029 =  ( n3773 ) ? ( bv_8_252_n17 ) : ( n4028 ) ;
assign n4030 =  ( n3771 ) ? ( bv_8_177_n295 ) : ( n4029 ) ;
assign n4031 =  ( n3769 ) ? ( bv_8_91_n557 ) : ( n4030 ) ;
assign n4032 =  ( n3767 ) ? ( bv_8_106_n516 ) : ( n4031 ) ;
assign n4033 =  ( n3765 ) ? ( bv_8_203_n205 ) : ( n4032 ) ;
assign n4034 =  ( n3763 ) ? ( bv_8_190_n252 ) : ( n4033 ) ;
assign n4035 =  ( n3761 ) ? ( bv_8_57_n559 ) : ( n4034 ) ;
assign n4036 =  ( n3759 ) ? ( bv_8_74_n555 ) : ( n4035 ) ;
assign n4037 =  ( n3757 ) ? ( bv_8_76_n552 ) : ( n4036 ) ;
assign n4038 =  ( n3755 ) ? ( bv_8_88_n549 ) : ( n4037 ) ;
assign n4039 =  ( n3753 ) ? ( bv_8_207_n190 ) : ( n4038 ) ;
assign n4040 =  ( n3751 ) ? ( bv_8_208_n186 ) : ( n4039 ) ;
assign n4041 =  ( n3749 ) ? ( bv_8_239_n69 ) : ( n4040 ) ;
assign n4042 =  ( n3747 ) ? ( bv_8_170_n318 ) : ( n4041 ) ;
assign n4043 =  ( n3745 ) ? ( bv_8_251_n21 ) : ( n4042 ) ;
assign n4044 =  ( n3743 ) ? ( bv_8_67_n535 ) : ( n4043 ) ;
assign n4045 =  ( n3741 ) ? ( bv_8_77_n532 ) : ( n4044 ) ;
assign n4046 =  ( n3739 ) ? ( bv_8_51_n529 ) : ( n4045 ) ;
assign n4047 =  ( n3737 ) ? ( bv_8_133_n435 ) : ( n4046 ) ;
assign n4048 =  ( n3735 ) ? ( bv_8_69_n523 ) : ( n4047 ) ;
assign n4049 =  ( n3733 ) ? ( bv_8_249_n29 ) : ( n4048 ) ;
assign n4050 =  ( n3731 ) ? ( bv_8_2_n518 ) : ( n4049 ) ;
assign n4051 =  ( n3729 ) ? ( bv_8_127_n455 ) : ( n4050 ) ;
assign n4052 =  ( n3727 ) ? ( bv_8_80_n511 ) : ( n4051 ) ;
assign n4053 =  ( n3725 ) ? ( bv_8_60_n508 ) : ( n4052 ) ;
assign n4054 =  ( n3723 ) ? ( bv_8_159_n355 ) : ( n4053 ) ;
assign n4055 =  ( n3721 ) ? ( bv_8_168_n323 ) : ( n4054 ) ;
assign n4056 =  ( n3719 ) ? ( bv_8_81_n499 ) : ( n4055 ) ;
assign n4057 =  ( n3717 ) ? ( bv_8_163_n341 ) : ( n4056 ) ;
assign n4058 =  ( n3715 ) ? ( bv_8_64_n493 ) : ( n4057 ) ;
assign n4059 =  ( n3713 ) ? ( bv_8_143_n406 ) : ( n4058 ) ;
assign n4060 =  ( n3711 ) ? ( bv_8_146_n396 ) : ( n4059 ) ;
assign n4061 =  ( n3709 ) ? ( bv_8_157_n361 ) : ( n4060 ) ;
assign n4062 =  ( n3707 ) ? ( bv_8_56_n482 ) : ( n4061 ) ;
assign n4063 =  ( n3705 ) ? ( bv_8_245_n45 ) : ( n4062 ) ;
assign n4064 =  ( n3703 ) ? ( bv_8_188_n259 ) : ( n4063 ) ;
assign n4065 =  ( n3701 ) ? ( bv_8_182_n278 ) : ( n4064 ) ;
assign n4066 =  ( n3699 ) ? ( bv_8_218_n148 ) : ( n4065 ) ;
assign n4067 =  ( n3697 ) ? ( bv_8_33_n469 ) : ( n4066 ) ;
assign n4068 =  ( n3695 ) ? ( bv_8_16_n465 ) : ( n4067 ) ;
assign n4069 =  ( n3693 ) ? ( bv_8_255_n5 ) : ( n4068 ) ;
assign n4070 =  ( n3691 ) ? ( bv_8_243_n53 ) : ( n4069 ) ;
assign n4071 =  ( n3689 ) ? ( bv_8_210_n178 ) : ( n4070 ) ;
assign n4072 =  ( n3687 ) ? ( bv_8_205_n197 ) : ( n4071 ) ;
assign n4073 =  ( n3685 ) ? ( bv_8_12_n450 ) : ( n4072 ) ;
assign n4074 =  ( n3683 ) ? ( bv_8_19_n447 ) : ( n4073 ) ;
assign n4075 =  ( n3681 ) ? ( bv_8_236_n81 ) : ( n4074 ) ;
assign n4076 =  ( n3679 ) ? ( bv_8_95_n440 ) : ( n4075 ) ;
assign n4077 =  ( n3677 ) ? ( bv_8_151_n379 ) : ( n4076 ) ;
assign n4078 =  ( n3675 ) ? ( bv_8_68_n433 ) : ( n4077 ) ;
assign n4079 =  ( n3673 ) ? ( bv_8_23_n430 ) : ( n4078 ) ;
assign n4080 =  ( n3671 ) ? ( bv_8_196_n230 ) : ( n4079 ) ;
assign n4081 =  ( n3669 ) ? ( bv_8_167_n326 ) : ( n4080 ) ;
assign n4082 =  ( n3667 ) ? ( bv_8_126_n423 ) : ( n4081 ) ;
assign n4083 =  ( n3665 ) ? ( bv_8_61_n420 ) : ( n4082 ) ;
assign n4084 =  ( n3663 ) ? ( bv_8_100_n417 ) : ( n4083 ) ;
assign n4085 =  ( n3661 ) ? ( bv_8_93_n414 ) : ( n4084 ) ;
assign n4086 =  ( n3659 ) ? ( bv_8_25_n411 ) : ( n4085 ) ;
assign n4087 =  ( n3657 ) ? ( bv_8_115_n408 ) : ( n4086 ) ;
assign n4088 =  ( n3655 ) ? ( bv_8_96_n404 ) : ( n4087 ) ;
assign n4089 =  ( n3653 ) ? ( bv_8_129_n401 ) : ( n4088 ) ;
assign n4090 =  ( n3651 ) ? ( bv_8_79_n398 ) : ( n4089 ) ;
assign n4091 =  ( n3649 ) ? ( bv_8_220_n140 ) : ( n4090 ) ;
assign n4092 =  ( n3647 ) ? ( bv_8_34_n391 ) : ( n4091 ) ;
assign n4093 =  ( n3645 ) ? ( bv_8_42_n388 ) : ( n4092 ) ;
assign n4094 =  ( n3643 ) ? ( bv_8_144_n385 ) : ( n4093 ) ;
assign n4095 =  ( n3641 ) ? ( bv_8_136_n381 ) : ( n4094 ) ;
assign n4096 =  ( n3639 ) ? ( bv_8_70_n377 ) : ( n4095 ) ;
assign n4097 =  ( n3637 ) ? ( bv_8_238_n73 ) : ( n4096 ) ;
assign n4098 =  ( n3635 ) ? ( bv_8_184_n270 ) : ( n4097 ) ;
assign n4099 =  ( n3633 ) ? ( bv_8_20_n369 ) : ( n4098 ) ;
assign n4100 =  ( n3631 ) ? ( bv_8_222_n132 ) : ( n4099 ) ;
assign n4101 =  ( n3629 ) ? ( bv_8_94_n363 ) : ( n4100 ) ;
assign n4102 =  ( n3627 ) ? ( bv_8_11_n359 ) : ( n4101 ) ;
assign n4103 =  ( n3625 ) ? ( bv_8_219_n144 ) : ( n4102 ) ;
assign n4104 =  ( n3623 ) ? ( bv_8_224_n126 ) : ( n4103 ) ;
assign n4105 =  ( n3621 ) ? ( bv_8_50_n350 ) : ( n4104 ) ;
assign n4106 =  ( n3619 ) ? ( bv_8_58_n347 ) : ( n4105 ) ;
assign n4107 =  ( n3617 ) ? ( bv_8_10_n343 ) : ( n4106 ) ;
assign n4108 =  ( n3615 ) ? ( bv_8_73_n339 ) : ( n4107 ) ;
assign n4109 =  ( n3613 ) ? ( bv_8_6_n335 ) : ( n4108 ) ;
assign n4110 =  ( n3611 ) ? ( bv_8_36_n331 ) : ( n4109 ) ;
assign n4111 =  ( n3609 ) ? ( bv_8_92_n328 ) : ( n4110 ) ;
assign n4112 =  ( n3607 ) ? ( bv_8_194_n238 ) : ( n4111 ) ;
assign n4113 =  ( n3605 ) ? ( bv_8_211_n174 ) : ( n4112 ) ;
assign n4114 =  ( n3603 ) ? ( bv_8_172_n310 ) : ( n4113 ) ;
assign n4115 =  ( n3601 ) ? ( bv_8_98_n316 ) : ( n4114 ) ;
assign n4116 =  ( n3599 ) ? ( bv_8_145_n312 ) : ( n4115 ) ;
assign n4117 =  ( n3597 ) ? ( bv_8_149_n308 ) : ( n4116 ) ;
assign n4118 =  ( n3595 ) ? ( bv_8_228_n111 ) : ( n4117 ) ;
assign n4119 =  ( n3593 ) ? ( bv_8_121_n302 ) : ( n4118 ) ;
assign n4120 =  ( n3591 ) ? ( bv_8_231_n100 ) : ( n4119 ) ;
assign n4121 =  ( n3589 ) ? ( bv_8_200_n216 ) : ( n4120 ) ;
assign n4122 =  ( n3587 ) ? ( bv_8_55_n293 ) : ( n4121 ) ;
assign n4123 =  ( n3585 ) ? ( bv_8_109_n289 ) : ( n4122 ) ;
assign n4124 =  ( n3583 ) ? ( bv_8_141_n285 ) : ( n4123 ) ;
assign n4125 =  ( n3581 ) ? ( bv_8_213_n166 ) : ( n4124 ) ;
assign n4126 =  ( n3579 ) ? ( bv_8_78_n280 ) : ( n4125 ) ;
assign n4127 =  ( n3577 ) ? ( bv_8_169_n276 ) : ( n4126 ) ;
assign n4128 =  ( n3575 ) ? ( bv_8_108_n272 ) : ( n4127 ) ;
assign n4129 =  ( n3573 ) ? ( bv_8_86_n268 ) : ( n4128 ) ;
assign n4130 =  ( n3571 ) ? ( bv_8_244_n49 ) : ( n4129 ) ;
assign n4131 =  ( n3569 ) ? ( bv_8_234_n89 ) : ( n4130 ) ;
assign n4132 =  ( n3567 ) ? ( bv_8_101_n261 ) : ( n4131 ) ;
assign n4133 =  ( n3565 ) ? ( bv_8_122_n257 ) : ( n4132 ) ;
assign n4134 =  ( n3563 ) ? ( bv_8_174_n254 ) : ( n4133 ) ;
assign n4135 =  ( n3561 ) ? ( bv_8_8_n250 ) : ( n4134 ) ;
assign n4136 =  ( n3559 ) ? ( bv_8_186_n247 ) : ( n4135 ) ;
assign n4137 =  ( n3557 ) ? ( bv_8_120_n243 ) : ( n4136 ) ;
assign n4138 =  ( n3555 ) ? ( bv_8_37_n240 ) : ( n4137 ) ;
assign n4139 =  ( n3553 ) ? ( bv_8_46_n236 ) : ( n4138 ) ;
assign n4140 =  ( n3551 ) ? ( bv_8_28_n232 ) : ( n4139 ) ;
assign n4141 =  ( n3549 ) ? ( bv_8_166_n228 ) : ( n4140 ) ;
assign n4142 =  ( n3547 ) ? ( bv_8_180_n224 ) : ( n4141 ) ;
assign n4143 =  ( n3545 ) ? ( bv_8_198_n221 ) : ( n4142 ) ;
assign n4144 =  ( n3543 ) ? ( bv_8_232_n96 ) : ( n4143 ) ;
assign n4145 =  ( n3541 ) ? ( bv_8_221_n136 ) : ( n4144 ) ;
assign n4146 =  ( n3539 ) ? ( bv_8_116_n211 ) : ( n4145 ) ;
assign n4147 =  ( n3537 ) ? ( bv_8_31_n207 ) : ( n4146 ) ;
assign n4148 =  ( n3535 ) ? ( bv_8_75_n203 ) : ( n4147 ) ;
assign n4149 =  ( n3533 ) ? ( bv_8_189_n199 ) : ( n4148 ) ;
assign n4150 =  ( n3531 ) ? ( bv_8_139_n195 ) : ( n4149 ) ;
assign n4151 =  ( n3529 ) ? ( bv_8_138_n192 ) : ( n4150 ) ;
assign n4152 =  ( n3527 ) ? ( bv_8_112_n188 ) : ( n4151 ) ;
assign n4153 =  ( n3525 ) ? ( bv_8_62_n184 ) : ( n4152 ) ;
assign n4154 =  ( n3523 ) ? ( bv_8_181_n180 ) : ( n4153 ) ;
assign n4155 =  ( n3521 ) ? ( bv_8_102_n176 ) : ( n4154 ) ;
assign n4156 =  ( n3519 ) ? ( bv_8_72_n172 ) : ( n4155 ) ;
assign n4157 =  ( n3517 ) ? ( bv_8_3_n168 ) : ( n4156 ) ;
assign n4158 =  ( n3515 ) ? ( bv_8_246_n41 ) : ( n4157 ) ;
assign n4159 =  ( n3513 ) ? ( bv_8_14_n161 ) : ( n4158 ) ;
assign n4160 =  ( n3511 ) ? ( bv_8_97_n157 ) : ( n4159 ) ;
assign n4161 =  ( n3509 ) ? ( bv_8_53_n153 ) : ( n4160 ) ;
assign n4162 =  ( n3507 ) ? ( bv_8_87_n150 ) : ( n4161 ) ;
assign n4163 =  ( n3505 ) ? ( bv_8_185_n146 ) : ( n4162 ) ;
assign n4164 =  ( n3503 ) ? ( bv_8_134_n142 ) : ( n4163 ) ;
assign n4165 =  ( n3501 ) ? ( bv_8_193_n138 ) : ( n4164 ) ;
assign n4166 =  ( n3499 ) ? ( bv_8_29_n134 ) : ( n4165 ) ;
assign n4167 =  ( n3497 ) ? ( bv_8_158_n130 ) : ( n4166 ) ;
assign n4168 =  ( n3495 ) ? ( bv_8_225_n123 ) : ( n4167 ) ;
assign n4169 =  ( n3493 ) ? ( bv_8_248_n33 ) : ( n4168 ) ;
assign n4170 =  ( n3491 ) ? ( bv_8_152_n121 ) : ( n4169 ) ;
assign n4171 =  ( n3489 ) ? ( bv_8_17_n117 ) : ( n4170 ) ;
assign n4172 =  ( n3487 ) ? ( bv_8_105_n113 ) : ( n4171 ) ;
assign n4173 =  ( n3485 ) ? ( bv_8_217_n109 ) : ( n4172 ) ;
assign n4174 =  ( n3483 ) ? ( bv_8_142_n105 ) : ( n4173 ) ;
assign n4175 =  ( n3481 ) ? ( bv_8_148_n102 ) : ( n4174 ) ;
assign n4176 =  ( n3479 ) ? ( bv_8_155_n98 ) : ( n4175 ) ;
assign n4177 =  ( n3477 ) ? ( bv_8_30_n94 ) : ( n4176 ) ;
assign n4178 =  ( n3475 ) ? ( bv_8_135_n91 ) : ( n4177 ) ;
assign n4179 =  ( n3473 ) ? ( bv_8_233_n87 ) : ( n4178 ) ;
assign n4180 =  ( n3471 ) ? ( bv_8_206_n83 ) : ( n4179 ) ;
assign n4181 =  ( n3469 ) ? ( bv_8_85_n79 ) : ( n4180 ) ;
assign n4182 =  ( n3467 ) ? ( bv_8_40_n75 ) : ( n4181 ) ;
assign n4183 =  ( n3465 ) ? ( bv_8_223_n71 ) : ( n4182 ) ;
assign n4184 =  ( n3463 ) ? ( bv_8_140_n67 ) : ( n4183 ) ;
assign n4185 =  ( n3461 ) ? ( bv_8_161_n63 ) : ( n4184 ) ;
assign n4186 =  ( n3459 ) ? ( bv_8_137_n59 ) : ( n4185 ) ;
assign n4187 =  ( n3457 ) ? ( bv_8_13_n55 ) : ( n4186 ) ;
assign n4188 =  ( n3455 ) ? ( bv_8_191_n51 ) : ( n4187 ) ;
assign n4189 =  ( n3453 ) ? ( bv_8_230_n47 ) : ( n4188 ) ;
assign n4190 =  ( n3451 ) ? ( bv_8_66_n43 ) : ( n4189 ) ;
assign n4191 =  ( n3449 ) ? ( bv_8_104_n39 ) : ( n4190 ) ;
assign n4192 =  ( n3447 ) ? ( bv_8_65_n35 ) : ( n4191 ) ;
assign n4193 =  ( n3445 ) ? ( bv_8_153_n31 ) : ( n4192 ) ;
assign n4194 =  ( n3443 ) ? ( bv_8_45_n27 ) : ( n4193 ) ;
assign n4195 =  ( n3441 ) ? ( bv_8_15_n23 ) : ( n4194 ) ;
assign n4196 =  ( n3439 ) ? ( bv_8_176_n19 ) : ( n4195 ) ;
assign n4197 =  ( n3437 ) ? ( bv_8_84_n15 ) : ( n4196 ) ;
assign n4198 =  ( n3435 ) ? ( bv_8_187_n11 ) : ( n4197 ) ;
assign n4199 =  ( n3433 ) ? ( bv_8_22_n7 ) : ( n4198 ) ;
assign n4200 =  ( n3431 ) ^ ( n4199 )  ;
assign n4201 = in[119:112] ;
assign n4202 = in[15:8] ;
assign n4203 =  ( n4202 ) == ( bv_8_255_n5 )  ;
assign n4204 = in[15:8] ;
assign n4205 =  ( n4204 ) == ( bv_8_254_n9 )  ;
assign n4206 = in[15:8] ;
assign n4207 =  ( n4206 ) == ( bv_8_253_n13 )  ;
assign n4208 = in[15:8] ;
assign n4209 =  ( n4208 ) == ( bv_8_252_n17 )  ;
assign n4210 = in[15:8] ;
assign n4211 =  ( n4210 ) == ( bv_8_251_n21 )  ;
assign n4212 = in[15:8] ;
assign n4213 =  ( n4212 ) == ( bv_8_250_n25 )  ;
assign n4214 = in[15:8] ;
assign n4215 =  ( n4214 ) == ( bv_8_249_n29 )  ;
assign n4216 = in[15:8] ;
assign n4217 =  ( n4216 ) == ( bv_8_248_n33 )  ;
assign n4218 = in[15:8] ;
assign n4219 =  ( n4218 ) == ( bv_8_247_n37 )  ;
assign n4220 = in[15:8] ;
assign n4221 =  ( n4220 ) == ( bv_8_246_n41 )  ;
assign n4222 = in[15:8] ;
assign n4223 =  ( n4222 ) == ( bv_8_245_n45 )  ;
assign n4224 = in[15:8] ;
assign n4225 =  ( n4224 ) == ( bv_8_244_n49 )  ;
assign n4226 = in[15:8] ;
assign n4227 =  ( n4226 ) == ( bv_8_243_n53 )  ;
assign n4228 = in[15:8] ;
assign n4229 =  ( n4228 ) == ( bv_8_242_n57 )  ;
assign n4230 = in[15:8] ;
assign n4231 =  ( n4230 ) == ( bv_8_241_n61 )  ;
assign n4232 = in[15:8] ;
assign n4233 =  ( n4232 ) == ( bv_8_240_n65 )  ;
assign n4234 = in[15:8] ;
assign n4235 =  ( n4234 ) == ( bv_8_239_n69 )  ;
assign n4236 = in[15:8] ;
assign n4237 =  ( n4236 ) == ( bv_8_238_n73 )  ;
assign n4238 = in[15:8] ;
assign n4239 =  ( n4238 ) == ( bv_8_237_n77 )  ;
assign n4240 = in[15:8] ;
assign n4241 =  ( n4240 ) == ( bv_8_236_n81 )  ;
assign n4242 = in[15:8] ;
assign n4243 =  ( n4242 ) == ( bv_8_235_n85 )  ;
assign n4244 = in[15:8] ;
assign n4245 =  ( n4244 ) == ( bv_8_234_n89 )  ;
assign n4246 = in[15:8] ;
assign n4247 =  ( n4246 ) == ( bv_8_233_n87 )  ;
assign n4248 = in[15:8] ;
assign n4249 =  ( n4248 ) == ( bv_8_232_n96 )  ;
assign n4250 = in[15:8] ;
assign n4251 =  ( n4250 ) == ( bv_8_231_n100 )  ;
assign n4252 = in[15:8] ;
assign n4253 =  ( n4252 ) == ( bv_8_230_n47 )  ;
assign n4254 = in[15:8] ;
assign n4255 =  ( n4254 ) == ( bv_8_229_n107 )  ;
assign n4256 = in[15:8] ;
assign n4257 =  ( n4256 ) == ( bv_8_228_n111 )  ;
assign n4258 = in[15:8] ;
assign n4259 =  ( n4258 ) == ( bv_8_227_n115 )  ;
assign n4260 = in[15:8] ;
assign n4261 =  ( n4260 ) == ( bv_8_226_n119 )  ;
assign n4262 = in[15:8] ;
assign n4263 =  ( n4262 ) == ( bv_8_225_n123 )  ;
assign n4264 = in[15:8] ;
assign n4265 =  ( n4264 ) == ( bv_8_224_n126 )  ;
assign n4266 = in[15:8] ;
assign n4267 =  ( n4266 ) == ( bv_8_223_n71 )  ;
assign n4268 = in[15:8] ;
assign n4269 =  ( n4268 ) == ( bv_8_222_n132 )  ;
assign n4270 = in[15:8] ;
assign n4271 =  ( n4270 ) == ( bv_8_221_n136 )  ;
assign n4272 = in[15:8] ;
assign n4273 =  ( n4272 ) == ( bv_8_220_n140 )  ;
assign n4274 = in[15:8] ;
assign n4275 =  ( n4274 ) == ( bv_8_219_n144 )  ;
assign n4276 = in[15:8] ;
assign n4277 =  ( n4276 ) == ( bv_8_218_n148 )  ;
assign n4278 = in[15:8] ;
assign n4279 =  ( n4278 ) == ( bv_8_217_n109 )  ;
assign n4280 = in[15:8] ;
assign n4281 =  ( n4280 ) == ( bv_8_216_n155 )  ;
assign n4282 = in[15:8] ;
assign n4283 =  ( n4282 ) == ( bv_8_215_n159 )  ;
assign n4284 = in[15:8] ;
assign n4285 =  ( n4284 ) == ( bv_8_214_n163 )  ;
assign n4286 = in[15:8] ;
assign n4287 =  ( n4286 ) == ( bv_8_213_n166 )  ;
assign n4288 = in[15:8] ;
assign n4289 =  ( n4288 ) == ( bv_8_212_n170 )  ;
assign n4290 = in[15:8] ;
assign n4291 =  ( n4290 ) == ( bv_8_211_n174 )  ;
assign n4292 = in[15:8] ;
assign n4293 =  ( n4292 ) == ( bv_8_210_n178 )  ;
assign n4294 = in[15:8] ;
assign n4295 =  ( n4294 ) == ( bv_8_209_n182 )  ;
assign n4296 = in[15:8] ;
assign n4297 =  ( n4296 ) == ( bv_8_208_n186 )  ;
assign n4298 = in[15:8] ;
assign n4299 =  ( n4298 ) == ( bv_8_207_n190 )  ;
assign n4300 = in[15:8] ;
assign n4301 =  ( n4300 ) == ( bv_8_206_n83 )  ;
assign n4302 = in[15:8] ;
assign n4303 =  ( n4302 ) == ( bv_8_205_n197 )  ;
assign n4304 = in[15:8] ;
assign n4305 =  ( n4304 ) == ( bv_8_204_n201 )  ;
assign n4306 = in[15:8] ;
assign n4307 =  ( n4306 ) == ( bv_8_203_n205 )  ;
assign n4308 = in[15:8] ;
assign n4309 =  ( n4308 ) == ( bv_8_202_n209 )  ;
assign n4310 = in[15:8] ;
assign n4311 =  ( n4310 ) == ( bv_8_201_n213 )  ;
assign n4312 = in[15:8] ;
assign n4313 =  ( n4312 ) == ( bv_8_200_n216 )  ;
assign n4314 = in[15:8] ;
assign n4315 =  ( n4314 ) == ( bv_8_199_n219 )  ;
assign n4316 = in[15:8] ;
assign n4317 =  ( n4316 ) == ( bv_8_198_n221 )  ;
assign n4318 = in[15:8] ;
assign n4319 =  ( n4318 ) == ( bv_8_197_n226 )  ;
assign n4320 = in[15:8] ;
assign n4321 =  ( n4320 ) == ( bv_8_196_n230 )  ;
assign n4322 = in[15:8] ;
assign n4323 =  ( n4322 ) == ( bv_8_195_n234 )  ;
assign n4324 = in[15:8] ;
assign n4325 =  ( n4324 ) == ( bv_8_194_n238 )  ;
assign n4326 = in[15:8] ;
assign n4327 =  ( n4326 ) == ( bv_8_193_n138 )  ;
assign n4328 = in[15:8] ;
assign n4329 =  ( n4328 ) == ( bv_8_192_n245 )  ;
assign n4330 = in[15:8] ;
assign n4331 =  ( n4330 ) == ( bv_8_191_n51 )  ;
assign n4332 = in[15:8] ;
assign n4333 =  ( n4332 ) == ( bv_8_190_n252 )  ;
assign n4334 = in[15:8] ;
assign n4335 =  ( n4334 ) == ( bv_8_189_n199 )  ;
assign n4336 = in[15:8] ;
assign n4337 =  ( n4336 ) == ( bv_8_188_n259 )  ;
assign n4338 = in[15:8] ;
assign n4339 =  ( n4338 ) == ( bv_8_187_n11 )  ;
assign n4340 = in[15:8] ;
assign n4341 =  ( n4340 ) == ( bv_8_186_n247 )  ;
assign n4342 = in[15:8] ;
assign n4343 =  ( n4342 ) == ( bv_8_185_n146 )  ;
assign n4344 = in[15:8] ;
assign n4345 =  ( n4344 ) == ( bv_8_184_n270 )  ;
assign n4346 = in[15:8] ;
assign n4347 =  ( n4346 ) == ( bv_8_183_n274 )  ;
assign n4348 = in[15:8] ;
assign n4349 =  ( n4348 ) == ( bv_8_182_n278 )  ;
assign n4350 = in[15:8] ;
assign n4351 =  ( n4350 ) == ( bv_8_181_n180 )  ;
assign n4352 = in[15:8] ;
assign n4353 =  ( n4352 ) == ( bv_8_180_n224 )  ;
assign n4354 = in[15:8] ;
assign n4355 =  ( n4354 ) == ( bv_8_179_n287 )  ;
assign n4356 = in[15:8] ;
assign n4357 =  ( n4356 ) == ( bv_8_178_n291 )  ;
assign n4358 = in[15:8] ;
assign n4359 =  ( n4358 ) == ( bv_8_177_n295 )  ;
assign n4360 = in[15:8] ;
assign n4361 =  ( n4360 ) == ( bv_8_176_n19 )  ;
assign n4362 = in[15:8] ;
assign n4363 =  ( n4362 ) == ( bv_8_175_n300 )  ;
assign n4364 = in[15:8] ;
assign n4365 =  ( n4364 ) == ( bv_8_174_n254 )  ;
assign n4366 = in[15:8] ;
assign n4367 =  ( n4366 ) == ( bv_8_173_n306 )  ;
assign n4368 = in[15:8] ;
assign n4369 =  ( n4368 ) == ( bv_8_172_n310 )  ;
assign n4370 = in[15:8] ;
assign n4371 =  ( n4370 ) == ( bv_8_171_n314 )  ;
assign n4372 = in[15:8] ;
assign n4373 =  ( n4372 ) == ( bv_8_170_n318 )  ;
assign n4374 = in[15:8] ;
assign n4375 =  ( n4374 ) == ( bv_8_169_n276 )  ;
assign n4376 = in[15:8] ;
assign n4377 =  ( n4376 ) == ( bv_8_168_n323 )  ;
assign n4378 = in[15:8] ;
assign n4379 =  ( n4378 ) == ( bv_8_167_n326 )  ;
assign n4380 = in[15:8] ;
assign n4381 =  ( n4380 ) == ( bv_8_166_n228 )  ;
assign n4382 = in[15:8] ;
assign n4383 =  ( n4382 ) == ( bv_8_165_n333 )  ;
assign n4384 = in[15:8] ;
assign n4385 =  ( n4384 ) == ( bv_8_164_n337 )  ;
assign n4386 = in[15:8] ;
assign n4387 =  ( n4386 ) == ( bv_8_163_n341 )  ;
assign n4388 = in[15:8] ;
assign n4389 =  ( n4388 ) == ( bv_8_162_n345 )  ;
assign n4390 = in[15:8] ;
assign n4391 =  ( n4390 ) == ( bv_8_161_n63 )  ;
assign n4392 = in[15:8] ;
assign n4393 =  ( n4392 ) == ( bv_8_160_n352 )  ;
assign n4394 = in[15:8] ;
assign n4395 =  ( n4394 ) == ( bv_8_159_n355 )  ;
assign n4396 = in[15:8] ;
assign n4397 =  ( n4396 ) == ( bv_8_158_n130 )  ;
assign n4398 = in[15:8] ;
assign n4399 =  ( n4398 ) == ( bv_8_157_n361 )  ;
assign n4400 = in[15:8] ;
assign n4401 =  ( n4400 ) == ( bv_8_156_n365 )  ;
assign n4402 = in[15:8] ;
assign n4403 =  ( n4402 ) == ( bv_8_155_n98 )  ;
assign n4404 = in[15:8] ;
assign n4405 =  ( n4404 ) == ( bv_8_154_n371 )  ;
assign n4406 = in[15:8] ;
assign n4407 =  ( n4406 ) == ( bv_8_153_n31 )  ;
assign n4408 = in[15:8] ;
assign n4409 =  ( n4408 ) == ( bv_8_152_n121 )  ;
assign n4410 = in[15:8] ;
assign n4411 =  ( n4410 ) == ( bv_8_151_n379 )  ;
assign n4412 = in[15:8] ;
assign n4413 =  ( n4412 ) == ( bv_8_150_n383 )  ;
assign n4414 = in[15:8] ;
assign n4415 =  ( n4414 ) == ( bv_8_149_n308 )  ;
assign n4416 = in[15:8] ;
assign n4417 =  ( n4416 ) == ( bv_8_148_n102 )  ;
assign n4418 = in[15:8] ;
assign n4419 =  ( n4418 ) == ( bv_8_147_n393 )  ;
assign n4420 = in[15:8] ;
assign n4421 =  ( n4420 ) == ( bv_8_146_n396 )  ;
assign n4422 = in[15:8] ;
assign n4423 =  ( n4422 ) == ( bv_8_145_n312 )  ;
assign n4424 = in[15:8] ;
assign n4425 =  ( n4424 ) == ( bv_8_144_n385 )  ;
assign n4426 = in[15:8] ;
assign n4427 =  ( n4426 ) == ( bv_8_143_n406 )  ;
assign n4428 = in[15:8] ;
assign n4429 =  ( n4428 ) == ( bv_8_142_n105 )  ;
assign n4430 = in[15:8] ;
assign n4431 =  ( n4430 ) == ( bv_8_141_n285 )  ;
assign n4432 = in[15:8] ;
assign n4433 =  ( n4432 ) == ( bv_8_140_n67 )  ;
assign n4434 = in[15:8] ;
assign n4435 =  ( n4434 ) == ( bv_8_139_n195 )  ;
assign n4436 = in[15:8] ;
assign n4437 =  ( n4436 ) == ( bv_8_138_n192 )  ;
assign n4438 = in[15:8] ;
assign n4439 =  ( n4438 ) == ( bv_8_137_n59 )  ;
assign n4440 = in[15:8] ;
assign n4441 =  ( n4440 ) == ( bv_8_136_n381 )  ;
assign n4442 = in[15:8] ;
assign n4443 =  ( n4442 ) == ( bv_8_135_n91 )  ;
assign n4444 = in[15:8] ;
assign n4445 =  ( n4444 ) == ( bv_8_134_n142 )  ;
assign n4446 = in[15:8] ;
assign n4447 =  ( n4446 ) == ( bv_8_133_n435 )  ;
assign n4448 = in[15:8] ;
assign n4449 =  ( n4448 ) == ( bv_8_132_n438 )  ;
assign n4450 = in[15:8] ;
assign n4451 =  ( n4450 ) == ( bv_8_131_n442 )  ;
assign n4452 = in[15:8] ;
assign n4453 =  ( n4452 ) == ( bv_8_130_n445 )  ;
assign n4454 = in[15:8] ;
assign n4455 =  ( n4454 ) == ( bv_8_129_n401 )  ;
assign n4456 = in[15:8] ;
assign n4457 =  ( n4456 ) == ( bv_8_128_n452 )  ;
assign n4458 = in[15:8] ;
assign n4459 =  ( n4458 ) == ( bv_8_127_n455 )  ;
assign n4460 = in[15:8] ;
assign n4461 =  ( n4460 ) == ( bv_8_126_n423 )  ;
assign n4462 = in[15:8] ;
assign n4463 =  ( n4462 ) == ( bv_8_125_n460 )  ;
assign n4464 = in[15:8] ;
assign n4465 =  ( n4464 ) == ( bv_8_124_n463 )  ;
assign n4466 = in[15:8] ;
assign n4467 =  ( n4466 ) == ( bv_8_123_n467 )  ;
assign n4468 = in[15:8] ;
assign n4469 =  ( n4468 ) == ( bv_8_122_n257 )  ;
assign n4470 = in[15:8] ;
assign n4471 =  ( n4470 ) == ( bv_8_121_n302 )  ;
assign n4472 = in[15:8] ;
assign n4473 =  ( n4472 ) == ( bv_8_120_n243 )  ;
assign n4474 = in[15:8] ;
assign n4475 =  ( n4474 ) == ( bv_8_119_n477 )  ;
assign n4476 = in[15:8] ;
assign n4477 =  ( n4476 ) == ( bv_8_118_n480 )  ;
assign n4478 = in[15:8] ;
assign n4479 =  ( n4478 ) == ( bv_8_117_n484 )  ;
assign n4480 = in[15:8] ;
assign n4481 =  ( n4480 ) == ( bv_8_116_n211 )  ;
assign n4482 = in[15:8] ;
assign n4483 =  ( n4482 ) == ( bv_8_115_n408 )  ;
assign n4484 = in[15:8] ;
assign n4485 =  ( n4484 ) == ( bv_8_114_n491 )  ;
assign n4486 = in[15:8] ;
assign n4487 =  ( n4486 ) == ( bv_8_113_n495 )  ;
assign n4488 = in[15:8] ;
assign n4489 =  ( n4488 ) == ( bv_8_112_n188 )  ;
assign n4490 = in[15:8] ;
assign n4491 =  ( n4490 ) == ( bv_8_111_n501 )  ;
assign n4492 = in[15:8] ;
assign n4493 =  ( n4492 ) == ( bv_8_110_n504 )  ;
assign n4494 = in[15:8] ;
assign n4495 =  ( n4494 ) == ( bv_8_109_n289 )  ;
assign n4496 = in[15:8] ;
assign n4497 =  ( n4496 ) == ( bv_8_108_n272 )  ;
assign n4498 = in[15:8] ;
assign n4499 =  ( n4498 ) == ( bv_8_107_n513 )  ;
assign n4500 = in[15:8] ;
assign n4501 =  ( n4500 ) == ( bv_8_106_n516 )  ;
assign n4502 = in[15:8] ;
assign n4503 =  ( n4502 ) == ( bv_8_105_n113 )  ;
assign n4504 = in[15:8] ;
assign n4505 =  ( n4504 ) == ( bv_8_104_n39 )  ;
assign n4506 = in[15:8] ;
assign n4507 =  ( n4506 ) == ( bv_8_103_n525 )  ;
assign n4508 = in[15:8] ;
assign n4509 =  ( n4508 ) == ( bv_8_102_n176 )  ;
assign n4510 = in[15:8] ;
assign n4511 =  ( n4510 ) == ( bv_8_101_n261 )  ;
assign n4512 = in[15:8] ;
assign n4513 =  ( n4512 ) == ( bv_8_100_n417 )  ;
assign n4514 = in[15:8] ;
assign n4515 =  ( n4514 ) == ( bv_8_99_n537 )  ;
assign n4516 = in[15:8] ;
assign n4517 =  ( n4516 ) == ( bv_8_98_n316 )  ;
assign n4518 = in[15:8] ;
assign n4519 =  ( n4518 ) == ( bv_8_97_n157 )  ;
assign n4520 = in[15:8] ;
assign n4521 =  ( n4520 ) == ( bv_8_96_n404 )  ;
assign n4522 = in[15:8] ;
assign n4523 =  ( n4522 ) == ( bv_8_95_n440 )  ;
assign n4524 = in[15:8] ;
assign n4525 =  ( n4524 ) == ( bv_8_94_n363 )  ;
assign n4526 = in[15:8] ;
assign n4527 =  ( n4526 ) == ( bv_8_93_n414 )  ;
assign n4528 = in[15:8] ;
assign n4529 =  ( n4528 ) == ( bv_8_92_n328 )  ;
assign n4530 = in[15:8] ;
assign n4531 =  ( n4530 ) == ( bv_8_91_n557 )  ;
assign n4532 = in[15:8] ;
assign n4533 =  ( n4532 ) == ( bv_8_90_n561 )  ;
assign n4534 = in[15:8] ;
assign n4535 =  ( n4534 ) == ( bv_8_89_n564 )  ;
assign n4536 = in[15:8] ;
assign n4537 =  ( n4536 ) == ( bv_8_88_n549 )  ;
assign n4538 = in[15:8] ;
assign n4539 =  ( n4538 ) == ( bv_8_87_n150 )  ;
assign n4540 = in[15:8] ;
assign n4541 =  ( n4540 ) == ( bv_8_86_n268 )  ;
assign n4542 = in[15:8] ;
assign n4543 =  ( n4542 ) == ( bv_8_85_n79 )  ;
assign n4544 = in[15:8] ;
assign n4545 =  ( n4544 ) == ( bv_8_84_n15 )  ;
assign n4546 = in[15:8] ;
assign n4547 =  ( n4546 ) == ( bv_8_83_n578 )  ;
assign n4548 = in[15:8] ;
assign n4549 =  ( n4548 ) == ( bv_8_82_n581 )  ;
assign n4550 = in[15:8] ;
assign n4551 =  ( n4550 ) == ( bv_8_81_n499 )  ;
assign n4552 = in[15:8] ;
assign n4553 =  ( n4552 ) == ( bv_8_80_n511 )  ;
assign n4554 = in[15:8] ;
assign n4555 =  ( n4554 ) == ( bv_8_79_n398 )  ;
assign n4556 = in[15:8] ;
assign n4557 =  ( n4556 ) == ( bv_8_78_n280 )  ;
assign n4558 = in[15:8] ;
assign n4559 =  ( n4558 ) == ( bv_8_77_n532 )  ;
assign n4560 = in[15:8] ;
assign n4561 =  ( n4560 ) == ( bv_8_76_n552 )  ;
assign n4562 = in[15:8] ;
assign n4563 =  ( n4562 ) == ( bv_8_75_n203 )  ;
assign n4564 = in[15:8] ;
assign n4565 =  ( n4564 ) == ( bv_8_74_n555 )  ;
assign n4566 = in[15:8] ;
assign n4567 =  ( n4566 ) == ( bv_8_73_n339 )  ;
assign n4568 = in[15:8] ;
assign n4569 =  ( n4568 ) == ( bv_8_72_n172 )  ;
assign n4570 = in[15:8] ;
assign n4571 =  ( n4570 ) == ( bv_8_71_n608 )  ;
assign n4572 = in[15:8] ;
assign n4573 =  ( n4572 ) == ( bv_8_70_n377 )  ;
assign n4574 = in[15:8] ;
assign n4575 =  ( n4574 ) == ( bv_8_69_n523 )  ;
assign n4576 = in[15:8] ;
assign n4577 =  ( n4576 ) == ( bv_8_68_n433 )  ;
assign n4578 = in[15:8] ;
assign n4579 =  ( n4578 ) == ( bv_8_67_n535 )  ;
assign n4580 = in[15:8] ;
assign n4581 =  ( n4580 ) == ( bv_8_66_n43 )  ;
assign n4582 = in[15:8] ;
assign n4583 =  ( n4582 ) == ( bv_8_65_n35 )  ;
assign n4584 = in[15:8] ;
assign n4585 =  ( n4584 ) == ( bv_8_64_n493 )  ;
assign n4586 = in[15:8] ;
assign n4587 =  ( n4586 ) == ( bv_8_63_n629 )  ;
assign n4588 = in[15:8] ;
assign n4589 =  ( n4588 ) == ( bv_8_62_n184 )  ;
assign n4590 = in[15:8] ;
assign n4591 =  ( n4590 ) == ( bv_8_61_n420 )  ;
assign n4592 = in[15:8] ;
assign n4593 =  ( n4592 ) == ( bv_8_60_n508 )  ;
assign n4594 = in[15:8] ;
assign n4595 =  ( n4594 ) == ( bv_8_59_n604 )  ;
assign n4596 = in[15:8] ;
assign n4597 =  ( n4596 ) == ( bv_8_58_n347 )  ;
assign n4598 = in[15:8] ;
assign n4599 =  ( n4598 ) == ( bv_8_57_n559 )  ;
assign n4600 = in[15:8] ;
assign n4601 =  ( n4600 ) == ( bv_8_56_n482 )  ;
assign n4602 = in[15:8] ;
assign n4603 =  ( n4602 ) == ( bv_8_55_n293 )  ;
assign n4604 = in[15:8] ;
assign n4605 =  ( n4604 ) == ( bv_8_54_n651 )  ;
assign n4606 = in[15:8] ;
assign n4607 =  ( n4606 ) == ( bv_8_53_n153 )  ;
assign n4608 = in[15:8] ;
assign n4609 =  ( n4608 ) == ( bv_8_52_n657 )  ;
assign n4610 = in[15:8] ;
assign n4611 =  ( n4610 ) == ( bv_8_51_n529 )  ;
assign n4612 = in[15:8] ;
assign n4613 =  ( n4612 ) == ( bv_8_50_n350 )  ;
assign n4614 = in[15:8] ;
assign n4615 =  ( n4614 ) == ( bv_8_49_n666 )  ;
assign n4616 = in[15:8] ;
assign n4617 =  ( n4616 ) == ( bv_8_48_n669 )  ;
assign n4618 = in[15:8] ;
assign n4619 =  ( n4618 ) == ( bv_8_47_n592 )  ;
assign n4620 = in[15:8] ;
assign n4621 =  ( n4620 ) == ( bv_8_46_n236 )  ;
assign n4622 = in[15:8] ;
assign n4623 =  ( n4622 ) == ( bv_8_45_n27 )  ;
assign n4624 = in[15:8] ;
assign n4625 =  ( n4624 ) == ( bv_8_44_n622 )  ;
assign n4626 = in[15:8] ;
assign n4627 =  ( n4626 ) == ( bv_8_43_n682 )  ;
assign n4628 = in[15:8] ;
assign n4629 =  ( n4628 ) == ( bv_8_42_n388 )  ;
assign n4630 = in[15:8] ;
assign n4631 =  ( n4630 ) == ( bv_8_41_n597 )  ;
assign n4632 = in[15:8] ;
assign n4633 =  ( n4632 ) == ( bv_8_40_n75 )  ;
assign n4634 = in[15:8] ;
assign n4635 =  ( n4634 ) == ( bv_8_39_n635 )  ;
assign n4636 = in[15:8] ;
assign n4637 =  ( n4636 ) == ( bv_8_38_n693 )  ;
assign n4638 = in[15:8] ;
assign n4639 =  ( n4638 ) == ( bv_8_37_n240 )  ;
assign n4640 = in[15:8] ;
assign n4641 =  ( n4640 ) == ( bv_8_36_n331 )  ;
assign n4642 = in[15:8] ;
assign n4643 =  ( n4642 ) == ( bv_8_35_n664 )  ;
assign n4644 = in[15:8] ;
assign n4645 =  ( n4644 ) == ( bv_8_34_n391 )  ;
assign n4646 = in[15:8] ;
assign n4647 =  ( n4646 ) == ( bv_8_33_n469 )  ;
assign n4648 = in[15:8] ;
assign n4649 =  ( n4648 ) == ( bv_8_32_n576 )  ;
assign n4650 = in[15:8] ;
assign n4651 =  ( n4650 ) == ( bv_8_31_n207 )  ;
assign n4652 = in[15:8] ;
assign n4653 =  ( n4652 ) == ( bv_8_30_n94 )  ;
assign n4654 = in[15:8] ;
assign n4655 =  ( n4654 ) == ( bv_8_29_n134 )  ;
assign n4656 = in[15:8] ;
assign n4657 =  ( n4656 ) == ( bv_8_28_n232 )  ;
assign n4658 = in[15:8] ;
assign n4659 =  ( n4658 ) == ( bv_8_27_n616 )  ;
assign n4660 = in[15:8] ;
assign n4661 =  ( n4660 ) == ( bv_8_26_n619 )  ;
assign n4662 = in[15:8] ;
assign n4663 =  ( n4662 ) == ( bv_8_25_n411 )  ;
assign n4664 = in[15:8] ;
assign n4665 =  ( n4664 ) == ( bv_8_24_n659 )  ;
assign n4666 = in[15:8] ;
assign n4667 =  ( n4666 ) == ( bv_8_23_n430 )  ;
assign n4668 = in[15:8] ;
assign n4669 =  ( n4668 ) == ( bv_8_22_n7 )  ;
assign n4670 = in[15:8] ;
assign n4671 =  ( n4670 ) == ( bv_8_21_n674 )  ;
assign n4672 = in[15:8] ;
assign n4673 =  ( n4672 ) == ( bv_8_20_n369 )  ;
assign n4674 = in[15:8] ;
assign n4675 =  ( n4674 ) == ( bv_8_19_n447 )  ;
assign n4676 = in[15:8] ;
assign n4677 =  ( n4676 ) == ( bv_8_18_n644 )  ;
assign n4678 = in[15:8] ;
assign n4679 =  ( n4678 ) == ( bv_8_17_n117 )  ;
assign n4680 = in[15:8] ;
assign n4681 =  ( n4680 ) == ( bv_8_16_n465 )  ;
assign n4682 = in[15:8] ;
assign n4683 =  ( n4682 ) == ( bv_8_15_n23 )  ;
assign n4684 = in[15:8] ;
assign n4685 =  ( n4684 ) == ( bv_8_14_n161 )  ;
assign n4686 = in[15:8] ;
assign n4687 =  ( n4686 ) == ( bv_8_13_n55 )  ;
assign n4688 = in[15:8] ;
assign n4689 =  ( n4688 ) == ( bv_8_12_n450 )  ;
assign n4690 = in[15:8] ;
assign n4691 =  ( n4690 ) == ( bv_8_11_n359 )  ;
assign n4692 = in[15:8] ;
assign n4693 =  ( n4692 ) == ( bv_8_10_n343 )  ;
assign n4694 = in[15:8] ;
assign n4695 =  ( n4694 ) == ( bv_8_9_n627 )  ;
assign n4696 = in[15:8] ;
assign n4697 =  ( n4696 ) == ( bv_8_8_n250 )  ;
assign n4698 = in[15:8] ;
assign n4699 =  ( n4698 ) == ( bv_8_7_n647 )  ;
assign n4700 = in[15:8] ;
assign n4701 =  ( n4700 ) == ( bv_8_6_n335 )  ;
assign n4702 = in[15:8] ;
assign n4703 =  ( n4702 ) == ( bv_8_5_n653 )  ;
assign n4704 = in[15:8] ;
assign n4705 =  ( n4704 ) == ( bv_8_4_n671 )  ;
assign n4706 = in[15:8] ;
assign n4707 =  ( n4706 ) == ( bv_8_3_n168 )  ;
assign n4708 = in[15:8] ;
assign n4709 =  ( n4708 ) == ( bv_8_2_n518 )  ;
assign n4710 = in[15:8] ;
assign n4711 =  ( n4710 ) == ( bv_8_1_n753 )  ;
assign n4712 = in[15:8] ;
assign n4713 =  ( n4712 ) == ( bv_8_0_n583 )  ;
assign n4714 =  ( n4713 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n4715 =  ( n4711 ) ? ( bv_8_124_n463 ) : ( n4714 ) ;
assign n4716 =  ( n4709 ) ? ( bv_8_119_n477 ) : ( n4715 ) ;
assign n4717 =  ( n4707 ) ? ( bv_8_123_n467 ) : ( n4716 ) ;
assign n4718 =  ( n4705 ) ? ( bv_8_242_n57 ) : ( n4717 ) ;
assign n4719 =  ( n4703 ) ? ( bv_8_107_n513 ) : ( n4718 ) ;
assign n4720 =  ( n4701 ) ? ( bv_8_111_n501 ) : ( n4719 ) ;
assign n4721 =  ( n4699 ) ? ( bv_8_197_n226 ) : ( n4720 ) ;
assign n4722 =  ( n4697 ) ? ( bv_8_48_n669 ) : ( n4721 ) ;
assign n4723 =  ( n4695 ) ? ( bv_8_1_n753 ) : ( n4722 ) ;
assign n4724 =  ( n4693 ) ? ( bv_8_103_n525 ) : ( n4723 ) ;
assign n4725 =  ( n4691 ) ? ( bv_8_43_n682 ) : ( n4724 ) ;
assign n4726 =  ( n4689 ) ? ( bv_8_254_n9 ) : ( n4725 ) ;
assign n4727 =  ( n4687 ) ? ( bv_8_215_n159 ) : ( n4726 ) ;
assign n4728 =  ( n4685 ) ? ( bv_8_171_n314 ) : ( n4727 ) ;
assign n4729 =  ( n4683 ) ? ( bv_8_118_n480 ) : ( n4728 ) ;
assign n4730 =  ( n4681 ) ? ( bv_8_202_n209 ) : ( n4729 ) ;
assign n4731 =  ( n4679 ) ? ( bv_8_130_n445 ) : ( n4730 ) ;
assign n4732 =  ( n4677 ) ? ( bv_8_201_n213 ) : ( n4731 ) ;
assign n4733 =  ( n4675 ) ? ( bv_8_125_n460 ) : ( n4732 ) ;
assign n4734 =  ( n4673 ) ? ( bv_8_250_n25 ) : ( n4733 ) ;
assign n4735 =  ( n4671 ) ? ( bv_8_89_n564 ) : ( n4734 ) ;
assign n4736 =  ( n4669 ) ? ( bv_8_71_n608 ) : ( n4735 ) ;
assign n4737 =  ( n4667 ) ? ( bv_8_240_n65 ) : ( n4736 ) ;
assign n4738 =  ( n4665 ) ? ( bv_8_173_n306 ) : ( n4737 ) ;
assign n4739 =  ( n4663 ) ? ( bv_8_212_n170 ) : ( n4738 ) ;
assign n4740 =  ( n4661 ) ? ( bv_8_162_n345 ) : ( n4739 ) ;
assign n4741 =  ( n4659 ) ? ( bv_8_175_n300 ) : ( n4740 ) ;
assign n4742 =  ( n4657 ) ? ( bv_8_156_n365 ) : ( n4741 ) ;
assign n4743 =  ( n4655 ) ? ( bv_8_164_n337 ) : ( n4742 ) ;
assign n4744 =  ( n4653 ) ? ( bv_8_114_n491 ) : ( n4743 ) ;
assign n4745 =  ( n4651 ) ? ( bv_8_192_n245 ) : ( n4744 ) ;
assign n4746 =  ( n4649 ) ? ( bv_8_183_n274 ) : ( n4745 ) ;
assign n4747 =  ( n4647 ) ? ( bv_8_253_n13 ) : ( n4746 ) ;
assign n4748 =  ( n4645 ) ? ( bv_8_147_n393 ) : ( n4747 ) ;
assign n4749 =  ( n4643 ) ? ( bv_8_38_n693 ) : ( n4748 ) ;
assign n4750 =  ( n4641 ) ? ( bv_8_54_n651 ) : ( n4749 ) ;
assign n4751 =  ( n4639 ) ? ( bv_8_63_n629 ) : ( n4750 ) ;
assign n4752 =  ( n4637 ) ? ( bv_8_247_n37 ) : ( n4751 ) ;
assign n4753 =  ( n4635 ) ? ( bv_8_204_n201 ) : ( n4752 ) ;
assign n4754 =  ( n4633 ) ? ( bv_8_52_n657 ) : ( n4753 ) ;
assign n4755 =  ( n4631 ) ? ( bv_8_165_n333 ) : ( n4754 ) ;
assign n4756 =  ( n4629 ) ? ( bv_8_229_n107 ) : ( n4755 ) ;
assign n4757 =  ( n4627 ) ? ( bv_8_241_n61 ) : ( n4756 ) ;
assign n4758 =  ( n4625 ) ? ( bv_8_113_n495 ) : ( n4757 ) ;
assign n4759 =  ( n4623 ) ? ( bv_8_216_n155 ) : ( n4758 ) ;
assign n4760 =  ( n4621 ) ? ( bv_8_49_n666 ) : ( n4759 ) ;
assign n4761 =  ( n4619 ) ? ( bv_8_21_n674 ) : ( n4760 ) ;
assign n4762 =  ( n4617 ) ? ( bv_8_4_n671 ) : ( n4761 ) ;
assign n4763 =  ( n4615 ) ? ( bv_8_199_n219 ) : ( n4762 ) ;
assign n4764 =  ( n4613 ) ? ( bv_8_35_n664 ) : ( n4763 ) ;
assign n4765 =  ( n4611 ) ? ( bv_8_195_n234 ) : ( n4764 ) ;
assign n4766 =  ( n4609 ) ? ( bv_8_24_n659 ) : ( n4765 ) ;
assign n4767 =  ( n4607 ) ? ( bv_8_150_n383 ) : ( n4766 ) ;
assign n4768 =  ( n4605 ) ? ( bv_8_5_n653 ) : ( n4767 ) ;
assign n4769 =  ( n4603 ) ? ( bv_8_154_n371 ) : ( n4768 ) ;
assign n4770 =  ( n4601 ) ? ( bv_8_7_n647 ) : ( n4769 ) ;
assign n4771 =  ( n4599 ) ? ( bv_8_18_n644 ) : ( n4770 ) ;
assign n4772 =  ( n4597 ) ? ( bv_8_128_n452 ) : ( n4771 ) ;
assign n4773 =  ( n4595 ) ? ( bv_8_226_n119 ) : ( n4772 ) ;
assign n4774 =  ( n4593 ) ? ( bv_8_235_n85 ) : ( n4773 ) ;
assign n4775 =  ( n4591 ) ? ( bv_8_39_n635 ) : ( n4774 ) ;
assign n4776 =  ( n4589 ) ? ( bv_8_178_n291 ) : ( n4775 ) ;
assign n4777 =  ( n4587 ) ? ( bv_8_117_n484 ) : ( n4776 ) ;
assign n4778 =  ( n4585 ) ? ( bv_8_9_n627 ) : ( n4777 ) ;
assign n4779 =  ( n4583 ) ? ( bv_8_131_n442 ) : ( n4778 ) ;
assign n4780 =  ( n4581 ) ? ( bv_8_44_n622 ) : ( n4779 ) ;
assign n4781 =  ( n4579 ) ? ( bv_8_26_n619 ) : ( n4780 ) ;
assign n4782 =  ( n4577 ) ? ( bv_8_27_n616 ) : ( n4781 ) ;
assign n4783 =  ( n4575 ) ? ( bv_8_110_n504 ) : ( n4782 ) ;
assign n4784 =  ( n4573 ) ? ( bv_8_90_n561 ) : ( n4783 ) ;
assign n4785 =  ( n4571 ) ? ( bv_8_160_n352 ) : ( n4784 ) ;
assign n4786 =  ( n4569 ) ? ( bv_8_82_n581 ) : ( n4785 ) ;
assign n4787 =  ( n4567 ) ? ( bv_8_59_n604 ) : ( n4786 ) ;
assign n4788 =  ( n4565 ) ? ( bv_8_214_n163 ) : ( n4787 ) ;
assign n4789 =  ( n4563 ) ? ( bv_8_179_n287 ) : ( n4788 ) ;
assign n4790 =  ( n4561 ) ? ( bv_8_41_n597 ) : ( n4789 ) ;
assign n4791 =  ( n4559 ) ? ( bv_8_227_n115 ) : ( n4790 ) ;
assign n4792 =  ( n4557 ) ? ( bv_8_47_n592 ) : ( n4791 ) ;
assign n4793 =  ( n4555 ) ? ( bv_8_132_n438 ) : ( n4792 ) ;
assign n4794 =  ( n4553 ) ? ( bv_8_83_n578 ) : ( n4793 ) ;
assign n4795 =  ( n4551 ) ? ( bv_8_209_n182 ) : ( n4794 ) ;
assign n4796 =  ( n4549 ) ? ( bv_8_0_n583 ) : ( n4795 ) ;
assign n4797 =  ( n4547 ) ? ( bv_8_237_n77 ) : ( n4796 ) ;
assign n4798 =  ( n4545 ) ? ( bv_8_32_n576 ) : ( n4797 ) ;
assign n4799 =  ( n4543 ) ? ( bv_8_252_n17 ) : ( n4798 ) ;
assign n4800 =  ( n4541 ) ? ( bv_8_177_n295 ) : ( n4799 ) ;
assign n4801 =  ( n4539 ) ? ( bv_8_91_n557 ) : ( n4800 ) ;
assign n4802 =  ( n4537 ) ? ( bv_8_106_n516 ) : ( n4801 ) ;
assign n4803 =  ( n4535 ) ? ( bv_8_203_n205 ) : ( n4802 ) ;
assign n4804 =  ( n4533 ) ? ( bv_8_190_n252 ) : ( n4803 ) ;
assign n4805 =  ( n4531 ) ? ( bv_8_57_n559 ) : ( n4804 ) ;
assign n4806 =  ( n4529 ) ? ( bv_8_74_n555 ) : ( n4805 ) ;
assign n4807 =  ( n4527 ) ? ( bv_8_76_n552 ) : ( n4806 ) ;
assign n4808 =  ( n4525 ) ? ( bv_8_88_n549 ) : ( n4807 ) ;
assign n4809 =  ( n4523 ) ? ( bv_8_207_n190 ) : ( n4808 ) ;
assign n4810 =  ( n4521 ) ? ( bv_8_208_n186 ) : ( n4809 ) ;
assign n4811 =  ( n4519 ) ? ( bv_8_239_n69 ) : ( n4810 ) ;
assign n4812 =  ( n4517 ) ? ( bv_8_170_n318 ) : ( n4811 ) ;
assign n4813 =  ( n4515 ) ? ( bv_8_251_n21 ) : ( n4812 ) ;
assign n4814 =  ( n4513 ) ? ( bv_8_67_n535 ) : ( n4813 ) ;
assign n4815 =  ( n4511 ) ? ( bv_8_77_n532 ) : ( n4814 ) ;
assign n4816 =  ( n4509 ) ? ( bv_8_51_n529 ) : ( n4815 ) ;
assign n4817 =  ( n4507 ) ? ( bv_8_133_n435 ) : ( n4816 ) ;
assign n4818 =  ( n4505 ) ? ( bv_8_69_n523 ) : ( n4817 ) ;
assign n4819 =  ( n4503 ) ? ( bv_8_249_n29 ) : ( n4818 ) ;
assign n4820 =  ( n4501 ) ? ( bv_8_2_n518 ) : ( n4819 ) ;
assign n4821 =  ( n4499 ) ? ( bv_8_127_n455 ) : ( n4820 ) ;
assign n4822 =  ( n4497 ) ? ( bv_8_80_n511 ) : ( n4821 ) ;
assign n4823 =  ( n4495 ) ? ( bv_8_60_n508 ) : ( n4822 ) ;
assign n4824 =  ( n4493 ) ? ( bv_8_159_n355 ) : ( n4823 ) ;
assign n4825 =  ( n4491 ) ? ( bv_8_168_n323 ) : ( n4824 ) ;
assign n4826 =  ( n4489 ) ? ( bv_8_81_n499 ) : ( n4825 ) ;
assign n4827 =  ( n4487 ) ? ( bv_8_163_n341 ) : ( n4826 ) ;
assign n4828 =  ( n4485 ) ? ( bv_8_64_n493 ) : ( n4827 ) ;
assign n4829 =  ( n4483 ) ? ( bv_8_143_n406 ) : ( n4828 ) ;
assign n4830 =  ( n4481 ) ? ( bv_8_146_n396 ) : ( n4829 ) ;
assign n4831 =  ( n4479 ) ? ( bv_8_157_n361 ) : ( n4830 ) ;
assign n4832 =  ( n4477 ) ? ( bv_8_56_n482 ) : ( n4831 ) ;
assign n4833 =  ( n4475 ) ? ( bv_8_245_n45 ) : ( n4832 ) ;
assign n4834 =  ( n4473 ) ? ( bv_8_188_n259 ) : ( n4833 ) ;
assign n4835 =  ( n4471 ) ? ( bv_8_182_n278 ) : ( n4834 ) ;
assign n4836 =  ( n4469 ) ? ( bv_8_218_n148 ) : ( n4835 ) ;
assign n4837 =  ( n4467 ) ? ( bv_8_33_n469 ) : ( n4836 ) ;
assign n4838 =  ( n4465 ) ? ( bv_8_16_n465 ) : ( n4837 ) ;
assign n4839 =  ( n4463 ) ? ( bv_8_255_n5 ) : ( n4838 ) ;
assign n4840 =  ( n4461 ) ? ( bv_8_243_n53 ) : ( n4839 ) ;
assign n4841 =  ( n4459 ) ? ( bv_8_210_n178 ) : ( n4840 ) ;
assign n4842 =  ( n4457 ) ? ( bv_8_205_n197 ) : ( n4841 ) ;
assign n4843 =  ( n4455 ) ? ( bv_8_12_n450 ) : ( n4842 ) ;
assign n4844 =  ( n4453 ) ? ( bv_8_19_n447 ) : ( n4843 ) ;
assign n4845 =  ( n4451 ) ? ( bv_8_236_n81 ) : ( n4844 ) ;
assign n4846 =  ( n4449 ) ? ( bv_8_95_n440 ) : ( n4845 ) ;
assign n4847 =  ( n4447 ) ? ( bv_8_151_n379 ) : ( n4846 ) ;
assign n4848 =  ( n4445 ) ? ( bv_8_68_n433 ) : ( n4847 ) ;
assign n4849 =  ( n4443 ) ? ( bv_8_23_n430 ) : ( n4848 ) ;
assign n4850 =  ( n4441 ) ? ( bv_8_196_n230 ) : ( n4849 ) ;
assign n4851 =  ( n4439 ) ? ( bv_8_167_n326 ) : ( n4850 ) ;
assign n4852 =  ( n4437 ) ? ( bv_8_126_n423 ) : ( n4851 ) ;
assign n4853 =  ( n4435 ) ? ( bv_8_61_n420 ) : ( n4852 ) ;
assign n4854 =  ( n4433 ) ? ( bv_8_100_n417 ) : ( n4853 ) ;
assign n4855 =  ( n4431 ) ? ( bv_8_93_n414 ) : ( n4854 ) ;
assign n4856 =  ( n4429 ) ? ( bv_8_25_n411 ) : ( n4855 ) ;
assign n4857 =  ( n4427 ) ? ( bv_8_115_n408 ) : ( n4856 ) ;
assign n4858 =  ( n4425 ) ? ( bv_8_96_n404 ) : ( n4857 ) ;
assign n4859 =  ( n4423 ) ? ( bv_8_129_n401 ) : ( n4858 ) ;
assign n4860 =  ( n4421 ) ? ( bv_8_79_n398 ) : ( n4859 ) ;
assign n4861 =  ( n4419 ) ? ( bv_8_220_n140 ) : ( n4860 ) ;
assign n4862 =  ( n4417 ) ? ( bv_8_34_n391 ) : ( n4861 ) ;
assign n4863 =  ( n4415 ) ? ( bv_8_42_n388 ) : ( n4862 ) ;
assign n4864 =  ( n4413 ) ? ( bv_8_144_n385 ) : ( n4863 ) ;
assign n4865 =  ( n4411 ) ? ( bv_8_136_n381 ) : ( n4864 ) ;
assign n4866 =  ( n4409 ) ? ( bv_8_70_n377 ) : ( n4865 ) ;
assign n4867 =  ( n4407 ) ? ( bv_8_238_n73 ) : ( n4866 ) ;
assign n4868 =  ( n4405 ) ? ( bv_8_184_n270 ) : ( n4867 ) ;
assign n4869 =  ( n4403 ) ? ( bv_8_20_n369 ) : ( n4868 ) ;
assign n4870 =  ( n4401 ) ? ( bv_8_222_n132 ) : ( n4869 ) ;
assign n4871 =  ( n4399 ) ? ( bv_8_94_n363 ) : ( n4870 ) ;
assign n4872 =  ( n4397 ) ? ( bv_8_11_n359 ) : ( n4871 ) ;
assign n4873 =  ( n4395 ) ? ( bv_8_219_n144 ) : ( n4872 ) ;
assign n4874 =  ( n4393 ) ? ( bv_8_224_n126 ) : ( n4873 ) ;
assign n4875 =  ( n4391 ) ? ( bv_8_50_n350 ) : ( n4874 ) ;
assign n4876 =  ( n4389 ) ? ( bv_8_58_n347 ) : ( n4875 ) ;
assign n4877 =  ( n4387 ) ? ( bv_8_10_n343 ) : ( n4876 ) ;
assign n4878 =  ( n4385 ) ? ( bv_8_73_n339 ) : ( n4877 ) ;
assign n4879 =  ( n4383 ) ? ( bv_8_6_n335 ) : ( n4878 ) ;
assign n4880 =  ( n4381 ) ? ( bv_8_36_n331 ) : ( n4879 ) ;
assign n4881 =  ( n4379 ) ? ( bv_8_92_n328 ) : ( n4880 ) ;
assign n4882 =  ( n4377 ) ? ( bv_8_194_n238 ) : ( n4881 ) ;
assign n4883 =  ( n4375 ) ? ( bv_8_211_n174 ) : ( n4882 ) ;
assign n4884 =  ( n4373 ) ? ( bv_8_172_n310 ) : ( n4883 ) ;
assign n4885 =  ( n4371 ) ? ( bv_8_98_n316 ) : ( n4884 ) ;
assign n4886 =  ( n4369 ) ? ( bv_8_145_n312 ) : ( n4885 ) ;
assign n4887 =  ( n4367 ) ? ( bv_8_149_n308 ) : ( n4886 ) ;
assign n4888 =  ( n4365 ) ? ( bv_8_228_n111 ) : ( n4887 ) ;
assign n4889 =  ( n4363 ) ? ( bv_8_121_n302 ) : ( n4888 ) ;
assign n4890 =  ( n4361 ) ? ( bv_8_231_n100 ) : ( n4889 ) ;
assign n4891 =  ( n4359 ) ? ( bv_8_200_n216 ) : ( n4890 ) ;
assign n4892 =  ( n4357 ) ? ( bv_8_55_n293 ) : ( n4891 ) ;
assign n4893 =  ( n4355 ) ? ( bv_8_109_n289 ) : ( n4892 ) ;
assign n4894 =  ( n4353 ) ? ( bv_8_141_n285 ) : ( n4893 ) ;
assign n4895 =  ( n4351 ) ? ( bv_8_213_n166 ) : ( n4894 ) ;
assign n4896 =  ( n4349 ) ? ( bv_8_78_n280 ) : ( n4895 ) ;
assign n4897 =  ( n4347 ) ? ( bv_8_169_n276 ) : ( n4896 ) ;
assign n4898 =  ( n4345 ) ? ( bv_8_108_n272 ) : ( n4897 ) ;
assign n4899 =  ( n4343 ) ? ( bv_8_86_n268 ) : ( n4898 ) ;
assign n4900 =  ( n4341 ) ? ( bv_8_244_n49 ) : ( n4899 ) ;
assign n4901 =  ( n4339 ) ? ( bv_8_234_n89 ) : ( n4900 ) ;
assign n4902 =  ( n4337 ) ? ( bv_8_101_n261 ) : ( n4901 ) ;
assign n4903 =  ( n4335 ) ? ( bv_8_122_n257 ) : ( n4902 ) ;
assign n4904 =  ( n4333 ) ? ( bv_8_174_n254 ) : ( n4903 ) ;
assign n4905 =  ( n4331 ) ? ( bv_8_8_n250 ) : ( n4904 ) ;
assign n4906 =  ( n4329 ) ? ( bv_8_186_n247 ) : ( n4905 ) ;
assign n4907 =  ( n4327 ) ? ( bv_8_120_n243 ) : ( n4906 ) ;
assign n4908 =  ( n4325 ) ? ( bv_8_37_n240 ) : ( n4907 ) ;
assign n4909 =  ( n4323 ) ? ( bv_8_46_n236 ) : ( n4908 ) ;
assign n4910 =  ( n4321 ) ? ( bv_8_28_n232 ) : ( n4909 ) ;
assign n4911 =  ( n4319 ) ? ( bv_8_166_n228 ) : ( n4910 ) ;
assign n4912 =  ( n4317 ) ? ( bv_8_180_n224 ) : ( n4911 ) ;
assign n4913 =  ( n4315 ) ? ( bv_8_198_n221 ) : ( n4912 ) ;
assign n4914 =  ( n4313 ) ? ( bv_8_232_n96 ) : ( n4913 ) ;
assign n4915 =  ( n4311 ) ? ( bv_8_221_n136 ) : ( n4914 ) ;
assign n4916 =  ( n4309 ) ? ( bv_8_116_n211 ) : ( n4915 ) ;
assign n4917 =  ( n4307 ) ? ( bv_8_31_n207 ) : ( n4916 ) ;
assign n4918 =  ( n4305 ) ? ( bv_8_75_n203 ) : ( n4917 ) ;
assign n4919 =  ( n4303 ) ? ( bv_8_189_n199 ) : ( n4918 ) ;
assign n4920 =  ( n4301 ) ? ( bv_8_139_n195 ) : ( n4919 ) ;
assign n4921 =  ( n4299 ) ? ( bv_8_138_n192 ) : ( n4920 ) ;
assign n4922 =  ( n4297 ) ? ( bv_8_112_n188 ) : ( n4921 ) ;
assign n4923 =  ( n4295 ) ? ( bv_8_62_n184 ) : ( n4922 ) ;
assign n4924 =  ( n4293 ) ? ( bv_8_181_n180 ) : ( n4923 ) ;
assign n4925 =  ( n4291 ) ? ( bv_8_102_n176 ) : ( n4924 ) ;
assign n4926 =  ( n4289 ) ? ( bv_8_72_n172 ) : ( n4925 ) ;
assign n4927 =  ( n4287 ) ? ( bv_8_3_n168 ) : ( n4926 ) ;
assign n4928 =  ( n4285 ) ? ( bv_8_246_n41 ) : ( n4927 ) ;
assign n4929 =  ( n4283 ) ? ( bv_8_14_n161 ) : ( n4928 ) ;
assign n4930 =  ( n4281 ) ? ( bv_8_97_n157 ) : ( n4929 ) ;
assign n4931 =  ( n4279 ) ? ( bv_8_53_n153 ) : ( n4930 ) ;
assign n4932 =  ( n4277 ) ? ( bv_8_87_n150 ) : ( n4931 ) ;
assign n4933 =  ( n4275 ) ? ( bv_8_185_n146 ) : ( n4932 ) ;
assign n4934 =  ( n4273 ) ? ( bv_8_134_n142 ) : ( n4933 ) ;
assign n4935 =  ( n4271 ) ? ( bv_8_193_n138 ) : ( n4934 ) ;
assign n4936 =  ( n4269 ) ? ( bv_8_29_n134 ) : ( n4935 ) ;
assign n4937 =  ( n4267 ) ? ( bv_8_158_n130 ) : ( n4936 ) ;
assign n4938 =  ( n4265 ) ? ( bv_8_225_n123 ) : ( n4937 ) ;
assign n4939 =  ( n4263 ) ? ( bv_8_248_n33 ) : ( n4938 ) ;
assign n4940 =  ( n4261 ) ? ( bv_8_152_n121 ) : ( n4939 ) ;
assign n4941 =  ( n4259 ) ? ( bv_8_17_n117 ) : ( n4940 ) ;
assign n4942 =  ( n4257 ) ? ( bv_8_105_n113 ) : ( n4941 ) ;
assign n4943 =  ( n4255 ) ? ( bv_8_217_n109 ) : ( n4942 ) ;
assign n4944 =  ( n4253 ) ? ( bv_8_142_n105 ) : ( n4943 ) ;
assign n4945 =  ( n4251 ) ? ( bv_8_148_n102 ) : ( n4944 ) ;
assign n4946 =  ( n4249 ) ? ( bv_8_155_n98 ) : ( n4945 ) ;
assign n4947 =  ( n4247 ) ? ( bv_8_30_n94 ) : ( n4946 ) ;
assign n4948 =  ( n4245 ) ? ( bv_8_135_n91 ) : ( n4947 ) ;
assign n4949 =  ( n4243 ) ? ( bv_8_233_n87 ) : ( n4948 ) ;
assign n4950 =  ( n4241 ) ? ( bv_8_206_n83 ) : ( n4949 ) ;
assign n4951 =  ( n4239 ) ? ( bv_8_85_n79 ) : ( n4950 ) ;
assign n4952 =  ( n4237 ) ? ( bv_8_40_n75 ) : ( n4951 ) ;
assign n4953 =  ( n4235 ) ? ( bv_8_223_n71 ) : ( n4952 ) ;
assign n4954 =  ( n4233 ) ? ( bv_8_140_n67 ) : ( n4953 ) ;
assign n4955 =  ( n4231 ) ? ( bv_8_161_n63 ) : ( n4954 ) ;
assign n4956 =  ( n4229 ) ? ( bv_8_137_n59 ) : ( n4955 ) ;
assign n4957 =  ( n4227 ) ? ( bv_8_13_n55 ) : ( n4956 ) ;
assign n4958 =  ( n4225 ) ? ( bv_8_191_n51 ) : ( n4957 ) ;
assign n4959 =  ( n4223 ) ? ( bv_8_230_n47 ) : ( n4958 ) ;
assign n4960 =  ( n4221 ) ? ( bv_8_66_n43 ) : ( n4959 ) ;
assign n4961 =  ( n4219 ) ? ( bv_8_104_n39 ) : ( n4960 ) ;
assign n4962 =  ( n4217 ) ? ( bv_8_65_n35 ) : ( n4961 ) ;
assign n4963 =  ( n4215 ) ? ( bv_8_153_n31 ) : ( n4962 ) ;
assign n4964 =  ( n4213 ) ? ( bv_8_45_n27 ) : ( n4963 ) ;
assign n4965 =  ( n4211 ) ? ( bv_8_15_n23 ) : ( n4964 ) ;
assign n4966 =  ( n4209 ) ? ( bv_8_176_n19 ) : ( n4965 ) ;
assign n4967 =  ( n4207 ) ? ( bv_8_84_n15 ) : ( n4966 ) ;
assign n4968 =  ( n4205 ) ? ( bv_8_187_n11 ) : ( n4967 ) ;
assign n4969 =  ( n4203 ) ? ( bv_8_22_n7 ) : ( n4968 ) ;
assign n4970 =  ( n4201 ) ^ ( n4969 )  ;
assign n4971 =  { ( n4200 ) , ( n4970 ) }  ;
assign n4972 = in[111:104] ;
assign n4973 = in[7:0] ;
assign n4974 =  ( n4973 ) == ( bv_8_255_n5 )  ;
assign n4975 = in[7:0] ;
assign n4976 =  ( n4975 ) == ( bv_8_254_n9 )  ;
assign n4977 = in[7:0] ;
assign n4978 =  ( n4977 ) == ( bv_8_253_n13 )  ;
assign n4979 = in[7:0] ;
assign n4980 =  ( n4979 ) == ( bv_8_252_n17 )  ;
assign n4981 = in[7:0] ;
assign n4982 =  ( n4981 ) == ( bv_8_251_n21 )  ;
assign n4983 = in[7:0] ;
assign n4984 =  ( n4983 ) == ( bv_8_250_n25 )  ;
assign n4985 = in[7:0] ;
assign n4986 =  ( n4985 ) == ( bv_8_249_n29 )  ;
assign n4987 = in[7:0] ;
assign n4988 =  ( n4987 ) == ( bv_8_248_n33 )  ;
assign n4989 = in[7:0] ;
assign n4990 =  ( n4989 ) == ( bv_8_247_n37 )  ;
assign n4991 = in[7:0] ;
assign n4992 =  ( n4991 ) == ( bv_8_246_n41 )  ;
assign n4993 = in[7:0] ;
assign n4994 =  ( n4993 ) == ( bv_8_245_n45 )  ;
assign n4995 = in[7:0] ;
assign n4996 =  ( n4995 ) == ( bv_8_244_n49 )  ;
assign n4997 = in[7:0] ;
assign n4998 =  ( n4997 ) == ( bv_8_243_n53 )  ;
assign n4999 = in[7:0] ;
assign n5000 =  ( n4999 ) == ( bv_8_242_n57 )  ;
assign n5001 = in[7:0] ;
assign n5002 =  ( n5001 ) == ( bv_8_241_n61 )  ;
assign n5003 = in[7:0] ;
assign n5004 =  ( n5003 ) == ( bv_8_240_n65 )  ;
assign n5005 = in[7:0] ;
assign n5006 =  ( n5005 ) == ( bv_8_239_n69 )  ;
assign n5007 = in[7:0] ;
assign n5008 =  ( n5007 ) == ( bv_8_238_n73 )  ;
assign n5009 = in[7:0] ;
assign n5010 =  ( n5009 ) == ( bv_8_237_n77 )  ;
assign n5011 = in[7:0] ;
assign n5012 =  ( n5011 ) == ( bv_8_236_n81 )  ;
assign n5013 = in[7:0] ;
assign n5014 =  ( n5013 ) == ( bv_8_235_n85 )  ;
assign n5015 = in[7:0] ;
assign n5016 =  ( n5015 ) == ( bv_8_234_n89 )  ;
assign n5017 = in[7:0] ;
assign n5018 =  ( n5017 ) == ( bv_8_233_n87 )  ;
assign n5019 = in[7:0] ;
assign n5020 =  ( n5019 ) == ( bv_8_232_n96 )  ;
assign n5021 = in[7:0] ;
assign n5022 =  ( n5021 ) == ( bv_8_231_n100 )  ;
assign n5023 = in[7:0] ;
assign n5024 =  ( n5023 ) == ( bv_8_230_n47 )  ;
assign n5025 = in[7:0] ;
assign n5026 =  ( n5025 ) == ( bv_8_229_n107 )  ;
assign n5027 = in[7:0] ;
assign n5028 =  ( n5027 ) == ( bv_8_228_n111 )  ;
assign n5029 = in[7:0] ;
assign n5030 =  ( n5029 ) == ( bv_8_227_n115 )  ;
assign n5031 = in[7:0] ;
assign n5032 =  ( n5031 ) == ( bv_8_226_n119 )  ;
assign n5033 = in[7:0] ;
assign n5034 =  ( n5033 ) == ( bv_8_225_n123 )  ;
assign n5035 = in[7:0] ;
assign n5036 =  ( n5035 ) == ( bv_8_224_n126 )  ;
assign n5037 = in[7:0] ;
assign n5038 =  ( n5037 ) == ( bv_8_223_n71 )  ;
assign n5039 = in[7:0] ;
assign n5040 =  ( n5039 ) == ( bv_8_222_n132 )  ;
assign n5041 = in[7:0] ;
assign n5042 =  ( n5041 ) == ( bv_8_221_n136 )  ;
assign n5043 = in[7:0] ;
assign n5044 =  ( n5043 ) == ( bv_8_220_n140 )  ;
assign n5045 = in[7:0] ;
assign n5046 =  ( n5045 ) == ( bv_8_219_n144 )  ;
assign n5047 = in[7:0] ;
assign n5048 =  ( n5047 ) == ( bv_8_218_n148 )  ;
assign n5049 = in[7:0] ;
assign n5050 =  ( n5049 ) == ( bv_8_217_n109 )  ;
assign n5051 = in[7:0] ;
assign n5052 =  ( n5051 ) == ( bv_8_216_n155 )  ;
assign n5053 = in[7:0] ;
assign n5054 =  ( n5053 ) == ( bv_8_215_n159 )  ;
assign n5055 = in[7:0] ;
assign n5056 =  ( n5055 ) == ( bv_8_214_n163 )  ;
assign n5057 = in[7:0] ;
assign n5058 =  ( n5057 ) == ( bv_8_213_n166 )  ;
assign n5059 = in[7:0] ;
assign n5060 =  ( n5059 ) == ( bv_8_212_n170 )  ;
assign n5061 = in[7:0] ;
assign n5062 =  ( n5061 ) == ( bv_8_211_n174 )  ;
assign n5063 = in[7:0] ;
assign n5064 =  ( n5063 ) == ( bv_8_210_n178 )  ;
assign n5065 = in[7:0] ;
assign n5066 =  ( n5065 ) == ( bv_8_209_n182 )  ;
assign n5067 = in[7:0] ;
assign n5068 =  ( n5067 ) == ( bv_8_208_n186 )  ;
assign n5069 = in[7:0] ;
assign n5070 =  ( n5069 ) == ( bv_8_207_n190 )  ;
assign n5071 = in[7:0] ;
assign n5072 =  ( n5071 ) == ( bv_8_206_n83 )  ;
assign n5073 = in[7:0] ;
assign n5074 =  ( n5073 ) == ( bv_8_205_n197 )  ;
assign n5075 = in[7:0] ;
assign n5076 =  ( n5075 ) == ( bv_8_204_n201 )  ;
assign n5077 = in[7:0] ;
assign n5078 =  ( n5077 ) == ( bv_8_203_n205 )  ;
assign n5079 = in[7:0] ;
assign n5080 =  ( n5079 ) == ( bv_8_202_n209 )  ;
assign n5081 = in[7:0] ;
assign n5082 =  ( n5081 ) == ( bv_8_201_n213 )  ;
assign n5083 = in[7:0] ;
assign n5084 =  ( n5083 ) == ( bv_8_200_n216 )  ;
assign n5085 = in[7:0] ;
assign n5086 =  ( n5085 ) == ( bv_8_199_n219 )  ;
assign n5087 = in[7:0] ;
assign n5088 =  ( n5087 ) == ( bv_8_198_n221 )  ;
assign n5089 = in[7:0] ;
assign n5090 =  ( n5089 ) == ( bv_8_197_n226 )  ;
assign n5091 = in[7:0] ;
assign n5092 =  ( n5091 ) == ( bv_8_196_n230 )  ;
assign n5093 = in[7:0] ;
assign n5094 =  ( n5093 ) == ( bv_8_195_n234 )  ;
assign n5095 = in[7:0] ;
assign n5096 =  ( n5095 ) == ( bv_8_194_n238 )  ;
assign n5097 = in[7:0] ;
assign n5098 =  ( n5097 ) == ( bv_8_193_n138 )  ;
assign n5099 = in[7:0] ;
assign n5100 =  ( n5099 ) == ( bv_8_192_n245 )  ;
assign n5101 = in[7:0] ;
assign n5102 =  ( n5101 ) == ( bv_8_191_n51 )  ;
assign n5103 = in[7:0] ;
assign n5104 =  ( n5103 ) == ( bv_8_190_n252 )  ;
assign n5105 = in[7:0] ;
assign n5106 =  ( n5105 ) == ( bv_8_189_n199 )  ;
assign n5107 = in[7:0] ;
assign n5108 =  ( n5107 ) == ( bv_8_188_n259 )  ;
assign n5109 = in[7:0] ;
assign n5110 =  ( n5109 ) == ( bv_8_187_n11 )  ;
assign n5111 = in[7:0] ;
assign n5112 =  ( n5111 ) == ( bv_8_186_n247 )  ;
assign n5113 = in[7:0] ;
assign n5114 =  ( n5113 ) == ( bv_8_185_n146 )  ;
assign n5115 = in[7:0] ;
assign n5116 =  ( n5115 ) == ( bv_8_184_n270 )  ;
assign n5117 = in[7:0] ;
assign n5118 =  ( n5117 ) == ( bv_8_183_n274 )  ;
assign n5119 = in[7:0] ;
assign n5120 =  ( n5119 ) == ( bv_8_182_n278 )  ;
assign n5121 = in[7:0] ;
assign n5122 =  ( n5121 ) == ( bv_8_181_n180 )  ;
assign n5123 = in[7:0] ;
assign n5124 =  ( n5123 ) == ( bv_8_180_n224 )  ;
assign n5125 = in[7:0] ;
assign n5126 =  ( n5125 ) == ( bv_8_179_n287 )  ;
assign n5127 = in[7:0] ;
assign n5128 =  ( n5127 ) == ( bv_8_178_n291 )  ;
assign n5129 = in[7:0] ;
assign n5130 =  ( n5129 ) == ( bv_8_177_n295 )  ;
assign n5131 = in[7:0] ;
assign n5132 =  ( n5131 ) == ( bv_8_176_n19 )  ;
assign n5133 = in[7:0] ;
assign n5134 =  ( n5133 ) == ( bv_8_175_n300 )  ;
assign n5135 = in[7:0] ;
assign n5136 =  ( n5135 ) == ( bv_8_174_n254 )  ;
assign n5137 = in[7:0] ;
assign n5138 =  ( n5137 ) == ( bv_8_173_n306 )  ;
assign n5139 = in[7:0] ;
assign n5140 =  ( n5139 ) == ( bv_8_172_n310 )  ;
assign n5141 = in[7:0] ;
assign n5142 =  ( n5141 ) == ( bv_8_171_n314 )  ;
assign n5143 = in[7:0] ;
assign n5144 =  ( n5143 ) == ( bv_8_170_n318 )  ;
assign n5145 = in[7:0] ;
assign n5146 =  ( n5145 ) == ( bv_8_169_n276 )  ;
assign n5147 = in[7:0] ;
assign n5148 =  ( n5147 ) == ( bv_8_168_n323 )  ;
assign n5149 = in[7:0] ;
assign n5150 =  ( n5149 ) == ( bv_8_167_n326 )  ;
assign n5151 = in[7:0] ;
assign n5152 =  ( n5151 ) == ( bv_8_166_n228 )  ;
assign n5153 = in[7:0] ;
assign n5154 =  ( n5153 ) == ( bv_8_165_n333 )  ;
assign n5155 = in[7:0] ;
assign n5156 =  ( n5155 ) == ( bv_8_164_n337 )  ;
assign n5157 = in[7:0] ;
assign n5158 =  ( n5157 ) == ( bv_8_163_n341 )  ;
assign n5159 = in[7:0] ;
assign n5160 =  ( n5159 ) == ( bv_8_162_n345 )  ;
assign n5161 = in[7:0] ;
assign n5162 =  ( n5161 ) == ( bv_8_161_n63 )  ;
assign n5163 = in[7:0] ;
assign n5164 =  ( n5163 ) == ( bv_8_160_n352 )  ;
assign n5165 = in[7:0] ;
assign n5166 =  ( n5165 ) == ( bv_8_159_n355 )  ;
assign n5167 = in[7:0] ;
assign n5168 =  ( n5167 ) == ( bv_8_158_n130 )  ;
assign n5169 = in[7:0] ;
assign n5170 =  ( n5169 ) == ( bv_8_157_n361 )  ;
assign n5171 = in[7:0] ;
assign n5172 =  ( n5171 ) == ( bv_8_156_n365 )  ;
assign n5173 = in[7:0] ;
assign n5174 =  ( n5173 ) == ( bv_8_155_n98 )  ;
assign n5175 = in[7:0] ;
assign n5176 =  ( n5175 ) == ( bv_8_154_n371 )  ;
assign n5177 = in[7:0] ;
assign n5178 =  ( n5177 ) == ( bv_8_153_n31 )  ;
assign n5179 = in[7:0] ;
assign n5180 =  ( n5179 ) == ( bv_8_152_n121 )  ;
assign n5181 = in[7:0] ;
assign n5182 =  ( n5181 ) == ( bv_8_151_n379 )  ;
assign n5183 = in[7:0] ;
assign n5184 =  ( n5183 ) == ( bv_8_150_n383 )  ;
assign n5185 = in[7:0] ;
assign n5186 =  ( n5185 ) == ( bv_8_149_n308 )  ;
assign n5187 = in[7:0] ;
assign n5188 =  ( n5187 ) == ( bv_8_148_n102 )  ;
assign n5189 = in[7:0] ;
assign n5190 =  ( n5189 ) == ( bv_8_147_n393 )  ;
assign n5191 = in[7:0] ;
assign n5192 =  ( n5191 ) == ( bv_8_146_n396 )  ;
assign n5193 = in[7:0] ;
assign n5194 =  ( n5193 ) == ( bv_8_145_n312 )  ;
assign n5195 = in[7:0] ;
assign n5196 =  ( n5195 ) == ( bv_8_144_n385 )  ;
assign n5197 = in[7:0] ;
assign n5198 =  ( n5197 ) == ( bv_8_143_n406 )  ;
assign n5199 = in[7:0] ;
assign n5200 =  ( n5199 ) == ( bv_8_142_n105 )  ;
assign n5201 = in[7:0] ;
assign n5202 =  ( n5201 ) == ( bv_8_141_n285 )  ;
assign n5203 = in[7:0] ;
assign n5204 =  ( n5203 ) == ( bv_8_140_n67 )  ;
assign n5205 = in[7:0] ;
assign n5206 =  ( n5205 ) == ( bv_8_139_n195 )  ;
assign n5207 = in[7:0] ;
assign n5208 =  ( n5207 ) == ( bv_8_138_n192 )  ;
assign n5209 = in[7:0] ;
assign n5210 =  ( n5209 ) == ( bv_8_137_n59 )  ;
assign n5211 = in[7:0] ;
assign n5212 =  ( n5211 ) == ( bv_8_136_n381 )  ;
assign n5213 = in[7:0] ;
assign n5214 =  ( n5213 ) == ( bv_8_135_n91 )  ;
assign n5215 = in[7:0] ;
assign n5216 =  ( n5215 ) == ( bv_8_134_n142 )  ;
assign n5217 = in[7:0] ;
assign n5218 =  ( n5217 ) == ( bv_8_133_n435 )  ;
assign n5219 = in[7:0] ;
assign n5220 =  ( n5219 ) == ( bv_8_132_n438 )  ;
assign n5221 = in[7:0] ;
assign n5222 =  ( n5221 ) == ( bv_8_131_n442 )  ;
assign n5223 = in[7:0] ;
assign n5224 =  ( n5223 ) == ( bv_8_130_n445 )  ;
assign n5225 = in[7:0] ;
assign n5226 =  ( n5225 ) == ( bv_8_129_n401 )  ;
assign n5227 = in[7:0] ;
assign n5228 =  ( n5227 ) == ( bv_8_128_n452 )  ;
assign n5229 = in[7:0] ;
assign n5230 =  ( n5229 ) == ( bv_8_127_n455 )  ;
assign n5231 = in[7:0] ;
assign n5232 =  ( n5231 ) == ( bv_8_126_n423 )  ;
assign n5233 = in[7:0] ;
assign n5234 =  ( n5233 ) == ( bv_8_125_n460 )  ;
assign n5235 = in[7:0] ;
assign n5236 =  ( n5235 ) == ( bv_8_124_n463 )  ;
assign n5237 = in[7:0] ;
assign n5238 =  ( n5237 ) == ( bv_8_123_n467 )  ;
assign n5239 = in[7:0] ;
assign n5240 =  ( n5239 ) == ( bv_8_122_n257 )  ;
assign n5241 = in[7:0] ;
assign n5242 =  ( n5241 ) == ( bv_8_121_n302 )  ;
assign n5243 = in[7:0] ;
assign n5244 =  ( n5243 ) == ( bv_8_120_n243 )  ;
assign n5245 = in[7:0] ;
assign n5246 =  ( n5245 ) == ( bv_8_119_n477 )  ;
assign n5247 = in[7:0] ;
assign n5248 =  ( n5247 ) == ( bv_8_118_n480 )  ;
assign n5249 = in[7:0] ;
assign n5250 =  ( n5249 ) == ( bv_8_117_n484 )  ;
assign n5251 = in[7:0] ;
assign n5252 =  ( n5251 ) == ( bv_8_116_n211 )  ;
assign n5253 = in[7:0] ;
assign n5254 =  ( n5253 ) == ( bv_8_115_n408 )  ;
assign n5255 = in[7:0] ;
assign n5256 =  ( n5255 ) == ( bv_8_114_n491 )  ;
assign n5257 = in[7:0] ;
assign n5258 =  ( n5257 ) == ( bv_8_113_n495 )  ;
assign n5259 = in[7:0] ;
assign n5260 =  ( n5259 ) == ( bv_8_112_n188 )  ;
assign n5261 = in[7:0] ;
assign n5262 =  ( n5261 ) == ( bv_8_111_n501 )  ;
assign n5263 = in[7:0] ;
assign n5264 =  ( n5263 ) == ( bv_8_110_n504 )  ;
assign n5265 = in[7:0] ;
assign n5266 =  ( n5265 ) == ( bv_8_109_n289 )  ;
assign n5267 = in[7:0] ;
assign n5268 =  ( n5267 ) == ( bv_8_108_n272 )  ;
assign n5269 = in[7:0] ;
assign n5270 =  ( n5269 ) == ( bv_8_107_n513 )  ;
assign n5271 = in[7:0] ;
assign n5272 =  ( n5271 ) == ( bv_8_106_n516 )  ;
assign n5273 = in[7:0] ;
assign n5274 =  ( n5273 ) == ( bv_8_105_n113 )  ;
assign n5275 = in[7:0] ;
assign n5276 =  ( n5275 ) == ( bv_8_104_n39 )  ;
assign n5277 = in[7:0] ;
assign n5278 =  ( n5277 ) == ( bv_8_103_n525 )  ;
assign n5279 = in[7:0] ;
assign n5280 =  ( n5279 ) == ( bv_8_102_n176 )  ;
assign n5281 = in[7:0] ;
assign n5282 =  ( n5281 ) == ( bv_8_101_n261 )  ;
assign n5283 = in[7:0] ;
assign n5284 =  ( n5283 ) == ( bv_8_100_n417 )  ;
assign n5285 = in[7:0] ;
assign n5286 =  ( n5285 ) == ( bv_8_99_n537 )  ;
assign n5287 = in[7:0] ;
assign n5288 =  ( n5287 ) == ( bv_8_98_n316 )  ;
assign n5289 = in[7:0] ;
assign n5290 =  ( n5289 ) == ( bv_8_97_n157 )  ;
assign n5291 = in[7:0] ;
assign n5292 =  ( n5291 ) == ( bv_8_96_n404 )  ;
assign n5293 = in[7:0] ;
assign n5294 =  ( n5293 ) == ( bv_8_95_n440 )  ;
assign n5295 = in[7:0] ;
assign n5296 =  ( n5295 ) == ( bv_8_94_n363 )  ;
assign n5297 = in[7:0] ;
assign n5298 =  ( n5297 ) == ( bv_8_93_n414 )  ;
assign n5299 = in[7:0] ;
assign n5300 =  ( n5299 ) == ( bv_8_92_n328 )  ;
assign n5301 = in[7:0] ;
assign n5302 =  ( n5301 ) == ( bv_8_91_n557 )  ;
assign n5303 = in[7:0] ;
assign n5304 =  ( n5303 ) == ( bv_8_90_n561 )  ;
assign n5305 = in[7:0] ;
assign n5306 =  ( n5305 ) == ( bv_8_89_n564 )  ;
assign n5307 = in[7:0] ;
assign n5308 =  ( n5307 ) == ( bv_8_88_n549 )  ;
assign n5309 = in[7:0] ;
assign n5310 =  ( n5309 ) == ( bv_8_87_n150 )  ;
assign n5311 = in[7:0] ;
assign n5312 =  ( n5311 ) == ( bv_8_86_n268 )  ;
assign n5313 = in[7:0] ;
assign n5314 =  ( n5313 ) == ( bv_8_85_n79 )  ;
assign n5315 = in[7:0] ;
assign n5316 =  ( n5315 ) == ( bv_8_84_n15 )  ;
assign n5317 = in[7:0] ;
assign n5318 =  ( n5317 ) == ( bv_8_83_n578 )  ;
assign n5319 = in[7:0] ;
assign n5320 =  ( n5319 ) == ( bv_8_82_n581 )  ;
assign n5321 = in[7:0] ;
assign n5322 =  ( n5321 ) == ( bv_8_81_n499 )  ;
assign n5323 = in[7:0] ;
assign n5324 =  ( n5323 ) == ( bv_8_80_n511 )  ;
assign n5325 = in[7:0] ;
assign n5326 =  ( n5325 ) == ( bv_8_79_n398 )  ;
assign n5327 = in[7:0] ;
assign n5328 =  ( n5327 ) == ( bv_8_78_n280 )  ;
assign n5329 = in[7:0] ;
assign n5330 =  ( n5329 ) == ( bv_8_77_n532 )  ;
assign n5331 = in[7:0] ;
assign n5332 =  ( n5331 ) == ( bv_8_76_n552 )  ;
assign n5333 = in[7:0] ;
assign n5334 =  ( n5333 ) == ( bv_8_75_n203 )  ;
assign n5335 = in[7:0] ;
assign n5336 =  ( n5335 ) == ( bv_8_74_n555 )  ;
assign n5337 = in[7:0] ;
assign n5338 =  ( n5337 ) == ( bv_8_73_n339 )  ;
assign n5339 = in[7:0] ;
assign n5340 =  ( n5339 ) == ( bv_8_72_n172 )  ;
assign n5341 = in[7:0] ;
assign n5342 =  ( n5341 ) == ( bv_8_71_n608 )  ;
assign n5343 = in[7:0] ;
assign n5344 =  ( n5343 ) == ( bv_8_70_n377 )  ;
assign n5345 = in[7:0] ;
assign n5346 =  ( n5345 ) == ( bv_8_69_n523 )  ;
assign n5347 = in[7:0] ;
assign n5348 =  ( n5347 ) == ( bv_8_68_n433 )  ;
assign n5349 = in[7:0] ;
assign n5350 =  ( n5349 ) == ( bv_8_67_n535 )  ;
assign n5351 = in[7:0] ;
assign n5352 =  ( n5351 ) == ( bv_8_66_n43 )  ;
assign n5353 = in[7:0] ;
assign n5354 =  ( n5353 ) == ( bv_8_65_n35 )  ;
assign n5355 = in[7:0] ;
assign n5356 =  ( n5355 ) == ( bv_8_64_n493 )  ;
assign n5357 = in[7:0] ;
assign n5358 =  ( n5357 ) == ( bv_8_63_n629 )  ;
assign n5359 = in[7:0] ;
assign n5360 =  ( n5359 ) == ( bv_8_62_n184 )  ;
assign n5361 = in[7:0] ;
assign n5362 =  ( n5361 ) == ( bv_8_61_n420 )  ;
assign n5363 = in[7:0] ;
assign n5364 =  ( n5363 ) == ( bv_8_60_n508 )  ;
assign n5365 = in[7:0] ;
assign n5366 =  ( n5365 ) == ( bv_8_59_n604 )  ;
assign n5367 = in[7:0] ;
assign n5368 =  ( n5367 ) == ( bv_8_58_n347 )  ;
assign n5369 = in[7:0] ;
assign n5370 =  ( n5369 ) == ( bv_8_57_n559 )  ;
assign n5371 = in[7:0] ;
assign n5372 =  ( n5371 ) == ( bv_8_56_n482 )  ;
assign n5373 = in[7:0] ;
assign n5374 =  ( n5373 ) == ( bv_8_55_n293 )  ;
assign n5375 = in[7:0] ;
assign n5376 =  ( n5375 ) == ( bv_8_54_n651 )  ;
assign n5377 = in[7:0] ;
assign n5378 =  ( n5377 ) == ( bv_8_53_n153 )  ;
assign n5379 = in[7:0] ;
assign n5380 =  ( n5379 ) == ( bv_8_52_n657 )  ;
assign n5381 = in[7:0] ;
assign n5382 =  ( n5381 ) == ( bv_8_51_n529 )  ;
assign n5383 = in[7:0] ;
assign n5384 =  ( n5383 ) == ( bv_8_50_n350 )  ;
assign n5385 = in[7:0] ;
assign n5386 =  ( n5385 ) == ( bv_8_49_n666 )  ;
assign n5387 = in[7:0] ;
assign n5388 =  ( n5387 ) == ( bv_8_48_n669 )  ;
assign n5389 = in[7:0] ;
assign n5390 =  ( n5389 ) == ( bv_8_47_n592 )  ;
assign n5391 = in[7:0] ;
assign n5392 =  ( n5391 ) == ( bv_8_46_n236 )  ;
assign n5393 = in[7:0] ;
assign n5394 =  ( n5393 ) == ( bv_8_45_n27 )  ;
assign n5395 = in[7:0] ;
assign n5396 =  ( n5395 ) == ( bv_8_44_n622 )  ;
assign n5397 = in[7:0] ;
assign n5398 =  ( n5397 ) == ( bv_8_43_n682 )  ;
assign n5399 = in[7:0] ;
assign n5400 =  ( n5399 ) == ( bv_8_42_n388 )  ;
assign n5401 = in[7:0] ;
assign n5402 =  ( n5401 ) == ( bv_8_41_n597 )  ;
assign n5403 = in[7:0] ;
assign n5404 =  ( n5403 ) == ( bv_8_40_n75 )  ;
assign n5405 = in[7:0] ;
assign n5406 =  ( n5405 ) == ( bv_8_39_n635 )  ;
assign n5407 = in[7:0] ;
assign n5408 =  ( n5407 ) == ( bv_8_38_n693 )  ;
assign n5409 = in[7:0] ;
assign n5410 =  ( n5409 ) == ( bv_8_37_n240 )  ;
assign n5411 = in[7:0] ;
assign n5412 =  ( n5411 ) == ( bv_8_36_n331 )  ;
assign n5413 = in[7:0] ;
assign n5414 =  ( n5413 ) == ( bv_8_35_n664 )  ;
assign n5415 = in[7:0] ;
assign n5416 =  ( n5415 ) == ( bv_8_34_n391 )  ;
assign n5417 = in[7:0] ;
assign n5418 =  ( n5417 ) == ( bv_8_33_n469 )  ;
assign n5419 = in[7:0] ;
assign n5420 =  ( n5419 ) == ( bv_8_32_n576 )  ;
assign n5421 = in[7:0] ;
assign n5422 =  ( n5421 ) == ( bv_8_31_n207 )  ;
assign n5423 = in[7:0] ;
assign n5424 =  ( n5423 ) == ( bv_8_30_n94 )  ;
assign n5425 = in[7:0] ;
assign n5426 =  ( n5425 ) == ( bv_8_29_n134 )  ;
assign n5427 = in[7:0] ;
assign n5428 =  ( n5427 ) == ( bv_8_28_n232 )  ;
assign n5429 = in[7:0] ;
assign n5430 =  ( n5429 ) == ( bv_8_27_n616 )  ;
assign n5431 = in[7:0] ;
assign n5432 =  ( n5431 ) == ( bv_8_26_n619 )  ;
assign n5433 = in[7:0] ;
assign n5434 =  ( n5433 ) == ( bv_8_25_n411 )  ;
assign n5435 = in[7:0] ;
assign n5436 =  ( n5435 ) == ( bv_8_24_n659 )  ;
assign n5437 = in[7:0] ;
assign n5438 =  ( n5437 ) == ( bv_8_23_n430 )  ;
assign n5439 = in[7:0] ;
assign n5440 =  ( n5439 ) == ( bv_8_22_n7 )  ;
assign n5441 = in[7:0] ;
assign n5442 =  ( n5441 ) == ( bv_8_21_n674 )  ;
assign n5443 = in[7:0] ;
assign n5444 =  ( n5443 ) == ( bv_8_20_n369 )  ;
assign n5445 = in[7:0] ;
assign n5446 =  ( n5445 ) == ( bv_8_19_n447 )  ;
assign n5447 = in[7:0] ;
assign n5448 =  ( n5447 ) == ( bv_8_18_n644 )  ;
assign n5449 = in[7:0] ;
assign n5450 =  ( n5449 ) == ( bv_8_17_n117 )  ;
assign n5451 = in[7:0] ;
assign n5452 =  ( n5451 ) == ( bv_8_16_n465 )  ;
assign n5453 = in[7:0] ;
assign n5454 =  ( n5453 ) == ( bv_8_15_n23 )  ;
assign n5455 = in[7:0] ;
assign n5456 =  ( n5455 ) == ( bv_8_14_n161 )  ;
assign n5457 = in[7:0] ;
assign n5458 =  ( n5457 ) == ( bv_8_13_n55 )  ;
assign n5459 = in[7:0] ;
assign n5460 =  ( n5459 ) == ( bv_8_12_n450 )  ;
assign n5461 = in[7:0] ;
assign n5462 =  ( n5461 ) == ( bv_8_11_n359 )  ;
assign n5463 = in[7:0] ;
assign n5464 =  ( n5463 ) == ( bv_8_10_n343 )  ;
assign n5465 = in[7:0] ;
assign n5466 =  ( n5465 ) == ( bv_8_9_n627 )  ;
assign n5467 = in[7:0] ;
assign n5468 =  ( n5467 ) == ( bv_8_8_n250 )  ;
assign n5469 = in[7:0] ;
assign n5470 =  ( n5469 ) == ( bv_8_7_n647 )  ;
assign n5471 = in[7:0] ;
assign n5472 =  ( n5471 ) == ( bv_8_6_n335 )  ;
assign n5473 = in[7:0] ;
assign n5474 =  ( n5473 ) == ( bv_8_5_n653 )  ;
assign n5475 = in[7:0] ;
assign n5476 =  ( n5475 ) == ( bv_8_4_n671 )  ;
assign n5477 = in[7:0] ;
assign n5478 =  ( n5477 ) == ( bv_8_3_n168 )  ;
assign n5479 = in[7:0] ;
assign n5480 =  ( n5479 ) == ( bv_8_2_n518 )  ;
assign n5481 = in[7:0] ;
assign n5482 =  ( n5481 ) == ( bv_8_1_n753 )  ;
assign n5483 = in[7:0] ;
assign n5484 =  ( n5483 ) == ( bv_8_0_n583 )  ;
assign n5485 =  ( n5484 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n5486 =  ( n5482 ) ? ( bv_8_124_n463 ) : ( n5485 ) ;
assign n5487 =  ( n5480 ) ? ( bv_8_119_n477 ) : ( n5486 ) ;
assign n5488 =  ( n5478 ) ? ( bv_8_123_n467 ) : ( n5487 ) ;
assign n5489 =  ( n5476 ) ? ( bv_8_242_n57 ) : ( n5488 ) ;
assign n5490 =  ( n5474 ) ? ( bv_8_107_n513 ) : ( n5489 ) ;
assign n5491 =  ( n5472 ) ? ( bv_8_111_n501 ) : ( n5490 ) ;
assign n5492 =  ( n5470 ) ? ( bv_8_197_n226 ) : ( n5491 ) ;
assign n5493 =  ( n5468 ) ? ( bv_8_48_n669 ) : ( n5492 ) ;
assign n5494 =  ( n5466 ) ? ( bv_8_1_n753 ) : ( n5493 ) ;
assign n5495 =  ( n5464 ) ? ( bv_8_103_n525 ) : ( n5494 ) ;
assign n5496 =  ( n5462 ) ? ( bv_8_43_n682 ) : ( n5495 ) ;
assign n5497 =  ( n5460 ) ? ( bv_8_254_n9 ) : ( n5496 ) ;
assign n5498 =  ( n5458 ) ? ( bv_8_215_n159 ) : ( n5497 ) ;
assign n5499 =  ( n5456 ) ? ( bv_8_171_n314 ) : ( n5498 ) ;
assign n5500 =  ( n5454 ) ? ( bv_8_118_n480 ) : ( n5499 ) ;
assign n5501 =  ( n5452 ) ? ( bv_8_202_n209 ) : ( n5500 ) ;
assign n5502 =  ( n5450 ) ? ( bv_8_130_n445 ) : ( n5501 ) ;
assign n5503 =  ( n5448 ) ? ( bv_8_201_n213 ) : ( n5502 ) ;
assign n5504 =  ( n5446 ) ? ( bv_8_125_n460 ) : ( n5503 ) ;
assign n5505 =  ( n5444 ) ? ( bv_8_250_n25 ) : ( n5504 ) ;
assign n5506 =  ( n5442 ) ? ( bv_8_89_n564 ) : ( n5505 ) ;
assign n5507 =  ( n5440 ) ? ( bv_8_71_n608 ) : ( n5506 ) ;
assign n5508 =  ( n5438 ) ? ( bv_8_240_n65 ) : ( n5507 ) ;
assign n5509 =  ( n5436 ) ? ( bv_8_173_n306 ) : ( n5508 ) ;
assign n5510 =  ( n5434 ) ? ( bv_8_212_n170 ) : ( n5509 ) ;
assign n5511 =  ( n5432 ) ? ( bv_8_162_n345 ) : ( n5510 ) ;
assign n5512 =  ( n5430 ) ? ( bv_8_175_n300 ) : ( n5511 ) ;
assign n5513 =  ( n5428 ) ? ( bv_8_156_n365 ) : ( n5512 ) ;
assign n5514 =  ( n5426 ) ? ( bv_8_164_n337 ) : ( n5513 ) ;
assign n5515 =  ( n5424 ) ? ( bv_8_114_n491 ) : ( n5514 ) ;
assign n5516 =  ( n5422 ) ? ( bv_8_192_n245 ) : ( n5515 ) ;
assign n5517 =  ( n5420 ) ? ( bv_8_183_n274 ) : ( n5516 ) ;
assign n5518 =  ( n5418 ) ? ( bv_8_253_n13 ) : ( n5517 ) ;
assign n5519 =  ( n5416 ) ? ( bv_8_147_n393 ) : ( n5518 ) ;
assign n5520 =  ( n5414 ) ? ( bv_8_38_n693 ) : ( n5519 ) ;
assign n5521 =  ( n5412 ) ? ( bv_8_54_n651 ) : ( n5520 ) ;
assign n5522 =  ( n5410 ) ? ( bv_8_63_n629 ) : ( n5521 ) ;
assign n5523 =  ( n5408 ) ? ( bv_8_247_n37 ) : ( n5522 ) ;
assign n5524 =  ( n5406 ) ? ( bv_8_204_n201 ) : ( n5523 ) ;
assign n5525 =  ( n5404 ) ? ( bv_8_52_n657 ) : ( n5524 ) ;
assign n5526 =  ( n5402 ) ? ( bv_8_165_n333 ) : ( n5525 ) ;
assign n5527 =  ( n5400 ) ? ( bv_8_229_n107 ) : ( n5526 ) ;
assign n5528 =  ( n5398 ) ? ( bv_8_241_n61 ) : ( n5527 ) ;
assign n5529 =  ( n5396 ) ? ( bv_8_113_n495 ) : ( n5528 ) ;
assign n5530 =  ( n5394 ) ? ( bv_8_216_n155 ) : ( n5529 ) ;
assign n5531 =  ( n5392 ) ? ( bv_8_49_n666 ) : ( n5530 ) ;
assign n5532 =  ( n5390 ) ? ( bv_8_21_n674 ) : ( n5531 ) ;
assign n5533 =  ( n5388 ) ? ( bv_8_4_n671 ) : ( n5532 ) ;
assign n5534 =  ( n5386 ) ? ( bv_8_199_n219 ) : ( n5533 ) ;
assign n5535 =  ( n5384 ) ? ( bv_8_35_n664 ) : ( n5534 ) ;
assign n5536 =  ( n5382 ) ? ( bv_8_195_n234 ) : ( n5535 ) ;
assign n5537 =  ( n5380 ) ? ( bv_8_24_n659 ) : ( n5536 ) ;
assign n5538 =  ( n5378 ) ? ( bv_8_150_n383 ) : ( n5537 ) ;
assign n5539 =  ( n5376 ) ? ( bv_8_5_n653 ) : ( n5538 ) ;
assign n5540 =  ( n5374 ) ? ( bv_8_154_n371 ) : ( n5539 ) ;
assign n5541 =  ( n5372 ) ? ( bv_8_7_n647 ) : ( n5540 ) ;
assign n5542 =  ( n5370 ) ? ( bv_8_18_n644 ) : ( n5541 ) ;
assign n5543 =  ( n5368 ) ? ( bv_8_128_n452 ) : ( n5542 ) ;
assign n5544 =  ( n5366 ) ? ( bv_8_226_n119 ) : ( n5543 ) ;
assign n5545 =  ( n5364 ) ? ( bv_8_235_n85 ) : ( n5544 ) ;
assign n5546 =  ( n5362 ) ? ( bv_8_39_n635 ) : ( n5545 ) ;
assign n5547 =  ( n5360 ) ? ( bv_8_178_n291 ) : ( n5546 ) ;
assign n5548 =  ( n5358 ) ? ( bv_8_117_n484 ) : ( n5547 ) ;
assign n5549 =  ( n5356 ) ? ( bv_8_9_n627 ) : ( n5548 ) ;
assign n5550 =  ( n5354 ) ? ( bv_8_131_n442 ) : ( n5549 ) ;
assign n5551 =  ( n5352 ) ? ( bv_8_44_n622 ) : ( n5550 ) ;
assign n5552 =  ( n5350 ) ? ( bv_8_26_n619 ) : ( n5551 ) ;
assign n5553 =  ( n5348 ) ? ( bv_8_27_n616 ) : ( n5552 ) ;
assign n5554 =  ( n5346 ) ? ( bv_8_110_n504 ) : ( n5553 ) ;
assign n5555 =  ( n5344 ) ? ( bv_8_90_n561 ) : ( n5554 ) ;
assign n5556 =  ( n5342 ) ? ( bv_8_160_n352 ) : ( n5555 ) ;
assign n5557 =  ( n5340 ) ? ( bv_8_82_n581 ) : ( n5556 ) ;
assign n5558 =  ( n5338 ) ? ( bv_8_59_n604 ) : ( n5557 ) ;
assign n5559 =  ( n5336 ) ? ( bv_8_214_n163 ) : ( n5558 ) ;
assign n5560 =  ( n5334 ) ? ( bv_8_179_n287 ) : ( n5559 ) ;
assign n5561 =  ( n5332 ) ? ( bv_8_41_n597 ) : ( n5560 ) ;
assign n5562 =  ( n5330 ) ? ( bv_8_227_n115 ) : ( n5561 ) ;
assign n5563 =  ( n5328 ) ? ( bv_8_47_n592 ) : ( n5562 ) ;
assign n5564 =  ( n5326 ) ? ( bv_8_132_n438 ) : ( n5563 ) ;
assign n5565 =  ( n5324 ) ? ( bv_8_83_n578 ) : ( n5564 ) ;
assign n5566 =  ( n5322 ) ? ( bv_8_209_n182 ) : ( n5565 ) ;
assign n5567 =  ( n5320 ) ? ( bv_8_0_n583 ) : ( n5566 ) ;
assign n5568 =  ( n5318 ) ? ( bv_8_237_n77 ) : ( n5567 ) ;
assign n5569 =  ( n5316 ) ? ( bv_8_32_n576 ) : ( n5568 ) ;
assign n5570 =  ( n5314 ) ? ( bv_8_252_n17 ) : ( n5569 ) ;
assign n5571 =  ( n5312 ) ? ( bv_8_177_n295 ) : ( n5570 ) ;
assign n5572 =  ( n5310 ) ? ( bv_8_91_n557 ) : ( n5571 ) ;
assign n5573 =  ( n5308 ) ? ( bv_8_106_n516 ) : ( n5572 ) ;
assign n5574 =  ( n5306 ) ? ( bv_8_203_n205 ) : ( n5573 ) ;
assign n5575 =  ( n5304 ) ? ( bv_8_190_n252 ) : ( n5574 ) ;
assign n5576 =  ( n5302 ) ? ( bv_8_57_n559 ) : ( n5575 ) ;
assign n5577 =  ( n5300 ) ? ( bv_8_74_n555 ) : ( n5576 ) ;
assign n5578 =  ( n5298 ) ? ( bv_8_76_n552 ) : ( n5577 ) ;
assign n5579 =  ( n5296 ) ? ( bv_8_88_n549 ) : ( n5578 ) ;
assign n5580 =  ( n5294 ) ? ( bv_8_207_n190 ) : ( n5579 ) ;
assign n5581 =  ( n5292 ) ? ( bv_8_208_n186 ) : ( n5580 ) ;
assign n5582 =  ( n5290 ) ? ( bv_8_239_n69 ) : ( n5581 ) ;
assign n5583 =  ( n5288 ) ? ( bv_8_170_n318 ) : ( n5582 ) ;
assign n5584 =  ( n5286 ) ? ( bv_8_251_n21 ) : ( n5583 ) ;
assign n5585 =  ( n5284 ) ? ( bv_8_67_n535 ) : ( n5584 ) ;
assign n5586 =  ( n5282 ) ? ( bv_8_77_n532 ) : ( n5585 ) ;
assign n5587 =  ( n5280 ) ? ( bv_8_51_n529 ) : ( n5586 ) ;
assign n5588 =  ( n5278 ) ? ( bv_8_133_n435 ) : ( n5587 ) ;
assign n5589 =  ( n5276 ) ? ( bv_8_69_n523 ) : ( n5588 ) ;
assign n5590 =  ( n5274 ) ? ( bv_8_249_n29 ) : ( n5589 ) ;
assign n5591 =  ( n5272 ) ? ( bv_8_2_n518 ) : ( n5590 ) ;
assign n5592 =  ( n5270 ) ? ( bv_8_127_n455 ) : ( n5591 ) ;
assign n5593 =  ( n5268 ) ? ( bv_8_80_n511 ) : ( n5592 ) ;
assign n5594 =  ( n5266 ) ? ( bv_8_60_n508 ) : ( n5593 ) ;
assign n5595 =  ( n5264 ) ? ( bv_8_159_n355 ) : ( n5594 ) ;
assign n5596 =  ( n5262 ) ? ( bv_8_168_n323 ) : ( n5595 ) ;
assign n5597 =  ( n5260 ) ? ( bv_8_81_n499 ) : ( n5596 ) ;
assign n5598 =  ( n5258 ) ? ( bv_8_163_n341 ) : ( n5597 ) ;
assign n5599 =  ( n5256 ) ? ( bv_8_64_n493 ) : ( n5598 ) ;
assign n5600 =  ( n5254 ) ? ( bv_8_143_n406 ) : ( n5599 ) ;
assign n5601 =  ( n5252 ) ? ( bv_8_146_n396 ) : ( n5600 ) ;
assign n5602 =  ( n5250 ) ? ( bv_8_157_n361 ) : ( n5601 ) ;
assign n5603 =  ( n5248 ) ? ( bv_8_56_n482 ) : ( n5602 ) ;
assign n5604 =  ( n5246 ) ? ( bv_8_245_n45 ) : ( n5603 ) ;
assign n5605 =  ( n5244 ) ? ( bv_8_188_n259 ) : ( n5604 ) ;
assign n5606 =  ( n5242 ) ? ( bv_8_182_n278 ) : ( n5605 ) ;
assign n5607 =  ( n5240 ) ? ( bv_8_218_n148 ) : ( n5606 ) ;
assign n5608 =  ( n5238 ) ? ( bv_8_33_n469 ) : ( n5607 ) ;
assign n5609 =  ( n5236 ) ? ( bv_8_16_n465 ) : ( n5608 ) ;
assign n5610 =  ( n5234 ) ? ( bv_8_255_n5 ) : ( n5609 ) ;
assign n5611 =  ( n5232 ) ? ( bv_8_243_n53 ) : ( n5610 ) ;
assign n5612 =  ( n5230 ) ? ( bv_8_210_n178 ) : ( n5611 ) ;
assign n5613 =  ( n5228 ) ? ( bv_8_205_n197 ) : ( n5612 ) ;
assign n5614 =  ( n5226 ) ? ( bv_8_12_n450 ) : ( n5613 ) ;
assign n5615 =  ( n5224 ) ? ( bv_8_19_n447 ) : ( n5614 ) ;
assign n5616 =  ( n5222 ) ? ( bv_8_236_n81 ) : ( n5615 ) ;
assign n5617 =  ( n5220 ) ? ( bv_8_95_n440 ) : ( n5616 ) ;
assign n5618 =  ( n5218 ) ? ( bv_8_151_n379 ) : ( n5617 ) ;
assign n5619 =  ( n5216 ) ? ( bv_8_68_n433 ) : ( n5618 ) ;
assign n5620 =  ( n5214 ) ? ( bv_8_23_n430 ) : ( n5619 ) ;
assign n5621 =  ( n5212 ) ? ( bv_8_196_n230 ) : ( n5620 ) ;
assign n5622 =  ( n5210 ) ? ( bv_8_167_n326 ) : ( n5621 ) ;
assign n5623 =  ( n5208 ) ? ( bv_8_126_n423 ) : ( n5622 ) ;
assign n5624 =  ( n5206 ) ? ( bv_8_61_n420 ) : ( n5623 ) ;
assign n5625 =  ( n5204 ) ? ( bv_8_100_n417 ) : ( n5624 ) ;
assign n5626 =  ( n5202 ) ? ( bv_8_93_n414 ) : ( n5625 ) ;
assign n5627 =  ( n5200 ) ? ( bv_8_25_n411 ) : ( n5626 ) ;
assign n5628 =  ( n5198 ) ? ( bv_8_115_n408 ) : ( n5627 ) ;
assign n5629 =  ( n5196 ) ? ( bv_8_96_n404 ) : ( n5628 ) ;
assign n5630 =  ( n5194 ) ? ( bv_8_129_n401 ) : ( n5629 ) ;
assign n5631 =  ( n5192 ) ? ( bv_8_79_n398 ) : ( n5630 ) ;
assign n5632 =  ( n5190 ) ? ( bv_8_220_n140 ) : ( n5631 ) ;
assign n5633 =  ( n5188 ) ? ( bv_8_34_n391 ) : ( n5632 ) ;
assign n5634 =  ( n5186 ) ? ( bv_8_42_n388 ) : ( n5633 ) ;
assign n5635 =  ( n5184 ) ? ( bv_8_144_n385 ) : ( n5634 ) ;
assign n5636 =  ( n5182 ) ? ( bv_8_136_n381 ) : ( n5635 ) ;
assign n5637 =  ( n5180 ) ? ( bv_8_70_n377 ) : ( n5636 ) ;
assign n5638 =  ( n5178 ) ? ( bv_8_238_n73 ) : ( n5637 ) ;
assign n5639 =  ( n5176 ) ? ( bv_8_184_n270 ) : ( n5638 ) ;
assign n5640 =  ( n5174 ) ? ( bv_8_20_n369 ) : ( n5639 ) ;
assign n5641 =  ( n5172 ) ? ( bv_8_222_n132 ) : ( n5640 ) ;
assign n5642 =  ( n5170 ) ? ( bv_8_94_n363 ) : ( n5641 ) ;
assign n5643 =  ( n5168 ) ? ( bv_8_11_n359 ) : ( n5642 ) ;
assign n5644 =  ( n5166 ) ? ( bv_8_219_n144 ) : ( n5643 ) ;
assign n5645 =  ( n5164 ) ? ( bv_8_224_n126 ) : ( n5644 ) ;
assign n5646 =  ( n5162 ) ? ( bv_8_50_n350 ) : ( n5645 ) ;
assign n5647 =  ( n5160 ) ? ( bv_8_58_n347 ) : ( n5646 ) ;
assign n5648 =  ( n5158 ) ? ( bv_8_10_n343 ) : ( n5647 ) ;
assign n5649 =  ( n5156 ) ? ( bv_8_73_n339 ) : ( n5648 ) ;
assign n5650 =  ( n5154 ) ? ( bv_8_6_n335 ) : ( n5649 ) ;
assign n5651 =  ( n5152 ) ? ( bv_8_36_n331 ) : ( n5650 ) ;
assign n5652 =  ( n5150 ) ? ( bv_8_92_n328 ) : ( n5651 ) ;
assign n5653 =  ( n5148 ) ? ( bv_8_194_n238 ) : ( n5652 ) ;
assign n5654 =  ( n5146 ) ? ( bv_8_211_n174 ) : ( n5653 ) ;
assign n5655 =  ( n5144 ) ? ( bv_8_172_n310 ) : ( n5654 ) ;
assign n5656 =  ( n5142 ) ? ( bv_8_98_n316 ) : ( n5655 ) ;
assign n5657 =  ( n5140 ) ? ( bv_8_145_n312 ) : ( n5656 ) ;
assign n5658 =  ( n5138 ) ? ( bv_8_149_n308 ) : ( n5657 ) ;
assign n5659 =  ( n5136 ) ? ( bv_8_228_n111 ) : ( n5658 ) ;
assign n5660 =  ( n5134 ) ? ( bv_8_121_n302 ) : ( n5659 ) ;
assign n5661 =  ( n5132 ) ? ( bv_8_231_n100 ) : ( n5660 ) ;
assign n5662 =  ( n5130 ) ? ( bv_8_200_n216 ) : ( n5661 ) ;
assign n5663 =  ( n5128 ) ? ( bv_8_55_n293 ) : ( n5662 ) ;
assign n5664 =  ( n5126 ) ? ( bv_8_109_n289 ) : ( n5663 ) ;
assign n5665 =  ( n5124 ) ? ( bv_8_141_n285 ) : ( n5664 ) ;
assign n5666 =  ( n5122 ) ? ( bv_8_213_n166 ) : ( n5665 ) ;
assign n5667 =  ( n5120 ) ? ( bv_8_78_n280 ) : ( n5666 ) ;
assign n5668 =  ( n5118 ) ? ( bv_8_169_n276 ) : ( n5667 ) ;
assign n5669 =  ( n5116 ) ? ( bv_8_108_n272 ) : ( n5668 ) ;
assign n5670 =  ( n5114 ) ? ( bv_8_86_n268 ) : ( n5669 ) ;
assign n5671 =  ( n5112 ) ? ( bv_8_244_n49 ) : ( n5670 ) ;
assign n5672 =  ( n5110 ) ? ( bv_8_234_n89 ) : ( n5671 ) ;
assign n5673 =  ( n5108 ) ? ( bv_8_101_n261 ) : ( n5672 ) ;
assign n5674 =  ( n5106 ) ? ( bv_8_122_n257 ) : ( n5673 ) ;
assign n5675 =  ( n5104 ) ? ( bv_8_174_n254 ) : ( n5674 ) ;
assign n5676 =  ( n5102 ) ? ( bv_8_8_n250 ) : ( n5675 ) ;
assign n5677 =  ( n5100 ) ? ( bv_8_186_n247 ) : ( n5676 ) ;
assign n5678 =  ( n5098 ) ? ( bv_8_120_n243 ) : ( n5677 ) ;
assign n5679 =  ( n5096 ) ? ( bv_8_37_n240 ) : ( n5678 ) ;
assign n5680 =  ( n5094 ) ? ( bv_8_46_n236 ) : ( n5679 ) ;
assign n5681 =  ( n5092 ) ? ( bv_8_28_n232 ) : ( n5680 ) ;
assign n5682 =  ( n5090 ) ? ( bv_8_166_n228 ) : ( n5681 ) ;
assign n5683 =  ( n5088 ) ? ( bv_8_180_n224 ) : ( n5682 ) ;
assign n5684 =  ( n5086 ) ? ( bv_8_198_n221 ) : ( n5683 ) ;
assign n5685 =  ( n5084 ) ? ( bv_8_232_n96 ) : ( n5684 ) ;
assign n5686 =  ( n5082 ) ? ( bv_8_221_n136 ) : ( n5685 ) ;
assign n5687 =  ( n5080 ) ? ( bv_8_116_n211 ) : ( n5686 ) ;
assign n5688 =  ( n5078 ) ? ( bv_8_31_n207 ) : ( n5687 ) ;
assign n5689 =  ( n5076 ) ? ( bv_8_75_n203 ) : ( n5688 ) ;
assign n5690 =  ( n5074 ) ? ( bv_8_189_n199 ) : ( n5689 ) ;
assign n5691 =  ( n5072 ) ? ( bv_8_139_n195 ) : ( n5690 ) ;
assign n5692 =  ( n5070 ) ? ( bv_8_138_n192 ) : ( n5691 ) ;
assign n5693 =  ( n5068 ) ? ( bv_8_112_n188 ) : ( n5692 ) ;
assign n5694 =  ( n5066 ) ? ( bv_8_62_n184 ) : ( n5693 ) ;
assign n5695 =  ( n5064 ) ? ( bv_8_181_n180 ) : ( n5694 ) ;
assign n5696 =  ( n5062 ) ? ( bv_8_102_n176 ) : ( n5695 ) ;
assign n5697 =  ( n5060 ) ? ( bv_8_72_n172 ) : ( n5696 ) ;
assign n5698 =  ( n5058 ) ? ( bv_8_3_n168 ) : ( n5697 ) ;
assign n5699 =  ( n5056 ) ? ( bv_8_246_n41 ) : ( n5698 ) ;
assign n5700 =  ( n5054 ) ? ( bv_8_14_n161 ) : ( n5699 ) ;
assign n5701 =  ( n5052 ) ? ( bv_8_97_n157 ) : ( n5700 ) ;
assign n5702 =  ( n5050 ) ? ( bv_8_53_n153 ) : ( n5701 ) ;
assign n5703 =  ( n5048 ) ? ( bv_8_87_n150 ) : ( n5702 ) ;
assign n5704 =  ( n5046 ) ? ( bv_8_185_n146 ) : ( n5703 ) ;
assign n5705 =  ( n5044 ) ? ( bv_8_134_n142 ) : ( n5704 ) ;
assign n5706 =  ( n5042 ) ? ( bv_8_193_n138 ) : ( n5705 ) ;
assign n5707 =  ( n5040 ) ? ( bv_8_29_n134 ) : ( n5706 ) ;
assign n5708 =  ( n5038 ) ? ( bv_8_158_n130 ) : ( n5707 ) ;
assign n5709 =  ( n5036 ) ? ( bv_8_225_n123 ) : ( n5708 ) ;
assign n5710 =  ( n5034 ) ? ( bv_8_248_n33 ) : ( n5709 ) ;
assign n5711 =  ( n5032 ) ? ( bv_8_152_n121 ) : ( n5710 ) ;
assign n5712 =  ( n5030 ) ? ( bv_8_17_n117 ) : ( n5711 ) ;
assign n5713 =  ( n5028 ) ? ( bv_8_105_n113 ) : ( n5712 ) ;
assign n5714 =  ( n5026 ) ? ( bv_8_217_n109 ) : ( n5713 ) ;
assign n5715 =  ( n5024 ) ? ( bv_8_142_n105 ) : ( n5714 ) ;
assign n5716 =  ( n5022 ) ? ( bv_8_148_n102 ) : ( n5715 ) ;
assign n5717 =  ( n5020 ) ? ( bv_8_155_n98 ) : ( n5716 ) ;
assign n5718 =  ( n5018 ) ? ( bv_8_30_n94 ) : ( n5717 ) ;
assign n5719 =  ( n5016 ) ? ( bv_8_135_n91 ) : ( n5718 ) ;
assign n5720 =  ( n5014 ) ? ( bv_8_233_n87 ) : ( n5719 ) ;
assign n5721 =  ( n5012 ) ? ( bv_8_206_n83 ) : ( n5720 ) ;
assign n5722 =  ( n5010 ) ? ( bv_8_85_n79 ) : ( n5721 ) ;
assign n5723 =  ( n5008 ) ? ( bv_8_40_n75 ) : ( n5722 ) ;
assign n5724 =  ( n5006 ) ? ( bv_8_223_n71 ) : ( n5723 ) ;
assign n5725 =  ( n5004 ) ? ( bv_8_140_n67 ) : ( n5724 ) ;
assign n5726 =  ( n5002 ) ? ( bv_8_161_n63 ) : ( n5725 ) ;
assign n5727 =  ( n5000 ) ? ( bv_8_137_n59 ) : ( n5726 ) ;
assign n5728 =  ( n4998 ) ? ( bv_8_13_n55 ) : ( n5727 ) ;
assign n5729 =  ( n4996 ) ? ( bv_8_191_n51 ) : ( n5728 ) ;
assign n5730 =  ( n4994 ) ? ( bv_8_230_n47 ) : ( n5729 ) ;
assign n5731 =  ( n4992 ) ? ( bv_8_66_n43 ) : ( n5730 ) ;
assign n5732 =  ( n4990 ) ? ( bv_8_104_n39 ) : ( n5731 ) ;
assign n5733 =  ( n4988 ) ? ( bv_8_65_n35 ) : ( n5732 ) ;
assign n5734 =  ( n4986 ) ? ( bv_8_153_n31 ) : ( n5733 ) ;
assign n5735 =  ( n4984 ) ? ( bv_8_45_n27 ) : ( n5734 ) ;
assign n5736 =  ( n4982 ) ? ( bv_8_15_n23 ) : ( n5735 ) ;
assign n5737 =  ( n4980 ) ? ( bv_8_176_n19 ) : ( n5736 ) ;
assign n5738 =  ( n4978 ) ? ( bv_8_84_n15 ) : ( n5737 ) ;
assign n5739 =  ( n4976 ) ? ( bv_8_187_n11 ) : ( n5738 ) ;
assign n5740 =  ( n4974 ) ? ( bv_8_22_n7 ) : ( n5739 ) ;
assign n5741 =  ( n4972 ) ^ ( n5740 )  ;
assign n5742 =  { ( n4971 ) , ( n5741 ) }  ;
assign n5743 = in[103:96] ;
assign n5744 = in[31:24] ;
assign n5745 =  ( n5744 ) == ( bv_8_255_n5 )  ;
assign n5746 = in[31:24] ;
assign n5747 =  ( n5746 ) == ( bv_8_254_n9 )  ;
assign n5748 = in[31:24] ;
assign n5749 =  ( n5748 ) == ( bv_8_253_n13 )  ;
assign n5750 = in[31:24] ;
assign n5751 =  ( n5750 ) == ( bv_8_252_n17 )  ;
assign n5752 = in[31:24] ;
assign n5753 =  ( n5752 ) == ( bv_8_251_n21 )  ;
assign n5754 = in[31:24] ;
assign n5755 =  ( n5754 ) == ( bv_8_250_n25 )  ;
assign n5756 = in[31:24] ;
assign n5757 =  ( n5756 ) == ( bv_8_249_n29 )  ;
assign n5758 = in[31:24] ;
assign n5759 =  ( n5758 ) == ( bv_8_248_n33 )  ;
assign n5760 = in[31:24] ;
assign n5761 =  ( n5760 ) == ( bv_8_247_n37 )  ;
assign n5762 = in[31:24] ;
assign n5763 =  ( n5762 ) == ( bv_8_246_n41 )  ;
assign n5764 = in[31:24] ;
assign n5765 =  ( n5764 ) == ( bv_8_245_n45 )  ;
assign n5766 = in[31:24] ;
assign n5767 =  ( n5766 ) == ( bv_8_244_n49 )  ;
assign n5768 = in[31:24] ;
assign n5769 =  ( n5768 ) == ( bv_8_243_n53 )  ;
assign n5770 = in[31:24] ;
assign n5771 =  ( n5770 ) == ( bv_8_242_n57 )  ;
assign n5772 = in[31:24] ;
assign n5773 =  ( n5772 ) == ( bv_8_241_n61 )  ;
assign n5774 = in[31:24] ;
assign n5775 =  ( n5774 ) == ( bv_8_240_n65 )  ;
assign n5776 = in[31:24] ;
assign n5777 =  ( n5776 ) == ( bv_8_239_n69 )  ;
assign n5778 = in[31:24] ;
assign n5779 =  ( n5778 ) == ( bv_8_238_n73 )  ;
assign n5780 = in[31:24] ;
assign n5781 =  ( n5780 ) == ( bv_8_237_n77 )  ;
assign n5782 = in[31:24] ;
assign n5783 =  ( n5782 ) == ( bv_8_236_n81 )  ;
assign n5784 = in[31:24] ;
assign n5785 =  ( n5784 ) == ( bv_8_235_n85 )  ;
assign n5786 = in[31:24] ;
assign n5787 =  ( n5786 ) == ( bv_8_234_n89 )  ;
assign n5788 = in[31:24] ;
assign n5789 =  ( n5788 ) == ( bv_8_233_n87 )  ;
assign n5790 = in[31:24] ;
assign n5791 =  ( n5790 ) == ( bv_8_232_n96 )  ;
assign n5792 = in[31:24] ;
assign n5793 =  ( n5792 ) == ( bv_8_231_n100 )  ;
assign n5794 = in[31:24] ;
assign n5795 =  ( n5794 ) == ( bv_8_230_n47 )  ;
assign n5796 = in[31:24] ;
assign n5797 =  ( n5796 ) == ( bv_8_229_n107 )  ;
assign n5798 = in[31:24] ;
assign n5799 =  ( n5798 ) == ( bv_8_228_n111 )  ;
assign n5800 = in[31:24] ;
assign n5801 =  ( n5800 ) == ( bv_8_227_n115 )  ;
assign n5802 = in[31:24] ;
assign n5803 =  ( n5802 ) == ( bv_8_226_n119 )  ;
assign n5804 = in[31:24] ;
assign n5805 =  ( n5804 ) == ( bv_8_225_n123 )  ;
assign n5806 = in[31:24] ;
assign n5807 =  ( n5806 ) == ( bv_8_224_n126 )  ;
assign n5808 = in[31:24] ;
assign n5809 =  ( n5808 ) == ( bv_8_223_n71 )  ;
assign n5810 = in[31:24] ;
assign n5811 =  ( n5810 ) == ( bv_8_222_n132 )  ;
assign n5812 = in[31:24] ;
assign n5813 =  ( n5812 ) == ( bv_8_221_n136 )  ;
assign n5814 = in[31:24] ;
assign n5815 =  ( n5814 ) == ( bv_8_220_n140 )  ;
assign n5816 = in[31:24] ;
assign n5817 =  ( n5816 ) == ( bv_8_219_n144 )  ;
assign n5818 = in[31:24] ;
assign n5819 =  ( n5818 ) == ( bv_8_218_n148 )  ;
assign n5820 = in[31:24] ;
assign n5821 =  ( n5820 ) == ( bv_8_217_n109 )  ;
assign n5822 = in[31:24] ;
assign n5823 =  ( n5822 ) == ( bv_8_216_n155 )  ;
assign n5824 = in[31:24] ;
assign n5825 =  ( n5824 ) == ( bv_8_215_n159 )  ;
assign n5826 = in[31:24] ;
assign n5827 =  ( n5826 ) == ( bv_8_214_n163 )  ;
assign n5828 = in[31:24] ;
assign n5829 =  ( n5828 ) == ( bv_8_213_n166 )  ;
assign n5830 = in[31:24] ;
assign n5831 =  ( n5830 ) == ( bv_8_212_n170 )  ;
assign n5832 = in[31:24] ;
assign n5833 =  ( n5832 ) == ( bv_8_211_n174 )  ;
assign n5834 = in[31:24] ;
assign n5835 =  ( n5834 ) == ( bv_8_210_n178 )  ;
assign n5836 = in[31:24] ;
assign n5837 =  ( n5836 ) == ( bv_8_209_n182 )  ;
assign n5838 = in[31:24] ;
assign n5839 =  ( n5838 ) == ( bv_8_208_n186 )  ;
assign n5840 = in[31:24] ;
assign n5841 =  ( n5840 ) == ( bv_8_207_n190 )  ;
assign n5842 = in[31:24] ;
assign n5843 =  ( n5842 ) == ( bv_8_206_n83 )  ;
assign n5844 = in[31:24] ;
assign n5845 =  ( n5844 ) == ( bv_8_205_n197 )  ;
assign n5846 = in[31:24] ;
assign n5847 =  ( n5846 ) == ( bv_8_204_n201 )  ;
assign n5848 = in[31:24] ;
assign n5849 =  ( n5848 ) == ( bv_8_203_n205 )  ;
assign n5850 = in[31:24] ;
assign n5851 =  ( n5850 ) == ( bv_8_202_n209 )  ;
assign n5852 = in[31:24] ;
assign n5853 =  ( n5852 ) == ( bv_8_201_n213 )  ;
assign n5854 = in[31:24] ;
assign n5855 =  ( n5854 ) == ( bv_8_200_n216 )  ;
assign n5856 = in[31:24] ;
assign n5857 =  ( n5856 ) == ( bv_8_199_n219 )  ;
assign n5858 = in[31:24] ;
assign n5859 =  ( n5858 ) == ( bv_8_198_n221 )  ;
assign n5860 = in[31:24] ;
assign n5861 =  ( n5860 ) == ( bv_8_197_n226 )  ;
assign n5862 = in[31:24] ;
assign n5863 =  ( n5862 ) == ( bv_8_196_n230 )  ;
assign n5864 = in[31:24] ;
assign n5865 =  ( n5864 ) == ( bv_8_195_n234 )  ;
assign n5866 = in[31:24] ;
assign n5867 =  ( n5866 ) == ( bv_8_194_n238 )  ;
assign n5868 = in[31:24] ;
assign n5869 =  ( n5868 ) == ( bv_8_193_n138 )  ;
assign n5870 = in[31:24] ;
assign n5871 =  ( n5870 ) == ( bv_8_192_n245 )  ;
assign n5872 = in[31:24] ;
assign n5873 =  ( n5872 ) == ( bv_8_191_n51 )  ;
assign n5874 = in[31:24] ;
assign n5875 =  ( n5874 ) == ( bv_8_190_n252 )  ;
assign n5876 = in[31:24] ;
assign n5877 =  ( n5876 ) == ( bv_8_189_n199 )  ;
assign n5878 = in[31:24] ;
assign n5879 =  ( n5878 ) == ( bv_8_188_n259 )  ;
assign n5880 = in[31:24] ;
assign n5881 =  ( n5880 ) == ( bv_8_187_n11 )  ;
assign n5882 = in[31:24] ;
assign n5883 =  ( n5882 ) == ( bv_8_186_n247 )  ;
assign n5884 = in[31:24] ;
assign n5885 =  ( n5884 ) == ( bv_8_185_n146 )  ;
assign n5886 = in[31:24] ;
assign n5887 =  ( n5886 ) == ( bv_8_184_n270 )  ;
assign n5888 = in[31:24] ;
assign n5889 =  ( n5888 ) == ( bv_8_183_n274 )  ;
assign n5890 = in[31:24] ;
assign n5891 =  ( n5890 ) == ( bv_8_182_n278 )  ;
assign n5892 = in[31:24] ;
assign n5893 =  ( n5892 ) == ( bv_8_181_n180 )  ;
assign n5894 = in[31:24] ;
assign n5895 =  ( n5894 ) == ( bv_8_180_n224 )  ;
assign n5896 = in[31:24] ;
assign n5897 =  ( n5896 ) == ( bv_8_179_n287 )  ;
assign n5898 = in[31:24] ;
assign n5899 =  ( n5898 ) == ( bv_8_178_n291 )  ;
assign n5900 = in[31:24] ;
assign n5901 =  ( n5900 ) == ( bv_8_177_n295 )  ;
assign n5902 = in[31:24] ;
assign n5903 =  ( n5902 ) == ( bv_8_176_n19 )  ;
assign n5904 = in[31:24] ;
assign n5905 =  ( n5904 ) == ( bv_8_175_n300 )  ;
assign n5906 = in[31:24] ;
assign n5907 =  ( n5906 ) == ( bv_8_174_n254 )  ;
assign n5908 = in[31:24] ;
assign n5909 =  ( n5908 ) == ( bv_8_173_n306 )  ;
assign n5910 = in[31:24] ;
assign n5911 =  ( n5910 ) == ( bv_8_172_n310 )  ;
assign n5912 = in[31:24] ;
assign n5913 =  ( n5912 ) == ( bv_8_171_n314 )  ;
assign n5914 = in[31:24] ;
assign n5915 =  ( n5914 ) == ( bv_8_170_n318 )  ;
assign n5916 = in[31:24] ;
assign n5917 =  ( n5916 ) == ( bv_8_169_n276 )  ;
assign n5918 = in[31:24] ;
assign n5919 =  ( n5918 ) == ( bv_8_168_n323 )  ;
assign n5920 = in[31:24] ;
assign n5921 =  ( n5920 ) == ( bv_8_167_n326 )  ;
assign n5922 = in[31:24] ;
assign n5923 =  ( n5922 ) == ( bv_8_166_n228 )  ;
assign n5924 = in[31:24] ;
assign n5925 =  ( n5924 ) == ( bv_8_165_n333 )  ;
assign n5926 = in[31:24] ;
assign n5927 =  ( n5926 ) == ( bv_8_164_n337 )  ;
assign n5928 = in[31:24] ;
assign n5929 =  ( n5928 ) == ( bv_8_163_n341 )  ;
assign n5930 = in[31:24] ;
assign n5931 =  ( n5930 ) == ( bv_8_162_n345 )  ;
assign n5932 = in[31:24] ;
assign n5933 =  ( n5932 ) == ( bv_8_161_n63 )  ;
assign n5934 = in[31:24] ;
assign n5935 =  ( n5934 ) == ( bv_8_160_n352 )  ;
assign n5936 = in[31:24] ;
assign n5937 =  ( n5936 ) == ( bv_8_159_n355 )  ;
assign n5938 = in[31:24] ;
assign n5939 =  ( n5938 ) == ( bv_8_158_n130 )  ;
assign n5940 = in[31:24] ;
assign n5941 =  ( n5940 ) == ( bv_8_157_n361 )  ;
assign n5942 = in[31:24] ;
assign n5943 =  ( n5942 ) == ( bv_8_156_n365 )  ;
assign n5944 = in[31:24] ;
assign n5945 =  ( n5944 ) == ( bv_8_155_n98 )  ;
assign n5946 = in[31:24] ;
assign n5947 =  ( n5946 ) == ( bv_8_154_n371 )  ;
assign n5948 = in[31:24] ;
assign n5949 =  ( n5948 ) == ( bv_8_153_n31 )  ;
assign n5950 = in[31:24] ;
assign n5951 =  ( n5950 ) == ( bv_8_152_n121 )  ;
assign n5952 = in[31:24] ;
assign n5953 =  ( n5952 ) == ( bv_8_151_n379 )  ;
assign n5954 = in[31:24] ;
assign n5955 =  ( n5954 ) == ( bv_8_150_n383 )  ;
assign n5956 = in[31:24] ;
assign n5957 =  ( n5956 ) == ( bv_8_149_n308 )  ;
assign n5958 = in[31:24] ;
assign n5959 =  ( n5958 ) == ( bv_8_148_n102 )  ;
assign n5960 = in[31:24] ;
assign n5961 =  ( n5960 ) == ( bv_8_147_n393 )  ;
assign n5962 = in[31:24] ;
assign n5963 =  ( n5962 ) == ( bv_8_146_n396 )  ;
assign n5964 = in[31:24] ;
assign n5965 =  ( n5964 ) == ( bv_8_145_n312 )  ;
assign n5966 = in[31:24] ;
assign n5967 =  ( n5966 ) == ( bv_8_144_n385 )  ;
assign n5968 = in[31:24] ;
assign n5969 =  ( n5968 ) == ( bv_8_143_n406 )  ;
assign n5970 = in[31:24] ;
assign n5971 =  ( n5970 ) == ( bv_8_142_n105 )  ;
assign n5972 = in[31:24] ;
assign n5973 =  ( n5972 ) == ( bv_8_141_n285 )  ;
assign n5974 = in[31:24] ;
assign n5975 =  ( n5974 ) == ( bv_8_140_n67 )  ;
assign n5976 = in[31:24] ;
assign n5977 =  ( n5976 ) == ( bv_8_139_n195 )  ;
assign n5978 = in[31:24] ;
assign n5979 =  ( n5978 ) == ( bv_8_138_n192 )  ;
assign n5980 = in[31:24] ;
assign n5981 =  ( n5980 ) == ( bv_8_137_n59 )  ;
assign n5982 = in[31:24] ;
assign n5983 =  ( n5982 ) == ( bv_8_136_n381 )  ;
assign n5984 = in[31:24] ;
assign n5985 =  ( n5984 ) == ( bv_8_135_n91 )  ;
assign n5986 = in[31:24] ;
assign n5987 =  ( n5986 ) == ( bv_8_134_n142 )  ;
assign n5988 = in[31:24] ;
assign n5989 =  ( n5988 ) == ( bv_8_133_n435 )  ;
assign n5990 = in[31:24] ;
assign n5991 =  ( n5990 ) == ( bv_8_132_n438 )  ;
assign n5992 = in[31:24] ;
assign n5993 =  ( n5992 ) == ( bv_8_131_n442 )  ;
assign n5994 = in[31:24] ;
assign n5995 =  ( n5994 ) == ( bv_8_130_n445 )  ;
assign n5996 = in[31:24] ;
assign n5997 =  ( n5996 ) == ( bv_8_129_n401 )  ;
assign n5998 = in[31:24] ;
assign n5999 =  ( n5998 ) == ( bv_8_128_n452 )  ;
assign n6000 = in[31:24] ;
assign n6001 =  ( n6000 ) == ( bv_8_127_n455 )  ;
assign n6002 = in[31:24] ;
assign n6003 =  ( n6002 ) == ( bv_8_126_n423 )  ;
assign n6004 = in[31:24] ;
assign n6005 =  ( n6004 ) == ( bv_8_125_n460 )  ;
assign n6006 = in[31:24] ;
assign n6007 =  ( n6006 ) == ( bv_8_124_n463 )  ;
assign n6008 = in[31:24] ;
assign n6009 =  ( n6008 ) == ( bv_8_123_n467 )  ;
assign n6010 = in[31:24] ;
assign n6011 =  ( n6010 ) == ( bv_8_122_n257 )  ;
assign n6012 = in[31:24] ;
assign n6013 =  ( n6012 ) == ( bv_8_121_n302 )  ;
assign n6014 = in[31:24] ;
assign n6015 =  ( n6014 ) == ( bv_8_120_n243 )  ;
assign n6016 = in[31:24] ;
assign n6017 =  ( n6016 ) == ( bv_8_119_n477 )  ;
assign n6018 = in[31:24] ;
assign n6019 =  ( n6018 ) == ( bv_8_118_n480 )  ;
assign n6020 = in[31:24] ;
assign n6021 =  ( n6020 ) == ( bv_8_117_n484 )  ;
assign n6022 = in[31:24] ;
assign n6023 =  ( n6022 ) == ( bv_8_116_n211 )  ;
assign n6024 = in[31:24] ;
assign n6025 =  ( n6024 ) == ( bv_8_115_n408 )  ;
assign n6026 = in[31:24] ;
assign n6027 =  ( n6026 ) == ( bv_8_114_n491 )  ;
assign n6028 = in[31:24] ;
assign n6029 =  ( n6028 ) == ( bv_8_113_n495 )  ;
assign n6030 = in[31:24] ;
assign n6031 =  ( n6030 ) == ( bv_8_112_n188 )  ;
assign n6032 = in[31:24] ;
assign n6033 =  ( n6032 ) == ( bv_8_111_n501 )  ;
assign n6034 = in[31:24] ;
assign n6035 =  ( n6034 ) == ( bv_8_110_n504 )  ;
assign n6036 = in[31:24] ;
assign n6037 =  ( n6036 ) == ( bv_8_109_n289 )  ;
assign n6038 = in[31:24] ;
assign n6039 =  ( n6038 ) == ( bv_8_108_n272 )  ;
assign n6040 = in[31:24] ;
assign n6041 =  ( n6040 ) == ( bv_8_107_n513 )  ;
assign n6042 = in[31:24] ;
assign n6043 =  ( n6042 ) == ( bv_8_106_n516 )  ;
assign n6044 = in[31:24] ;
assign n6045 =  ( n6044 ) == ( bv_8_105_n113 )  ;
assign n6046 = in[31:24] ;
assign n6047 =  ( n6046 ) == ( bv_8_104_n39 )  ;
assign n6048 = in[31:24] ;
assign n6049 =  ( n6048 ) == ( bv_8_103_n525 )  ;
assign n6050 = in[31:24] ;
assign n6051 =  ( n6050 ) == ( bv_8_102_n176 )  ;
assign n6052 = in[31:24] ;
assign n6053 =  ( n6052 ) == ( bv_8_101_n261 )  ;
assign n6054 = in[31:24] ;
assign n6055 =  ( n6054 ) == ( bv_8_100_n417 )  ;
assign n6056 = in[31:24] ;
assign n6057 =  ( n6056 ) == ( bv_8_99_n537 )  ;
assign n6058 = in[31:24] ;
assign n6059 =  ( n6058 ) == ( bv_8_98_n316 )  ;
assign n6060 = in[31:24] ;
assign n6061 =  ( n6060 ) == ( bv_8_97_n157 )  ;
assign n6062 = in[31:24] ;
assign n6063 =  ( n6062 ) == ( bv_8_96_n404 )  ;
assign n6064 = in[31:24] ;
assign n6065 =  ( n6064 ) == ( bv_8_95_n440 )  ;
assign n6066 = in[31:24] ;
assign n6067 =  ( n6066 ) == ( bv_8_94_n363 )  ;
assign n6068 = in[31:24] ;
assign n6069 =  ( n6068 ) == ( bv_8_93_n414 )  ;
assign n6070 = in[31:24] ;
assign n6071 =  ( n6070 ) == ( bv_8_92_n328 )  ;
assign n6072 = in[31:24] ;
assign n6073 =  ( n6072 ) == ( bv_8_91_n557 )  ;
assign n6074 = in[31:24] ;
assign n6075 =  ( n6074 ) == ( bv_8_90_n561 )  ;
assign n6076 = in[31:24] ;
assign n6077 =  ( n6076 ) == ( bv_8_89_n564 )  ;
assign n6078 = in[31:24] ;
assign n6079 =  ( n6078 ) == ( bv_8_88_n549 )  ;
assign n6080 = in[31:24] ;
assign n6081 =  ( n6080 ) == ( bv_8_87_n150 )  ;
assign n6082 = in[31:24] ;
assign n6083 =  ( n6082 ) == ( bv_8_86_n268 )  ;
assign n6084 = in[31:24] ;
assign n6085 =  ( n6084 ) == ( bv_8_85_n79 )  ;
assign n6086 = in[31:24] ;
assign n6087 =  ( n6086 ) == ( bv_8_84_n15 )  ;
assign n6088 = in[31:24] ;
assign n6089 =  ( n6088 ) == ( bv_8_83_n578 )  ;
assign n6090 = in[31:24] ;
assign n6091 =  ( n6090 ) == ( bv_8_82_n581 )  ;
assign n6092 = in[31:24] ;
assign n6093 =  ( n6092 ) == ( bv_8_81_n499 )  ;
assign n6094 = in[31:24] ;
assign n6095 =  ( n6094 ) == ( bv_8_80_n511 )  ;
assign n6096 = in[31:24] ;
assign n6097 =  ( n6096 ) == ( bv_8_79_n398 )  ;
assign n6098 = in[31:24] ;
assign n6099 =  ( n6098 ) == ( bv_8_78_n280 )  ;
assign n6100 = in[31:24] ;
assign n6101 =  ( n6100 ) == ( bv_8_77_n532 )  ;
assign n6102 = in[31:24] ;
assign n6103 =  ( n6102 ) == ( bv_8_76_n552 )  ;
assign n6104 = in[31:24] ;
assign n6105 =  ( n6104 ) == ( bv_8_75_n203 )  ;
assign n6106 = in[31:24] ;
assign n6107 =  ( n6106 ) == ( bv_8_74_n555 )  ;
assign n6108 = in[31:24] ;
assign n6109 =  ( n6108 ) == ( bv_8_73_n339 )  ;
assign n6110 = in[31:24] ;
assign n6111 =  ( n6110 ) == ( bv_8_72_n172 )  ;
assign n6112 = in[31:24] ;
assign n6113 =  ( n6112 ) == ( bv_8_71_n608 )  ;
assign n6114 = in[31:24] ;
assign n6115 =  ( n6114 ) == ( bv_8_70_n377 )  ;
assign n6116 = in[31:24] ;
assign n6117 =  ( n6116 ) == ( bv_8_69_n523 )  ;
assign n6118 = in[31:24] ;
assign n6119 =  ( n6118 ) == ( bv_8_68_n433 )  ;
assign n6120 = in[31:24] ;
assign n6121 =  ( n6120 ) == ( bv_8_67_n535 )  ;
assign n6122 = in[31:24] ;
assign n6123 =  ( n6122 ) == ( bv_8_66_n43 )  ;
assign n6124 = in[31:24] ;
assign n6125 =  ( n6124 ) == ( bv_8_65_n35 )  ;
assign n6126 = in[31:24] ;
assign n6127 =  ( n6126 ) == ( bv_8_64_n493 )  ;
assign n6128 = in[31:24] ;
assign n6129 =  ( n6128 ) == ( bv_8_63_n629 )  ;
assign n6130 = in[31:24] ;
assign n6131 =  ( n6130 ) == ( bv_8_62_n184 )  ;
assign n6132 = in[31:24] ;
assign n6133 =  ( n6132 ) == ( bv_8_61_n420 )  ;
assign n6134 = in[31:24] ;
assign n6135 =  ( n6134 ) == ( bv_8_60_n508 )  ;
assign n6136 = in[31:24] ;
assign n6137 =  ( n6136 ) == ( bv_8_59_n604 )  ;
assign n6138 = in[31:24] ;
assign n6139 =  ( n6138 ) == ( bv_8_58_n347 )  ;
assign n6140 = in[31:24] ;
assign n6141 =  ( n6140 ) == ( bv_8_57_n559 )  ;
assign n6142 = in[31:24] ;
assign n6143 =  ( n6142 ) == ( bv_8_56_n482 )  ;
assign n6144 = in[31:24] ;
assign n6145 =  ( n6144 ) == ( bv_8_55_n293 )  ;
assign n6146 = in[31:24] ;
assign n6147 =  ( n6146 ) == ( bv_8_54_n651 )  ;
assign n6148 = in[31:24] ;
assign n6149 =  ( n6148 ) == ( bv_8_53_n153 )  ;
assign n6150 = in[31:24] ;
assign n6151 =  ( n6150 ) == ( bv_8_52_n657 )  ;
assign n6152 = in[31:24] ;
assign n6153 =  ( n6152 ) == ( bv_8_51_n529 )  ;
assign n6154 = in[31:24] ;
assign n6155 =  ( n6154 ) == ( bv_8_50_n350 )  ;
assign n6156 = in[31:24] ;
assign n6157 =  ( n6156 ) == ( bv_8_49_n666 )  ;
assign n6158 = in[31:24] ;
assign n6159 =  ( n6158 ) == ( bv_8_48_n669 )  ;
assign n6160 = in[31:24] ;
assign n6161 =  ( n6160 ) == ( bv_8_47_n592 )  ;
assign n6162 = in[31:24] ;
assign n6163 =  ( n6162 ) == ( bv_8_46_n236 )  ;
assign n6164 = in[31:24] ;
assign n6165 =  ( n6164 ) == ( bv_8_45_n27 )  ;
assign n6166 = in[31:24] ;
assign n6167 =  ( n6166 ) == ( bv_8_44_n622 )  ;
assign n6168 = in[31:24] ;
assign n6169 =  ( n6168 ) == ( bv_8_43_n682 )  ;
assign n6170 = in[31:24] ;
assign n6171 =  ( n6170 ) == ( bv_8_42_n388 )  ;
assign n6172 = in[31:24] ;
assign n6173 =  ( n6172 ) == ( bv_8_41_n597 )  ;
assign n6174 = in[31:24] ;
assign n6175 =  ( n6174 ) == ( bv_8_40_n75 )  ;
assign n6176 = in[31:24] ;
assign n6177 =  ( n6176 ) == ( bv_8_39_n635 )  ;
assign n6178 = in[31:24] ;
assign n6179 =  ( n6178 ) == ( bv_8_38_n693 )  ;
assign n6180 = in[31:24] ;
assign n6181 =  ( n6180 ) == ( bv_8_37_n240 )  ;
assign n6182 = in[31:24] ;
assign n6183 =  ( n6182 ) == ( bv_8_36_n331 )  ;
assign n6184 = in[31:24] ;
assign n6185 =  ( n6184 ) == ( bv_8_35_n664 )  ;
assign n6186 = in[31:24] ;
assign n6187 =  ( n6186 ) == ( bv_8_34_n391 )  ;
assign n6188 = in[31:24] ;
assign n6189 =  ( n6188 ) == ( bv_8_33_n469 )  ;
assign n6190 = in[31:24] ;
assign n6191 =  ( n6190 ) == ( bv_8_32_n576 )  ;
assign n6192 = in[31:24] ;
assign n6193 =  ( n6192 ) == ( bv_8_31_n207 )  ;
assign n6194 = in[31:24] ;
assign n6195 =  ( n6194 ) == ( bv_8_30_n94 )  ;
assign n6196 = in[31:24] ;
assign n6197 =  ( n6196 ) == ( bv_8_29_n134 )  ;
assign n6198 = in[31:24] ;
assign n6199 =  ( n6198 ) == ( bv_8_28_n232 )  ;
assign n6200 = in[31:24] ;
assign n6201 =  ( n6200 ) == ( bv_8_27_n616 )  ;
assign n6202 = in[31:24] ;
assign n6203 =  ( n6202 ) == ( bv_8_26_n619 )  ;
assign n6204 = in[31:24] ;
assign n6205 =  ( n6204 ) == ( bv_8_25_n411 )  ;
assign n6206 = in[31:24] ;
assign n6207 =  ( n6206 ) == ( bv_8_24_n659 )  ;
assign n6208 = in[31:24] ;
assign n6209 =  ( n6208 ) == ( bv_8_23_n430 )  ;
assign n6210 = in[31:24] ;
assign n6211 =  ( n6210 ) == ( bv_8_22_n7 )  ;
assign n6212 = in[31:24] ;
assign n6213 =  ( n6212 ) == ( bv_8_21_n674 )  ;
assign n6214 = in[31:24] ;
assign n6215 =  ( n6214 ) == ( bv_8_20_n369 )  ;
assign n6216 = in[31:24] ;
assign n6217 =  ( n6216 ) == ( bv_8_19_n447 )  ;
assign n6218 = in[31:24] ;
assign n6219 =  ( n6218 ) == ( bv_8_18_n644 )  ;
assign n6220 = in[31:24] ;
assign n6221 =  ( n6220 ) == ( bv_8_17_n117 )  ;
assign n6222 = in[31:24] ;
assign n6223 =  ( n6222 ) == ( bv_8_16_n465 )  ;
assign n6224 = in[31:24] ;
assign n6225 =  ( n6224 ) == ( bv_8_15_n23 )  ;
assign n6226 = in[31:24] ;
assign n6227 =  ( n6226 ) == ( bv_8_14_n161 )  ;
assign n6228 = in[31:24] ;
assign n6229 =  ( n6228 ) == ( bv_8_13_n55 )  ;
assign n6230 = in[31:24] ;
assign n6231 =  ( n6230 ) == ( bv_8_12_n450 )  ;
assign n6232 = in[31:24] ;
assign n6233 =  ( n6232 ) == ( bv_8_11_n359 )  ;
assign n6234 = in[31:24] ;
assign n6235 =  ( n6234 ) == ( bv_8_10_n343 )  ;
assign n6236 = in[31:24] ;
assign n6237 =  ( n6236 ) == ( bv_8_9_n627 )  ;
assign n6238 = in[31:24] ;
assign n6239 =  ( n6238 ) == ( bv_8_8_n250 )  ;
assign n6240 = in[31:24] ;
assign n6241 =  ( n6240 ) == ( bv_8_7_n647 )  ;
assign n6242 = in[31:24] ;
assign n6243 =  ( n6242 ) == ( bv_8_6_n335 )  ;
assign n6244 = in[31:24] ;
assign n6245 =  ( n6244 ) == ( bv_8_5_n653 )  ;
assign n6246 = in[31:24] ;
assign n6247 =  ( n6246 ) == ( bv_8_4_n671 )  ;
assign n6248 = in[31:24] ;
assign n6249 =  ( n6248 ) == ( bv_8_3_n168 )  ;
assign n6250 = in[31:24] ;
assign n6251 =  ( n6250 ) == ( bv_8_2_n518 )  ;
assign n6252 = in[31:24] ;
assign n6253 =  ( n6252 ) == ( bv_8_1_n753 )  ;
assign n6254 = in[31:24] ;
assign n6255 =  ( n6254 ) == ( bv_8_0_n583 )  ;
assign n6256 =  ( n6255 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n6257 =  ( n6253 ) ? ( bv_8_124_n463 ) : ( n6256 ) ;
assign n6258 =  ( n6251 ) ? ( bv_8_119_n477 ) : ( n6257 ) ;
assign n6259 =  ( n6249 ) ? ( bv_8_123_n467 ) : ( n6258 ) ;
assign n6260 =  ( n6247 ) ? ( bv_8_242_n57 ) : ( n6259 ) ;
assign n6261 =  ( n6245 ) ? ( bv_8_107_n513 ) : ( n6260 ) ;
assign n6262 =  ( n6243 ) ? ( bv_8_111_n501 ) : ( n6261 ) ;
assign n6263 =  ( n6241 ) ? ( bv_8_197_n226 ) : ( n6262 ) ;
assign n6264 =  ( n6239 ) ? ( bv_8_48_n669 ) : ( n6263 ) ;
assign n6265 =  ( n6237 ) ? ( bv_8_1_n753 ) : ( n6264 ) ;
assign n6266 =  ( n6235 ) ? ( bv_8_103_n525 ) : ( n6265 ) ;
assign n6267 =  ( n6233 ) ? ( bv_8_43_n682 ) : ( n6266 ) ;
assign n6268 =  ( n6231 ) ? ( bv_8_254_n9 ) : ( n6267 ) ;
assign n6269 =  ( n6229 ) ? ( bv_8_215_n159 ) : ( n6268 ) ;
assign n6270 =  ( n6227 ) ? ( bv_8_171_n314 ) : ( n6269 ) ;
assign n6271 =  ( n6225 ) ? ( bv_8_118_n480 ) : ( n6270 ) ;
assign n6272 =  ( n6223 ) ? ( bv_8_202_n209 ) : ( n6271 ) ;
assign n6273 =  ( n6221 ) ? ( bv_8_130_n445 ) : ( n6272 ) ;
assign n6274 =  ( n6219 ) ? ( bv_8_201_n213 ) : ( n6273 ) ;
assign n6275 =  ( n6217 ) ? ( bv_8_125_n460 ) : ( n6274 ) ;
assign n6276 =  ( n6215 ) ? ( bv_8_250_n25 ) : ( n6275 ) ;
assign n6277 =  ( n6213 ) ? ( bv_8_89_n564 ) : ( n6276 ) ;
assign n6278 =  ( n6211 ) ? ( bv_8_71_n608 ) : ( n6277 ) ;
assign n6279 =  ( n6209 ) ? ( bv_8_240_n65 ) : ( n6278 ) ;
assign n6280 =  ( n6207 ) ? ( bv_8_173_n306 ) : ( n6279 ) ;
assign n6281 =  ( n6205 ) ? ( bv_8_212_n170 ) : ( n6280 ) ;
assign n6282 =  ( n6203 ) ? ( bv_8_162_n345 ) : ( n6281 ) ;
assign n6283 =  ( n6201 ) ? ( bv_8_175_n300 ) : ( n6282 ) ;
assign n6284 =  ( n6199 ) ? ( bv_8_156_n365 ) : ( n6283 ) ;
assign n6285 =  ( n6197 ) ? ( bv_8_164_n337 ) : ( n6284 ) ;
assign n6286 =  ( n6195 ) ? ( bv_8_114_n491 ) : ( n6285 ) ;
assign n6287 =  ( n6193 ) ? ( bv_8_192_n245 ) : ( n6286 ) ;
assign n6288 =  ( n6191 ) ? ( bv_8_183_n274 ) : ( n6287 ) ;
assign n6289 =  ( n6189 ) ? ( bv_8_253_n13 ) : ( n6288 ) ;
assign n6290 =  ( n6187 ) ? ( bv_8_147_n393 ) : ( n6289 ) ;
assign n6291 =  ( n6185 ) ? ( bv_8_38_n693 ) : ( n6290 ) ;
assign n6292 =  ( n6183 ) ? ( bv_8_54_n651 ) : ( n6291 ) ;
assign n6293 =  ( n6181 ) ? ( bv_8_63_n629 ) : ( n6292 ) ;
assign n6294 =  ( n6179 ) ? ( bv_8_247_n37 ) : ( n6293 ) ;
assign n6295 =  ( n6177 ) ? ( bv_8_204_n201 ) : ( n6294 ) ;
assign n6296 =  ( n6175 ) ? ( bv_8_52_n657 ) : ( n6295 ) ;
assign n6297 =  ( n6173 ) ? ( bv_8_165_n333 ) : ( n6296 ) ;
assign n6298 =  ( n6171 ) ? ( bv_8_229_n107 ) : ( n6297 ) ;
assign n6299 =  ( n6169 ) ? ( bv_8_241_n61 ) : ( n6298 ) ;
assign n6300 =  ( n6167 ) ? ( bv_8_113_n495 ) : ( n6299 ) ;
assign n6301 =  ( n6165 ) ? ( bv_8_216_n155 ) : ( n6300 ) ;
assign n6302 =  ( n6163 ) ? ( bv_8_49_n666 ) : ( n6301 ) ;
assign n6303 =  ( n6161 ) ? ( bv_8_21_n674 ) : ( n6302 ) ;
assign n6304 =  ( n6159 ) ? ( bv_8_4_n671 ) : ( n6303 ) ;
assign n6305 =  ( n6157 ) ? ( bv_8_199_n219 ) : ( n6304 ) ;
assign n6306 =  ( n6155 ) ? ( bv_8_35_n664 ) : ( n6305 ) ;
assign n6307 =  ( n6153 ) ? ( bv_8_195_n234 ) : ( n6306 ) ;
assign n6308 =  ( n6151 ) ? ( bv_8_24_n659 ) : ( n6307 ) ;
assign n6309 =  ( n6149 ) ? ( bv_8_150_n383 ) : ( n6308 ) ;
assign n6310 =  ( n6147 ) ? ( bv_8_5_n653 ) : ( n6309 ) ;
assign n6311 =  ( n6145 ) ? ( bv_8_154_n371 ) : ( n6310 ) ;
assign n6312 =  ( n6143 ) ? ( bv_8_7_n647 ) : ( n6311 ) ;
assign n6313 =  ( n6141 ) ? ( bv_8_18_n644 ) : ( n6312 ) ;
assign n6314 =  ( n6139 ) ? ( bv_8_128_n452 ) : ( n6313 ) ;
assign n6315 =  ( n6137 ) ? ( bv_8_226_n119 ) : ( n6314 ) ;
assign n6316 =  ( n6135 ) ? ( bv_8_235_n85 ) : ( n6315 ) ;
assign n6317 =  ( n6133 ) ? ( bv_8_39_n635 ) : ( n6316 ) ;
assign n6318 =  ( n6131 ) ? ( bv_8_178_n291 ) : ( n6317 ) ;
assign n6319 =  ( n6129 ) ? ( bv_8_117_n484 ) : ( n6318 ) ;
assign n6320 =  ( n6127 ) ? ( bv_8_9_n627 ) : ( n6319 ) ;
assign n6321 =  ( n6125 ) ? ( bv_8_131_n442 ) : ( n6320 ) ;
assign n6322 =  ( n6123 ) ? ( bv_8_44_n622 ) : ( n6321 ) ;
assign n6323 =  ( n6121 ) ? ( bv_8_26_n619 ) : ( n6322 ) ;
assign n6324 =  ( n6119 ) ? ( bv_8_27_n616 ) : ( n6323 ) ;
assign n6325 =  ( n6117 ) ? ( bv_8_110_n504 ) : ( n6324 ) ;
assign n6326 =  ( n6115 ) ? ( bv_8_90_n561 ) : ( n6325 ) ;
assign n6327 =  ( n6113 ) ? ( bv_8_160_n352 ) : ( n6326 ) ;
assign n6328 =  ( n6111 ) ? ( bv_8_82_n581 ) : ( n6327 ) ;
assign n6329 =  ( n6109 ) ? ( bv_8_59_n604 ) : ( n6328 ) ;
assign n6330 =  ( n6107 ) ? ( bv_8_214_n163 ) : ( n6329 ) ;
assign n6331 =  ( n6105 ) ? ( bv_8_179_n287 ) : ( n6330 ) ;
assign n6332 =  ( n6103 ) ? ( bv_8_41_n597 ) : ( n6331 ) ;
assign n6333 =  ( n6101 ) ? ( bv_8_227_n115 ) : ( n6332 ) ;
assign n6334 =  ( n6099 ) ? ( bv_8_47_n592 ) : ( n6333 ) ;
assign n6335 =  ( n6097 ) ? ( bv_8_132_n438 ) : ( n6334 ) ;
assign n6336 =  ( n6095 ) ? ( bv_8_83_n578 ) : ( n6335 ) ;
assign n6337 =  ( n6093 ) ? ( bv_8_209_n182 ) : ( n6336 ) ;
assign n6338 =  ( n6091 ) ? ( bv_8_0_n583 ) : ( n6337 ) ;
assign n6339 =  ( n6089 ) ? ( bv_8_237_n77 ) : ( n6338 ) ;
assign n6340 =  ( n6087 ) ? ( bv_8_32_n576 ) : ( n6339 ) ;
assign n6341 =  ( n6085 ) ? ( bv_8_252_n17 ) : ( n6340 ) ;
assign n6342 =  ( n6083 ) ? ( bv_8_177_n295 ) : ( n6341 ) ;
assign n6343 =  ( n6081 ) ? ( bv_8_91_n557 ) : ( n6342 ) ;
assign n6344 =  ( n6079 ) ? ( bv_8_106_n516 ) : ( n6343 ) ;
assign n6345 =  ( n6077 ) ? ( bv_8_203_n205 ) : ( n6344 ) ;
assign n6346 =  ( n6075 ) ? ( bv_8_190_n252 ) : ( n6345 ) ;
assign n6347 =  ( n6073 ) ? ( bv_8_57_n559 ) : ( n6346 ) ;
assign n6348 =  ( n6071 ) ? ( bv_8_74_n555 ) : ( n6347 ) ;
assign n6349 =  ( n6069 ) ? ( bv_8_76_n552 ) : ( n6348 ) ;
assign n6350 =  ( n6067 ) ? ( bv_8_88_n549 ) : ( n6349 ) ;
assign n6351 =  ( n6065 ) ? ( bv_8_207_n190 ) : ( n6350 ) ;
assign n6352 =  ( n6063 ) ? ( bv_8_208_n186 ) : ( n6351 ) ;
assign n6353 =  ( n6061 ) ? ( bv_8_239_n69 ) : ( n6352 ) ;
assign n6354 =  ( n6059 ) ? ( bv_8_170_n318 ) : ( n6353 ) ;
assign n6355 =  ( n6057 ) ? ( bv_8_251_n21 ) : ( n6354 ) ;
assign n6356 =  ( n6055 ) ? ( bv_8_67_n535 ) : ( n6355 ) ;
assign n6357 =  ( n6053 ) ? ( bv_8_77_n532 ) : ( n6356 ) ;
assign n6358 =  ( n6051 ) ? ( bv_8_51_n529 ) : ( n6357 ) ;
assign n6359 =  ( n6049 ) ? ( bv_8_133_n435 ) : ( n6358 ) ;
assign n6360 =  ( n6047 ) ? ( bv_8_69_n523 ) : ( n6359 ) ;
assign n6361 =  ( n6045 ) ? ( bv_8_249_n29 ) : ( n6360 ) ;
assign n6362 =  ( n6043 ) ? ( bv_8_2_n518 ) : ( n6361 ) ;
assign n6363 =  ( n6041 ) ? ( bv_8_127_n455 ) : ( n6362 ) ;
assign n6364 =  ( n6039 ) ? ( bv_8_80_n511 ) : ( n6363 ) ;
assign n6365 =  ( n6037 ) ? ( bv_8_60_n508 ) : ( n6364 ) ;
assign n6366 =  ( n6035 ) ? ( bv_8_159_n355 ) : ( n6365 ) ;
assign n6367 =  ( n6033 ) ? ( bv_8_168_n323 ) : ( n6366 ) ;
assign n6368 =  ( n6031 ) ? ( bv_8_81_n499 ) : ( n6367 ) ;
assign n6369 =  ( n6029 ) ? ( bv_8_163_n341 ) : ( n6368 ) ;
assign n6370 =  ( n6027 ) ? ( bv_8_64_n493 ) : ( n6369 ) ;
assign n6371 =  ( n6025 ) ? ( bv_8_143_n406 ) : ( n6370 ) ;
assign n6372 =  ( n6023 ) ? ( bv_8_146_n396 ) : ( n6371 ) ;
assign n6373 =  ( n6021 ) ? ( bv_8_157_n361 ) : ( n6372 ) ;
assign n6374 =  ( n6019 ) ? ( bv_8_56_n482 ) : ( n6373 ) ;
assign n6375 =  ( n6017 ) ? ( bv_8_245_n45 ) : ( n6374 ) ;
assign n6376 =  ( n6015 ) ? ( bv_8_188_n259 ) : ( n6375 ) ;
assign n6377 =  ( n6013 ) ? ( bv_8_182_n278 ) : ( n6376 ) ;
assign n6378 =  ( n6011 ) ? ( bv_8_218_n148 ) : ( n6377 ) ;
assign n6379 =  ( n6009 ) ? ( bv_8_33_n469 ) : ( n6378 ) ;
assign n6380 =  ( n6007 ) ? ( bv_8_16_n465 ) : ( n6379 ) ;
assign n6381 =  ( n6005 ) ? ( bv_8_255_n5 ) : ( n6380 ) ;
assign n6382 =  ( n6003 ) ? ( bv_8_243_n53 ) : ( n6381 ) ;
assign n6383 =  ( n6001 ) ? ( bv_8_210_n178 ) : ( n6382 ) ;
assign n6384 =  ( n5999 ) ? ( bv_8_205_n197 ) : ( n6383 ) ;
assign n6385 =  ( n5997 ) ? ( bv_8_12_n450 ) : ( n6384 ) ;
assign n6386 =  ( n5995 ) ? ( bv_8_19_n447 ) : ( n6385 ) ;
assign n6387 =  ( n5993 ) ? ( bv_8_236_n81 ) : ( n6386 ) ;
assign n6388 =  ( n5991 ) ? ( bv_8_95_n440 ) : ( n6387 ) ;
assign n6389 =  ( n5989 ) ? ( bv_8_151_n379 ) : ( n6388 ) ;
assign n6390 =  ( n5987 ) ? ( bv_8_68_n433 ) : ( n6389 ) ;
assign n6391 =  ( n5985 ) ? ( bv_8_23_n430 ) : ( n6390 ) ;
assign n6392 =  ( n5983 ) ? ( bv_8_196_n230 ) : ( n6391 ) ;
assign n6393 =  ( n5981 ) ? ( bv_8_167_n326 ) : ( n6392 ) ;
assign n6394 =  ( n5979 ) ? ( bv_8_126_n423 ) : ( n6393 ) ;
assign n6395 =  ( n5977 ) ? ( bv_8_61_n420 ) : ( n6394 ) ;
assign n6396 =  ( n5975 ) ? ( bv_8_100_n417 ) : ( n6395 ) ;
assign n6397 =  ( n5973 ) ? ( bv_8_93_n414 ) : ( n6396 ) ;
assign n6398 =  ( n5971 ) ? ( bv_8_25_n411 ) : ( n6397 ) ;
assign n6399 =  ( n5969 ) ? ( bv_8_115_n408 ) : ( n6398 ) ;
assign n6400 =  ( n5967 ) ? ( bv_8_96_n404 ) : ( n6399 ) ;
assign n6401 =  ( n5965 ) ? ( bv_8_129_n401 ) : ( n6400 ) ;
assign n6402 =  ( n5963 ) ? ( bv_8_79_n398 ) : ( n6401 ) ;
assign n6403 =  ( n5961 ) ? ( bv_8_220_n140 ) : ( n6402 ) ;
assign n6404 =  ( n5959 ) ? ( bv_8_34_n391 ) : ( n6403 ) ;
assign n6405 =  ( n5957 ) ? ( bv_8_42_n388 ) : ( n6404 ) ;
assign n6406 =  ( n5955 ) ? ( bv_8_144_n385 ) : ( n6405 ) ;
assign n6407 =  ( n5953 ) ? ( bv_8_136_n381 ) : ( n6406 ) ;
assign n6408 =  ( n5951 ) ? ( bv_8_70_n377 ) : ( n6407 ) ;
assign n6409 =  ( n5949 ) ? ( bv_8_238_n73 ) : ( n6408 ) ;
assign n6410 =  ( n5947 ) ? ( bv_8_184_n270 ) : ( n6409 ) ;
assign n6411 =  ( n5945 ) ? ( bv_8_20_n369 ) : ( n6410 ) ;
assign n6412 =  ( n5943 ) ? ( bv_8_222_n132 ) : ( n6411 ) ;
assign n6413 =  ( n5941 ) ? ( bv_8_94_n363 ) : ( n6412 ) ;
assign n6414 =  ( n5939 ) ? ( bv_8_11_n359 ) : ( n6413 ) ;
assign n6415 =  ( n5937 ) ? ( bv_8_219_n144 ) : ( n6414 ) ;
assign n6416 =  ( n5935 ) ? ( bv_8_224_n126 ) : ( n6415 ) ;
assign n6417 =  ( n5933 ) ? ( bv_8_50_n350 ) : ( n6416 ) ;
assign n6418 =  ( n5931 ) ? ( bv_8_58_n347 ) : ( n6417 ) ;
assign n6419 =  ( n5929 ) ? ( bv_8_10_n343 ) : ( n6418 ) ;
assign n6420 =  ( n5927 ) ? ( bv_8_73_n339 ) : ( n6419 ) ;
assign n6421 =  ( n5925 ) ? ( bv_8_6_n335 ) : ( n6420 ) ;
assign n6422 =  ( n5923 ) ? ( bv_8_36_n331 ) : ( n6421 ) ;
assign n6423 =  ( n5921 ) ? ( bv_8_92_n328 ) : ( n6422 ) ;
assign n6424 =  ( n5919 ) ? ( bv_8_194_n238 ) : ( n6423 ) ;
assign n6425 =  ( n5917 ) ? ( bv_8_211_n174 ) : ( n6424 ) ;
assign n6426 =  ( n5915 ) ? ( bv_8_172_n310 ) : ( n6425 ) ;
assign n6427 =  ( n5913 ) ? ( bv_8_98_n316 ) : ( n6426 ) ;
assign n6428 =  ( n5911 ) ? ( bv_8_145_n312 ) : ( n6427 ) ;
assign n6429 =  ( n5909 ) ? ( bv_8_149_n308 ) : ( n6428 ) ;
assign n6430 =  ( n5907 ) ? ( bv_8_228_n111 ) : ( n6429 ) ;
assign n6431 =  ( n5905 ) ? ( bv_8_121_n302 ) : ( n6430 ) ;
assign n6432 =  ( n5903 ) ? ( bv_8_231_n100 ) : ( n6431 ) ;
assign n6433 =  ( n5901 ) ? ( bv_8_200_n216 ) : ( n6432 ) ;
assign n6434 =  ( n5899 ) ? ( bv_8_55_n293 ) : ( n6433 ) ;
assign n6435 =  ( n5897 ) ? ( bv_8_109_n289 ) : ( n6434 ) ;
assign n6436 =  ( n5895 ) ? ( bv_8_141_n285 ) : ( n6435 ) ;
assign n6437 =  ( n5893 ) ? ( bv_8_213_n166 ) : ( n6436 ) ;
assign n6438 =  ( n5891 ) ? ( bv_8_78_n280 ) : ( n6437 ) ;
assign n6439 =  ( n5889 ) ? ( bv_8_169_n276 ) : ( n6438 ) ;
assign n6440 =  ( n5887 ) ? ( bv_8_108_n272 ) : ( n6439 ) ;
assign n6441 =  ( n5885 ) ? ( bv_8_86_n268 ) : ( n6440 ) ;
assign n6442 =  ( n5883 ) ? ( bv_8_244_n49 ) : ( n6441 ) ;
assign n6443 =  ( n5881 ) ? ( bv_8_234_n89 ) : ( n6442 ) ;
assign n6444 =  ( n5879 ) ? ( bv_8_101_n261 ) : ( n6443 ) ;
assign n6445 =  ( n5877 ) ? ( bv_8_122_n257 ) : ( n6444 ) ;
assign n6446 =  ( n5875 ) ? ( bv_8_174_n254 ) : ( n6445 ) ;
assign n6447 =  ( n5873 ) ? ( bv_8_8_n250 ) : ( n6446 ) ;
assign n6448 =  ( n5871 ) ? ( bv_8_186_n247 ) : ( n6447 ) ;
assign n6449 =  ( n5869 ) ? ( bv_8_120_n243 ) : ( n6448 ) ;
assign n6450 =  ( n5867 ) ? ( bv_8_37_n240 ) : ( n6449 ) ;
assign n6451 =  ( n5865 ) ? ( bv_8_46_n236 ) : ( n6450 ) ;
assign n6452 =  ( n5863 ) ? ( bv_8_28_n232 ) : ( n6451 ) ;
assign n6453 =  ( n5861 ) ? ( bv_8_166_n228 ) : ( n6452 ) ;
assign n6454 =  ( n5859 ) ? ( bv_8_180_n224 ) : ( n6453 ) ;
assign n6455 =  ( n5857 ) ? ( bv_8_198_n221 ) : ( n6454 ) ;
assign n6456 =  ( n5855 ) ? ( bv_8_232_n96 ) : ( n6455 ) ;
assign n6457 =  ( n5853 ) ? ( bv_8_221_n136 ) : ( n6456 ) ;
assign n6458 =  ( n5851 ) ? ( bv_8_116_n211 ) : ( n6457 ) ;
assign n6459 =  ( n5849 ) ? ( bv_8_31_n207 ) : ( n6458 ) ;
assign n6460 =  ( n5847 ) ? ( bv_8_75_n203 ) : ( n6459 ) ;
assign n6461 =  ( n5845 ) ? ( bv_8_189_n199 ) : ( n6460 ) ;
assign n6462 =  ( n5843 ) ? ( bv_8_139_n195 ) : ( n6461 ) ;
assign n6463 =  ( n5841 ) ? ( bv_8_138_n192 ) : ( n6462 ) ;
assign n6464 =  ( n5839 ) ? ( bv_8_112_n188 ) : ( n6463 ) ;
assign n6465 =  ( n5837 ) ? ( bv_8_62_n184 ) : ( n6464 ) ;
assign n6466 =  ( n5835 ) ? ( bv_8_181_n180 ) : ( n6465 ) ;
assign n6467 =  ( n5833 ) ? ( bv_8_102_n176 ) : ( n6466 ) ;
assign n6468 =  ( n5831 ) ? ( bv_8_72_n172 ) : ( n6467 ) ;
assign n6469 =  ( n5829 ) ? ( bv_8_3_n168 ) : ( n6468 ) ;
assign n6470 =  ( n5827 ) ? ( bv_8_246_n41 ) : ( n6469 ) ;
assign n6471 =  ( n5825 ) ? ( bv_8_14_n161 ) : ( n6470 ) ;
assign n6472 =  ( n5823 ) ? ( bv_8_97_n157 ) : ( n6471 ) ;
assign n6473 =  ( n5821 ) ? ( bv_8_53_n153 ) : ( n6472 ) ;
assign n6474 =  ( n5819 ) ? ( bv_8_87_n150 ) : ( n6473 ) ;
assign n6475 =  ( n5817 ) ? ( bv_8_185_n146 ) : ( n6474 ) ;
assign n6476 =  ( n5815 ) ? ( bv_8_134_n142 ) : ( n6475 ) ;
assign n6477 =  ( n5813 ) ? ( bv_8_193_n138 ) : ( n6476 ) ;
assign n6478 =  ( n5811 ) ? ( bv_8_29_n134 ) : ( n6477 ) ;
assign n6479 =  ( n5809 ) ? ( bv_8_158_n130 ) : ( n6478 ) ;
assign n6480 =  ( n5807 ) ? ( bv_8_225_n123 ) : ( n6479 ) ;
assign n6481 =  ( n5805 ) ? ( bv_8_248_n33 ) : ( n6480 ) ;
assign n6482 =  ( n5803 ) ? ( bv_8_152_n121 ) : ( n6481 ) ;
assign n6483 =  ( n5801 ) ? ( bv_8_17_n117 ) : ( n6482 ) ;
assign n6484 =  ( n5799 ) ? ( bv_8_105_n113 ) : ( n6483 ) ;
assign n6485 =  ( n5797 ) ? ( bv_8_217_n109 ) : ( n6484 ) ;
assign n6486 =  ( n5795 ) ? ( bv_8_142_n105 ) : ( n6485 ) ;
assign n6487 =  ( n5793 ) ? ( bv_8_148_n102 ) : ( n6486 ) ;
assign n6488 =  ( n5791 ) ? ( bv_8_155_n98 ) : ( n6487 ) ;
assign n6489 =  ( n5789 ) ? ( bv_8_30_n94 ) : ( n6488 ) ;
assign n6490 =  ( n5787 ) ? ( bv_8_135_n91 ) : ( n6489 ) ;
assign n6491 =  ( n5785 ) ? ( bv_8_233_n87 ) : ( n6490 ) ;
assign n6492 =  ( n5783 ) ? ( bv_8_206_n83 ) : ( n6491 ) ;
assign n6493 =  ( n5781 ) ? ( bv_8_85_n79 ) : ( n6492 ) ;
assign n6494 =  ( n5779 ) ? ( bv_8_40_n75 ) : ( n6493 ) ;
assign n6495 =  ( n5777 ) ? ( bv_8_223_n71 ) : ( n6494 ) ;
assign n6496 =  ( n5775 ) ? ( bv_8_140_n67 ) : ( n6495 ) ;
assign n6497 =  ( n5773 ) ? ( bv_8_161_n63 ) : ( n6496 ) ;
assign n6498 =  ( n5771 ) ? ( bv_8_137_n59 ) : ( n6497 ) ;
assign n6499 =  ( n5769 ) ? ( bv_8_13_n55 ) : ( n6498 ) ;
assign n6500 =  ( n5767 ) ? ( bv_8_191_n51 ) : ( n6499 ) ;
assign n6501 =  ( n5765 ) ? ( bv_8_230_n47 ) : ( n6500 ) ;
assign n6502 =  ( n5763 ) ? ( bv_8_66_n43 ) : ( n6501 ) ;
assign n6503 =  ( n5761 ) ? ( bv_8_104_n39 ) : ( n6502 ) ;
assign n6504 =  ( n5759 ) ? ( bv_8_65_n35 ) : ( n6503 ) ;
assign n6505 =  ( n5757 ) ? ( bv_8_153_n31 ) : ( n6504 ) ;
assign n6506 =  ( n5755 ) ? ( bv_8_45_n27 ) : ( n6505 ) ;
assign n6507 =  ( n5753 ) ? ( bv_8_15_n23 ) : ( n6506 ) ;
assign n6508 =  ( n5751 ) ? ( bv_8_176_n19 ) : ( n6507 ) ;
assign n6509 =  ( n5749 ) ? ( bv_8_84_n15 ) : ( n6508 ) ;
assign n6510 =  ( n5747 ) ? ( bv_8_187_n11 ) : ( n6509 ) ;
assign n6511 =  ( n5745 ) ? ( bv_8_22_n7 ) : ( n6510 ) ;
assign n6512 =  ( n5743 ) ^ ( n6511 )  ;
assign n6513 =  { ( n5742 ) , ( n6512 ) }  ;
assign n6514 = in[127:120] ;
assign n6515 =  ( n6514 ) ^ ( rcon )  ;
assign n6516 = in[95:88] ;
assign n6517 =  ( n6515 ) ^ ( n6516 )  ;
assign n6518 =  ( n6517 ) ^ ( n4199 )  ;
assign n6519 =  { ( n6513 ) , ( n6518 ) }  ;
assign n6520 = in[119:112] ;
assign n6521 = in[87:80] ;
assign n6522 =  ( n6520 ) ^ ( n6521 )  ;
assign n6523 =  ( n6522 ) ^ ( n4969 )  ;
assign n6524 =  { ( n6519 ) , ( n6523 ) }  ;
assign n6525 = in[111:104] ;
assign n6526 = in[79:72] ;
assign n6527 =  ( n6525 ) ^ ( n6526 )  ;
assign n6528 =  ( n6527 ) ^ ( n5740 )  ;
assign n6529 =  { ( n6524 ) , ( n6528 ) }  ;
assign n6530 = in[103:96] ;
assign n6531 = in[71:64] ;
assign n6532 =  ( n6530 ) ^ ( n6531 )  ;
assign n6533 =  ( n6532 ) ^ ( n6511 )  ;
assign n6534 =  { ( n6529 ) , ( n6533 ) }  ;
assign n6535 = in[127:120] ;
assign n6536 =  ( n6535 ) ^ ( rcon )  ;
assign n6537 = in[95:88] ;
assign n6538 =  ( n6536 ) ^ ( n6537 )  ;
assign n6539 = in[63:56] ;
assign n6540 =  ( n6538 ) ^ ( n6539 )  ;
assign n6541 =  ( n6540 ) ^ ( n4199 )  ;
assign n6542 =  { ( n6534 ) , ( n6541 ) }  ;
assign n6543 = in[119:112] ;
assign n6544 = in[87:80] ;
assign n6545 =  ( n6543 ) ^ ( n6544 )  ;
assign n6546 = in[55:48] ;
assign n6547 =  ( n6545 ) ^ ( n6546 )  ;
assign n6548 =  ( n6547 ) ^ ( n4969 )  ;
assign n6549 =  { ( n6542 ) , ( n6548 ) }  ;
assign n6550 = in[111:104] ;
assign n6551 = in[79:72] ;
assign n6552 =  ( n6550 ) ^ ( n6551 )  ;
assign n6553 = in[47:40] ;
assign n6554 =  ( n6552 ) ^ ( n6553 )  ;
assign n6555 =  ( n6554 ) ^ ( n5740 )  ;
assign n6556 =  { ( n6549 ) , ( n6555 ) }  ;
assign n6557 = in[103:96] ;
assign n6558 = in[71:64] ;
assign n6559 =  ( n6557 ) ^ ( n6558 )  ;
assign n6560 = in[39:32] ;
assign n6561 =  ( n6559 ) ^ ( n6560 )  ;
assign n6562 =  ( n6561 ) ^ ( n6511 )  ;
assign n6563 =  { ( n6556 ) , ( n6562 ) }  ;
assign n6564 = in[127:120] ;
assign n6565 =  ( n6564 ) ^ ( rcon )  ;
assign n6566 = in[95:88] ;
assign n6567 =  ( n6565 ) ^ ( n6566 )  ;
assign n6568 = in[63:56] ;
assign n6569 =  ( n6567 ) ^ ( n6568 )  ;
assign n6570 = in[31:24] ;
assign n6571 =  ( n6569 ) ^ ( n6570 )  ;
assign n6572 =  ( n6571 ) ^ ( n4199 )  ;
assign n6573 =  { ( n6563 ) , ( n6572 ) }  ;
assign n6574 = in[119:112] ;
assign n6575 = in[87:80] ;
assign n6576 =  ( n6574 ) ^ ( n6575 )  ;
assign n6577 = in[55:48] ;
assign n6578 =  ( n6576 ) ^ ( n6577 )  ;
assign n6579 = in[23:16] ;
assign n6580 =  ( n6578 ) ^ ( n6579 )  ;
assign n6581 =  ( n6580 ) ^ ( n4969 )  ;
assign n6582 =  { ( n6573 ) , ( n6581 ) }  ;
assign n6583 = in[111:104] ;
assign n6584 = in[79:72] ;
assign n6585 =  ( n6583 ) ^ ( n6584 )  ;
assign n6586 = in[47:40] ;
assign n6587 =  ( n6585 ) ^ ( n6586 )  ;
assign n6588 = in[15:8] ;
assign n6589 =  ( n6587 ) ^ ( n6588 )  ;
assign n6590 =  ( n6589 ) ^ ( n5740 )  ;
assign n6591 =  { ( n6582 ) , ( n6590 ) }  ;
assign n6592 = in[103:96] ;
assign n6593 = in[71:64] ;
assign n6594 =  ( n6592 ) ^ ( n6593 )  ;
assign n6595 = in[39:32] ;
assign n6596 =  ( n6594 ) ^ ( n6595 )  ;
assign n6597 = in[7:0] ;
assign n6598 =  ( n6596 ) ^ ( n6597 )  ;
assign n6599 =  ( n6598 ) ^ ( n6511 )  ;
assign n6600 =  { ( n6591 ) , ( n6599 ) }  ;
assign n6601 =  ( bv_128_0_n1 ) + ( n6600 )  ;
always @(posedge clk) begin
   if(rst) begin
       in <= in_randinit ;
       rcon <= rcon_randinit ;
       out_1 <= out_1_randinit ;
       out_2 <= out_2_randinit ;
       __COUNTER_start__n0 <= 0;
   end
   else if(__START__ && __ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           in <= in ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           rcon <= rcon ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           out_1 <= n3429 ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           out_2 <= n6601 ;
       end
   end
end
endmodule
