module NV_NVDLA_SDP_CORE_c_core(nvdla_core_clk, nvdla_core_rstn, chn_in_rsc_z, chn_in_rsc_vz, chn_in_rsc_lz, cfg_offset_rsc_z, cfg_scale_rsc_z, cfg_truncate_rsc_z, cfg_proc_precision_rsc_z, cfg_out_precision_rsc_z, cfg_mode_eql_rsc_z, chn_out_rsc_z, chn_out_rsc_vz, chn_out_rsc_lz, chn_in_rsci_oswt, chn_in_rsci_oswt_unreg, chn_out_rsci_oswt, chn_out_rsci_oswt_unreg);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24327" *)
  wire [2:0] _00000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [2:0] _00002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24374" *)
  wire [4:0] _00017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24432" *)
  wire _00074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24449" *)
  wire [9:0] _00106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24466" *)
  wire [14:0] _00138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24500" *)
  wire [23:0] _00170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24647" *)
  wire [10:0] _00186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24641" *)
  wire [2:0] _00202_;
  wire [15:0] _00203_;
  wire [15:0] _00204_;
  wire [15:0] _00205_;
  wire [15:0] _00206_;
  wire [15:0] _00207_;
  wire [15:0] _00208_;
  wire [15:0] _00209_;
  wire [15:0] _00210_;
  wire [15:0] _00211_;
  wire [15:0] _00212_;
  wire [15:0] _00213_;
  wire [15:0] _00214_;
  wire [15:0] _00215_;
  wire [15:0] _00216_;
  wire [15:0] _00217_;
  wire [15:0] _00218_;
  wire [3:0] _00219_;
  wire [3:0] _00220_;
  wire [3:0] _00221_;
  wire [3:0] _00222_;
  wire [3:0] _00223_;
  wire [3:0] _00224_;
  wire [3:0] _00225_;
  wire [3:0] _00226_;
  wire [3:0] _00227_;
  wire [3:0] _00228_;
  wire [3:0] _00229_;
  wire [3:0] _00230_;
  wire [3:0] _00231_;
  wire [3:0] _00232_;
  wire [3:0] _00233_;
  wire [3:0] _00234_;
  wire [3:0] _00235_;
  wire [3:0] _00236_;
  wire [3:0] _00237_;
  wire [3:0] _00238_;
  wire [3:0] _00239_;
  wire [3:0] _00240_;
  wire [3:0] _00241_;
  wire [3:0] _00242_;
  wire [3:0] _00243_;
  wire [3:0] _00244_;
  wire [3:0] _00245_;
  wire [3:0] _00246_;
  wire [3:0] _00247_;
  wire [3:0] _00248_;
  wire [3:0] _00249_;
  wire [3:0] _00250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17958" *)
  wire _00265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18365" *)
  wire _00266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18300" *)
  wire [14:0] _00267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire [9:0] _00268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17565" *)
  wire _00269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17613" *)
  wire _00270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17671" *)
  wire _00271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17719" *)
  wire _00272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17786" *)
  wire _00273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17842" *)
  wire _00274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16983" *)
  wire _00275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17041" *)
  wire _00276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17105" *)
  wire _00277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17205" *)
  wire _00278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17261" *)
  wire _00279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17329" *)
  wire _00280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17391" *)
  wire _00281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17447" *)
  wire _00282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17505" *)
  wire _00283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17898" *)
  wire _00284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16983" *)
  wire [14:0] _00285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17041" *)
  wire [14:0] _00286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17105" *)
  wire [14:0] _00287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17505" *)
  wire [14:0] _00288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20835" *)
  wire _00289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21020" *)
  wire _00290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21039" *)
  wire _00291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21059" *)
  wire _00292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21079" *)
  wire _00293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21098" *)
  wire _00294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21116" *)
  wire _00295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20853" *)
  wire _00296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20871" *)
  wire _00297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20889" *)
  wire _00298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20908" *)
  wire _00299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20927" *)
  wire _00300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20945" *)
  wire _00301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20964" *)
  wire _00302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20983" *)
  wire _00303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21002" *)
  wire _00304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _00305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19295" *)
  wire _00306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _00307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19325" *)
  wire _00308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19591" *)
  wire _00309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19356" *)
  wire _00310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21147" *)
  wire _00311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19387" *)
  wire _00312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19603" *)
  wire _00313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19387" *)
  wire _00314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19614" *)
  wire _00315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19474" *)
  wire _00316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18983" *)
  wire _00317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19023" *)
  wire _00318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19054" *)
  wire _00319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _00320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19099" *)
  wire _00321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19054" *)
  wire _00322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _00323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19161" *)
  wire _00324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _00325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19192" *)
  wire _00326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19591" *)
  wire _00327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19223" *)
  wire _00328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19254" *)
  wire _00329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19614" *)
  wire _00330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19474" *)
  wire _00331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19953" *)
  wire [4:0] _00332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19969" *)
  wire [4:0] _00333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19985" *)
  wire [4:0] _00334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20001" *)
  wire [4:0] _00335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20017" *)
  wire [4:0] _00336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20033" *)
  wire [4:0] _00337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19809" *)
  wire [4:0] _00338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19825" *)
  wire [4:0] _00339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19841" *)
  wire [4:0] _00340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19857" *)
  wire [4:0] _00341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19873" *)
  wire [4:0] _00342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19889" *)
  wire [4:0] _00343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19905" *)
  wire [4:0] _00344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19921" *)
  wire [4:0] _00345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19937" *)
  wire [4:0] _00346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20049" *)
  wire [4:0] _00347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19961" *)
  wire _00348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19977" *)
  wire _00349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19993" *)
  wire _00350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20009" *)
  wire _00351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20025" *)
  wire _00352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20041" *)
  wire _00353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19817" *)
  wire _00354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19833" *)
  wire _00355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19849" *)
  wire _00356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19865" *)
  wire _00357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19881" *)
  wire _00358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19897" *)
  wire _00359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19913" *)
  wire _00360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19929" *)
  wire _00361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19945" *)
  wire _00362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20057" *)
  wire _00363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15909" *)
  wire [2:0] _00364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15937" *)
  wire [2:0] _00365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15965" *)
  wire [2:0] _00366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15993" *)
  wire [2:0] _00367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16021" *)
  wire [2:0] _00368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16049" *)
  wire [2:0] _00369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16077" *)
  wire [2:0] _00370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16105" *)
  wire [2:0] _00371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15633" *)
  wire [2:0] _00372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15669" *)
  wire [2:0] _00373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15741" *)
  wire [2:0] _00374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15769" *)
  wire [2:0] _00375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15797" *)
  wire [2:0] _00376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15825" *)
  wire [2:0] _00377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15853" *)
  wire [2:0] _00378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15881" *)
  wire [2:0] _00379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15955" *)
  wire _00381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15983" *)
  wire _00383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16011" *)
  wire _00385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16039" *)
  wire _00387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16067" *)
  wire _00389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16095" *)
  wire _00391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15659" *)
  wire _00393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15731" *)
  wire _00395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15759" *)
  wire _00397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15787" *)
  wire _00399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15815" *)
  wire _00401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15843" *)
  wire _00403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15871" *)
  wire _00405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15899" *)
  wire _00407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15927" *)
  wire _00409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16123" *)
  wire _00411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20179" *)
  wire [4:0] _00430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20160" *)
  wire [4:0] _00433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20141" *)
  wire [4:0] _00436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20122" *)
  wire [4:0] _00439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20103" *)
  wire [4:0] _00442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20084" *)
  wire [4:0] _00445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20350" *)
  wire [4:0] _00448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20331" *)
  wire [4:0] _00451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20312" *)
  wire [4:0] _00454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20293" *)
  wire [4:0] _00457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20274" *)
  wire [4:0] _00460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20255" *)
  wire [4:0] _00463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20236" *)
  wire [4:0] _00466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20217" *)
  wire [4:0] _00469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20198" *)
  wire [4:0] _00472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [3:0] _00473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20065" *)
  wire [4:0] _00475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16872" *)
  wire [9:0] _00476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16883" *)
  wire [9:0] _00477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16894" *)
  wire [9:0] _00478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16905" *)
  wire [9:0] _00479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16916" *)
  wire [9:0] _00480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16927" *)
  wire [9:0] _00481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16713" *)
  wire [9:0] _00482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16732" *)
  wire [9:0] _00483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16755" *)
  wire [9:0] _00484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16766" *)
  wire [9:0] _00485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16777" *)
  wire [9:0] _00486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16796" *)
  wire [9:0] _00487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16827" *)
  wire [9:0] _00488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16838" *)
  wire [9:0] _00489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16849" *)
  wire [9:0] _00490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16946" *)
  wire [9:0] _00491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16507" *)
  wire [48:0] _00498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16429" *)
  wire [48:0] _00499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16429" *)
  wire [48:0] _00500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16444" *)
  wire [48:0] _00501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16490" *)
  wire [48:0] _00502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16429" *)
  wire [48:0] _00506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _00507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19761" *)
  wire _00511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17747" *)
  wire _00512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19428" *)
  wire _00513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20561" *)
  wire _00526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20441" *)
  wire [14:0] _00527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20429" *)
  wire [14:0] _00528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20417" *)
  wire [14:0] _00529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20405" *)
  wire [14:0] _00530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20393" *)
  wire [14:0] _00531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20381" *)
  wire [14:0] _00532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20549" *)
  wire [14:0] _00533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20537" *)
  wire [14:0] _00534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20525" *)
  wire [14:0] _00535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20513" *)
  wire [14:0] _00536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20501" *)
  wire [14:0] _00537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20489" *)
  wire [14:0] _00538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20477" *)
  wire [14:0] _00539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20465" *)
  wire [14:0] _00540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20453" *)
  wire [14:0] _00541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20369" *)
  wire [14:0] _00542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17537" *)
  wire [48:0] _00543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17585" *)
  wire [48:0] _00544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17633" *)
  wire [48:0] _00545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17691" *)
  wire [48:0] _00546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17739" *)
  wire [48:0] _00547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17806" *)
  wire [48:0] _00548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16965" *)
  wire [48:0] _00549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17013" *)
  wire [48:0] _00550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17087" *)
  wire [48:0] _00551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17137" *)
  wire [48:0] _00552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17235" *)
  wire [48:0] _00553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17291" *)
  wire [48:0] _00554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17363" *)
  wire [48:0] _00555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17411" *)
  wire [48:0] _00556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17487" *)
  wire [48:0] _00557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17862" *)
  wire [48:0] _00558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20804" *)
  wire _00559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20743" *)
  wire _00560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20743" *)
  wire _00561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20757" *)
  wire _00562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20768" *)
  wire _00563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20768" *)
  wire _00564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20793" *)
  wire _00565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20815" *)
  wire _00566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20682" *)
  wire _00567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20682" *)
  wire _00568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20696" *)
  wire _00569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20732" *)
  wire _00570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20707" *)
  wire _00571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20707" *)
  wire _00572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20721" *)
  wire _00573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20782" *)
  wire _00574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19420" *)
  wire _00583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18971" *)
  wire _00590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18971" *)
  wire _00594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18971" *)
  wire _00602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire [14:0] _00605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17555" *)
  wire [14:0] _00606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire [14:0] _00607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17603" *)
  wire [14:0] _00608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19751" *)
  wire [14:0] _00609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17651" *)
  wire [14:0] _00610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19761" *)
  wire [14:0] _00611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17709" *)
  wire [14:0] _00612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19761" *)
  wire [14:0] _00613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17759" *)
  wire [14:0] _00614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19781" *)
  wire [14:0] _00615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17824" *)
  wire [14:0] _00616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21157" *)
  wire [14:0] _00617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16973" *)
  wire [14:0] _00618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire [14:0] _00619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17031" *)
  wire [14:0] _00620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire [14:0] _00621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17095" *)
  wire [14:0] _00622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19761" *)
  wire [14:0] _00623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17155" *)
  wire [14:0] _00624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21184" *)
  wire [14:0] _00625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17243" *)
  wire [14:0] _00626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19705" *)
  wire [14:0] _00627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17309" *)
  wire [14:0] _00628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19705" *)
  wire [14:0] _00629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17381" *)
  wire [14:0] _00630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19719" *)
  wire [14:0] _00631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17429" *)
  wire [14:0] _00632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire [14:0] _00633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17495" *)
  wire [14:0] _00634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19791" *)
  wire [14:0] _00635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17880" *)
  wire [14:0] _00636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire _00637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17545" *)
  wire _00638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire _00640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17593" *)
  wire _00641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19751" *)
  wire _00643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17641" *)
  wire _00644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19761" *)
  wire _00646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17699" *)
  wire _00647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19761" *)
  wire _00649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17747" *)
  wire _00650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19781" *)
  wire _00652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17814" *)
  wire _00653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18806" *)
  wire _00656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19729" *)
  wire _00657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17021" *)
  wire _00658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18887" *)
  wire _00661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19761" *)
  wire _00662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17145" *)
  wire _00663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18904" *)
  wire _00666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19705" *)
  wire _00667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17299" *)
  wire _00668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19705" *)
  wire _00670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17371" *)
  wire _00671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19719" *)
  wire _00673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17419" *)
  wire _00674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18963" *)
  wire _00677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19791" *)
  wire _00678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17870" *)
  wire _00679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20671" *)
  wire _00681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20651" *)
  wire _00682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20630" *)
  wire _00683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18553" *)
  wire _00693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18115" *)
  wire _00694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18115" *)
  wire _00695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18153" *)
  wire _00696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18528" *)
  wire _00706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _00712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20661" *)
  wire _00713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20641" *)
  wire _00714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20620" *)
  wire _00715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire _00733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _00734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire [1:0] _00736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [1:0] _00737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19554" *)
  wire [1:0] _00738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19544" *)
  wire [1:0] _00739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17918" *)
  wire [1:0] _00740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16499" *)
  wire [1:0] _00741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19528" *)
  wire [1:0] _00742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17926" *)
  wire [1:0] _00743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19544" *)
  wire [1:0] _00744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19536" *)
  wire [1:0] _00745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [1:0] _00746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [1:0] _00747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire [1:0] _00748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17938" *)
  wire [1:0] _00749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19554" *)
  wire [1:0] _00750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [5:0] _00751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15641" *)
  wire [27:0] _00757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19801" *)
  wire _00766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire [28:0] _00768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20612" *)
  wire [15:0] _00771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16938" *)
  wire _00784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire [16:0] _00785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18195" *)
  wire [16:0] _00786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18292" *)
  wire [16:0] _00787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18357" *)
  wire [16:0] _00788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18434" *)
  wire [16:0] _00789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18520" *)
  wire [16:0] _00790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18600" *)
  wire [16:0] _00791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18648" *)
  wire [16:0] _00792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18672" *)
  wire [16:0] _00793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18624" *)
  wire [16:0] _00794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18579" *)
  wire [16:0] _00795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18499" *)
  wire [16:0] _00796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18410" *)
  wire [16:0] _00797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18037" *)
  wire [16:0] _00798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18336" *)
  wire [16:0] _00799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18145" *)
  wire [16:0] _00800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15088" *)
  wire _00801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15098" *)
  wire _00802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18955" *)
  wire _00803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15406" *)
  wire [3:0] _00806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15420" *)
  wire [3:0] _00811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15106" *)
  wire [3:0] _00816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15106" *)
  wire [3:0] _00817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15434" *)
  wire [3:0] _00823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15448" *)
  wire [3:0] _00830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15462" *)
  wire [3:0] _00835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15476" *)
  wire [3:0] _00840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15490" *)
  wire [3:0] _00845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15510" *)
  wire [3:0] _00850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15605" *)
  wire _00853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15490" *)
  wire [3:0] _00855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15605" *)
  wire _00857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15365" *)
  wire [3:0] _00875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15106" *)
  wire [3:0] _00880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15379" *)
  wire [3:0] _00885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15106" *)
  wire [3:0] _00890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15392" *)
  wire [3:0] _00895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire _00896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _00898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15136" *)
  wire [8:0] _00899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15088" *)
  wire _00900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18680" *)
  wire _00901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16807" *)
  wire [4:0] _00903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21211" *)
  wire _00904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _00905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17575" *)
  wire _00906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20993" *)
  wire _00907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21346" *)
  wire _00908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20187" *)
  wire _00909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15945" *)
  wire _00911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18696" *)
  wire _00914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16807" *)
  wire [4:0] _00916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21211" *)
  wire _00917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _00918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17623" *)
  wire _00919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21011" *)
  wire _00920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21356" *)
  wire _00921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20168" *)
  wire _00922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15973" *)
  wire _00924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18656" *)
  wire _00927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16860" *)
  wire [4:0] _00929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21221" *)
  wire _00930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19668" *)
  wire _00931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17681" *)
  wire _00932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21029" *)
  wire _00933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21366" *)
  wire _00934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20149" *)
  wire _00935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16001" *)
  wire _00937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18608" *)
  wire _00940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16807" *)
  wire [4:0] _00942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21165" *)
  wire _00943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19680" *)
  wire _00944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17729" *)
  wire _00945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21049" *)
  wire _00946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21376" *)
  wire _00947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20130" *)
  wire _00948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16029" *)
  wire _00950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18537" *)
  wire _00953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16860" *)
  wire [4:0] _00955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21230" *)
  wire _00956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19695" *)
  wire _00957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17796" *)
  wire _00958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21069" *)
  wire _00959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21386" *)
  wire _00960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20111" *)
  wire _00961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16057" *)
  wire _00963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18814" *)
  wire _00965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18468" *)
  wire _00967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16807" *)
  wire [4:0] _00969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21238" *)
  wire _00970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19680" *)
  wire _00971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17852" *)
  wire _00972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21088" *)
  wire _00973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21396" *)
  wire _00974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20092" *)
  wire _00975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16085" *)
  wire _00977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18374" *)
  wire _00980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16957" *)
  wire [4:0] _00982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21247" *)
  wire _00983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19680" *)
  wire _00984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17908" *)
  wire _00985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21107" *)
  wire _00986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21406" *)
  wire _00987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20073" *)
  wire _00988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16113" *)
  wire _00990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _00991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _00992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18024" *)
  wire _00993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _00994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16724" *)
  wire [4:0] _00995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17005" *)
  wire _00996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16995" *)
  wire _00997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20826" *)
  wire _00998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21256" *)
  wire _00999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20358" *)
  wire _01000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15649" *)
  wire _01002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19013" *)
  wire _01004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17938" *)
  wire _01006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18129" *)
  wire _01007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16743" *)
  wire [4:0] _01009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19626" *)
  wire _01010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17063" *)
  wire _01011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17053" *)
  wire _01012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20844" *)
  wire _01013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21266" *)
  wire _01014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20339" *)
  wire _01015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15721" *)
  wire _01017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17073" *)
  wire _01020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18179" *)
  wire _01021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16743" *)
  wire [4:0] _01023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19626" *)
  wire _01024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17127" *)
  wire _01025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17117" *)
  wire _01026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20862" *)
  wire _01027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21276" *)
  wire _01028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20320" *)
  wire _01029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15749" *)
  wire _01031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19089" *)
  wire _01033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17073" *)
  wire _01035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18276" *)
  wire _01036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16743" *)
  wire [4:0] _01038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21165" *)
  wire _01039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17215" *)
  wire _01041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20880" *)
  wire _01042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21286" *)
  wire _01043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20301" *)
  wire _01044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15777" *)
  wire _01046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17225" *)
  wire _01049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18344" *)
  wire _01050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16788" *)
  wire [4:0] _01052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21175" *)
  wire _01053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19659" *)
  wire _01054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17281" *)
  wire _01055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17271" *)
  wire _01056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20898" *)
  wire _01057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21296" *)
  wire _01058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20282" *)
  wire _01059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15805" *)
  wire _01061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19151" *)
  wire _01063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17477" *)
  wire _01065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18418" *)
  wire _01066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16807" *)
  wire [4:0] _01068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21192" *)
  wire _01069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17339" *)
  wire _01071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20918" *)
  wire _01072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21306" *)
  wire _01073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20263" *)
  wire _01074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15833" *)
  wire _01076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17349" *)
  wire _01079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18507" *)
  wire _01080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16807" *)
  wire [4:0] _01082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21192" *)
  wire _01083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17401" *)
  wire _01085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20936" *)
  wire _01086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21316" *)
  wire _01087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20244" *)
  wire _01088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15861" *)
  wire _01090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17349" *)
  wire _01093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18587" *)
  wire _01094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16807" *)
  wire [4:0] _01096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21202" *)
  wire _01097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19668" *)
  wire _01098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17457" *)
  wire _01099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20954" *)
  wire _01100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21326" *)
  wire _01101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20225" *)
  wire _01102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15889" *)
  wire _01104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17467" *)
  wire _01107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18632" *)
  wire _01108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18045" *)
  wire _01109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16860" *)
  wire [4:0] _01110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19626" *)
  wire _01111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17527" *)
  wire _01112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17517" *)
  wire _01113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20973" *)
  wire _01114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21336" *)
  wire _01115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20206" *)
  wire _01116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15917" *)
  wire _01118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16133" *)
  wire _01119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19285" *)
  wire _01120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17926" *)
  wire _01122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18895" *)
  wire _01123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18912" *)
  wire _01124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18922" *)
  wire _01125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18922" *)
  wire _01126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18943" *)
  wire _01127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18943" *)
  wire _01128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18868" *)
  wire _01129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18878" *)
  wire _01130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18934" *)
  wire _01131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18922" *)
  wire _01132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18943" *)
  wire _01133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18868" *)
  wire _01134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15677" *)
  wire _01135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16526" *)
  wire _01136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18712" *)
  wire _01137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15625" *)
  wire _01138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16518" *)
  wire _01139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17950" *)
  wire _01140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18454" *)
  wire [9:0] _01141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18314" *)
  wire [4:0] _01142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18454" *)
  wire [9:0] _01143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18314" *)
  wire [4:0] _01144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18400" *)
  wire [9:0] _01145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18390" *)
  wire [4:0] _01146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18571" *)
  wire [9:0] _01147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18563" *)
  wire [4:0] _01148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18490" *)
  wire [9:0] _01149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18481" *)
  wire [4:0] _01150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18400" *)
  wire [9:0] _01151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18390" *)
  wire [4:0] _01152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18170" *)
  wire [9:0] _01153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18162" *)
  wire [4:0] _01154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18264" *)
  wire [9:0] _01155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18252" *)
  wire [4:0] _01156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18264" *)
  wire [9:0] _01157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18252" *)
  wire [4:0] _01158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18454" *)
  wire [9:0] _01159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18442" *)
  wire [4:0] _01160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18454" *)
  wire [9:0] _01161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18442" *)
  wire [4:0] _01162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18326" *)
  wire [9:0] _01163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18442" *)
  wire [4:0] _01164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18264" *)
  wire [9:0] _01165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18252" *)
  wire [4:0] _01166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18326" *)
  wire [9:0] _01167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18314" *)
  wire [4:0] _01168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17193" *)
  wire [9:0] _01169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17193" *)
  wire [9:0] _01171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17661" *)
  wire [9:0] _01173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17661" *)
  wire [9:0] _01175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17778" *)
  wire [9:0] _01177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17769" *)
  wire [4:0] _01178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17834" *)
  wire [9:0] _01179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17193" *)
  wire [9:0] _01181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17253" *)
  wire [9:0] _01183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17319" *)
  wire [9:0] _01185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17319" *)
  wire [9:0] _01187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17439" *)
  wire [9:0] _01189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17890" *)
  wire [9:0] _01191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17165" *)
  wire [4:0] _01192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19316" *)
  wire [3:0] _01193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19304" *)
  wire _01194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19347" *)
  wire [3:0] _01195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19335" *)
  wire _01196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19378" *)
  wire [3:0] _01197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19366" *)
  wire _01198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19411" *)
  wire [3:0] _01199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19399" *)
  wire _01200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19448" *)
  wire [3:0] _01201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19436" *)
  wire _01202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19498" *)
  wire [3:0] _01203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19486" *)
  wire _01204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19004" *)
  wire [3:0] _01205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18993" *)
  wire _01206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19045" *)
  wire [3:0] _01207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19033" *)
  wire _01208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19080" *)
  wire [3:0] _01209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19068" *)
  wire _01210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19121" *)
  wire [3:0] _01211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19109" *)
  wire _01212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19142" *)
  wire [3:0] _01213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19130" *)
  wire _01214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19183" *)
  wire [3:0] _01215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19171" *)
  wire _01216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19214" *)
  wire [3:0] _01217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19202" *)
  wire _01218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19245" *)
  wire [3:0] _01219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19233" *)
  wire _01220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19276" *)
  wire [3:0] _01221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19264" *)
  wire _01222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19519" *)
  wire [3:0] _01223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19507" *)
  wire _01224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19457" *)
  wire [4:0] _01225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19466" *)
  wire [9:0] _01226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16507" *)
  wire [1:0] _01227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19572" *)
  wire [4:0] _01228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19582" *)
  wire [9:0] _01229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19564" *)
  wire _01230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15617" *)
  wire _01231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18912" *)
  wire _01232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15524" *)
  wire _01262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15605" *)
  wire _01263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15605" *)
  wire _01264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16983" *)
  wire _01265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17021" *)
  wire _01266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17041" *)
  wire _01267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17105" *)
  wire _01268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17145" *)
  wire _01269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17205" *)
  wire _01270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17261" *)
  wire _01271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17299" *)
  wire _01272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17329" *)
  wire _01273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17371" *)
  wire _01274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17391" *)
  wire _01275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17419" *)
  wire _01276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17447" *)
  wire _01277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17505" *)
  wire _01278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17545" *)
  wire _01279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17565" *)
  wire _01280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17593" *)
  wire _01281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17613" *)
  wire _01282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17641" *)
  wire _01283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17671" *)
  wire _01284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17699" *)
  wire _01285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17719" *)
  wire _01286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17747" *)
  wire _01287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17747" *)
  wire _01288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17786" *)
  wire _01289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17814" *)
  wire _01290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17842" *)
  wire _01291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17870" *)
  wire _01292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17898" *)
  wire _01293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18115" *)
  wire _01294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18115" *)
  wire _01295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18153" *)
  wire _01296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire _01308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18365" *)
  wire _01309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18528" *)
  wire _01310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18553" *)
  wire _01311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19023" *)
  wire _01312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19099" *)
  wire _01313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19161" *)
  wire _01314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19192" *)
  wire _01315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19223" *)
  wire _01316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19295" *)
  wire _01317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19325" *)
  wire _01318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19356" *)
  wire _01319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19387" *)
  wire _01320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19387" *)
  wire _01321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19474" *)
  wire _01322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19474" *)
  wire _01323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19591" *)
  wire _01324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19591" *)
  wire _01325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19603" *)
  wire _01326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19614" *)
  wire _01327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19614" *)
  wire _01328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19638" *)
  wire _01333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19659" *)
  wire _01334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19668" *)
  wire _01335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19668" *)
  wire _01336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19680" *)
  wire _01337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19680" *)
  wire _01338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19680" *)
  wire _01339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19695" *)
  wire _01340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20073" *)
  wire _01341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20092" *)
  wire _01342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20111" *)
  wire _01343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20130" *)
  wire _01344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20149" *)
  wire _01345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20168" *)
  wire _01346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20187" *)
  wire _01347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20206" *)
  wire _01348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20225" *)
  wire _01349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20244" *)
  wire _01350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20263" *)
  wire _01351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20282" *)
  wire _01352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20301" *)
  wire _01353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20320" *)
  wire _01354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20339" *)
  wire _01355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20358" *)
  wire _01356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20620" *)
  wire _01357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20630" *)
  wire _01358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20641" *)
  wire _01359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20651" *)
  wire _01360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20661" *)
  wire _01361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20671" *)
  wire _01362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20682" *)
  wire _01363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20682" *)
  wire _01364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20696" *)
  wire _01365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20707" *)
  wire _01366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20707" *)
  wire _01367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20721" *)
  wire _01368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20732" *)
  wire _01369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20743" *)
  wire _01370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20743" *)
  wire _01371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20757" *)
  wire _01372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20768" *)
  wire _01373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20768" *)
  wire _01374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20782" *)
  wire _01375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20793" *)
  wire _01376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20804" *)
  wire _01377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20815" *)
  wire _01378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _01379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _01380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _01381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _01382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21126" *)
  wire _01383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21147" *)
  wire _01384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16713" *)
  wire [9:0] _01385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16732" *)
  wire [9:0] _01386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16755" *)
  wire [9:0] _01387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16766" *)
  wire [9:0] _01388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16777" *)
  wire [9:0] _01389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16796" *)
  wire [9:0] _01390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16827" *)
  wire [9:0] _01391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16838" *)
  wire [9:0] _01392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16849" *)
  wire [9:0] _01393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16872" *)
  wire [9:0] _01394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16883" *)
  wire [9:0] _01395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16894" *)
  wire [9:0] _01396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16905" *)
  wire [9:0] _01397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16916" *)
  wire [9:0] _01398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16927" *)
  wire [9:0] _01399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16946" *)
  wire [9:0] _01400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18203" *)
  wire [9:0] _01401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16973" *)
  wire [14:0] _01402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16983" *)
  wire [14:0] _01403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17031" *)
  wire [14:0] _01404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17041" *)
  wire [14:0] _01405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17095" *)
  wire [14:0] _01406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17105" *)
  wire [14:0] _01407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17155" *)
  wire [14:0] _01408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17243" *)
  wire [14:0] _01409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17309" *)
  wire [14:0] _01410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17381" *)
  wire [14:0] _01411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17429" *)
  wire [14:0] _01412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17495" *)
  wire [14:0] _01413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17505" *)
  wire [14:0] _01414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17555" *)
  wire [14:0] _01415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17603" *)
  wire [14:0] _01416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17651" *)
  wire [14:0] _01417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17709" *)
  wire [14:0] _01418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17759" *)
  wire [14:0] _01419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17824" *)
  wire [14:0] _01420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17880" *)
  wire [14:0] _01421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16444" *)
  wire [48:0] _01422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16454" *)
  wire [48:0] _01432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10004" *)
  wire _01433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10010" *)
  wire _01434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10016" *)
  wire _01435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10022" *)
  wire _01436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10028" *)
  wire _01437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10034" *)
  wire _01438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10040" *)
  wire _01439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10046" *)
  wire _01440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10052" *)
  wire _01441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10058" *)
  wire _01442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10071" *)
  wire _01443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10071" *)
  wire _01444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10071" *)
  wire _01445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10075" *)
  wire _01446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10079" *)
  wire _01447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10079" *)
  wire _01448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10084" *)
  wire _01449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *)
  wire _01450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *)
  wire _01451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *)
  wire _01452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *)
  wire _01453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *)
  wire _01454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *)
  wire _01455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *)
  wire _01456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10094" *)
  wire _01457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10094" *)
  wire _01458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10104" *)
  wire _01459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10110" *)
  wire _01460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10125" *)
  wire _01461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11235" *)
  wire _01462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11261" *)
  wire _01463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11261" *)
  wire _01464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11281" *)
  wire _01465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11281" *)
  wire _01466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11295" *)
  wire _01467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11295" *)
  wire _01468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11309" *)
  wire _01469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11309" *)
  wire _01470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11323" *)
  wire _01471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11323" *)
  wire _01472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11337" *)
  wire _01473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11337" *)
  wire _01474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11351" *)
  wire _01475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11351" *)
  wire _01476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11365" *)
  wire _01477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11365" *)
  wire _01478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11379" *)
  wire _01479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11379" *)
  wire _01480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11393" *)
  wire _01481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11393" *)
  wire _01482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11407" *)
  wire _01483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11407" *)
  wire _01484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11639" *)
  wire _01485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11645" *)
  wire _01486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11651" *)
  wire _01487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11657" *)
  wire _01488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11663" *)
  wire _01489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11669" *)
  wire _01490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11675" *)
  wire _01491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11681" *)
  wire _01492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11687" *)
  wire _01493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11693" *)
  wire _01494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11700" *)
  wire _01495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11707" *)
  wire _01496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11714" *)
  wire _01497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11721" *)
  wire _01498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11728" *)
  wire _01499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11735" *)
  wire _01500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11738" *)
  wire _01501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11759" *)
  wire _01502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11765" *)
  wire _01503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11771" *)
  wire _01504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11777" *)
  wire _01505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11783" *)
  wire _01506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11789" *)
  wire _01507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11795" *)
  wire _01508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11801" *)
  wire _01509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11810" *)
  wire _01510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11816" *)
  wire _01511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11825" *)
  wire _01512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11831" *)
  wire _01513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11837" *)
  wire _01514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11843" *)
  wire _01515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11849" *)
  wire _01516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11855" *)
  wire _01517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14072" *)
  wire _01518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14073" *)
  wire _01519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14074" *)
  wire _01520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14075" *)
  wire _01521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14076" *)
  wire _01522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14077" *)
  wire _01523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14078" *)
  wire _01524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14079" *)
  wire _01525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14080" *)
  wire _01526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14081" *)
  wire _01527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14082" *)
  wire _01528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14083" *)
  wire _01529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14084" *)
  wire _01530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14085" *)
  wire _01531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14086" *)
  wire _01532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14087" *)
  wire _01533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14088" *)
  wire _01534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14089" *)
  wire _01535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14090" *)
  wire _01536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14093" *)
  wire _01537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14094" *)
  wire _01538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14095" *)
  wire _01539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14096" *)
  wire _01540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14097" *)
  wire _01541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14127" *)
  wire _01542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14145" *)
  wire _01543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14156" *)
  wire _01544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14172" *)
  wire _01545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14174" *)
  wire _01546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14180" *)
  wire _01547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14200" *)
  wire _01548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14203" *)
  wire _01549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14209" *)
  wire _01550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14232" *)
  wire _01551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14241" *)
  wire _01552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14246" *)
  wire _01553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14257" *)
  wire _01554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14261" *)
  wire _01555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14275" *)
  wire _01556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14281" *)
  wire _01557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14297" *)
  wire _01558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14298" *)
  wire _01559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14308" *)
  wire _01560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14312" *)
  wire _01561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14325" *)
  wire _01562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14329" *)
  wire _01563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14342" *)
  wire _01564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14346" *)
  wire _01565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14364" *)
  wire _01566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14373" *)
  wire _01567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14412" *)
  wire _01568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14440" *)
  wire _01569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14473" *)
  wire _01570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14473" *)
  wire _01571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14494" *)
  wire _01572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14507" *)
  wire _01573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14540" *)
  wire _01574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14561" *)
  wire _01575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14616" *)
  wire _01576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14656" *)
  wire _01577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14656" *)
  wire _01578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14677" *)
  wire _01579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14678" *)
  wire _01580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14680" *)
  wire _01581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14684" *)
  wire _01582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14702" *)
  wire _01583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14736" *)
  wire _01584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14737" *)
  wire _01585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14741" *)
  wire _01586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14743" *)
  wire _01587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14749" *)
  wire _01588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14750" *)
  wire _01589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14752" *)
  wire _01590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14767" *)
  wire _01591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14778" *)
  wire _01592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14778" *)
  wire _01593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14778" *)
  wire _01594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14781" *)
  wire _01595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14782" *)
  wire _01596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14782" *)
  wire _01597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14783" *)
  wire _01598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14784" *)
  wire _01599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14784" *)
  wire _01600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14784" *)
  wire _01601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14853" *)
  wire _01602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14854" *)
  wire _01603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14855" *)
  wire _01604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14855" *)
  wire _01605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14856" *)
  wire _01606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14857" *)
  wire _01607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14863" *)
  wire _01608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14870" *)
  wire _01609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14877" *)
  wire _01610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14881" *)
  wire _01611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14881" *)
  wire _01612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14887" *)
  wire _01613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14894" *)
  wire _01614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14901" *)
  wire _01615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14908" *)
  wire _01616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14915" *)
  wire _01617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14922" *)
  wire _01618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14929" *)
  wire _01619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14936" *)
  wire _01620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14990" *)
  wire _01621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15057" *)
  wire _01622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15057" *)
  wire _01623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15059" *)
  wire _01624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15059" *)
  wire _01625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15061" *)
  wire _01626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15061" *)
  wire _01627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15063" *)
  wire _01628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15063" *)
  wire _01629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15065" *)
  wire _01630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15065" *)
  wire _01631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15067" *)
  wire _01632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15067" *)
  wire _01633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15069" *)
  wire _01634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15069" *)
  wire _01635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15071" *)
  wire _01636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15071" *)
  wire _01637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15073" *)
  wire _01638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15073" *)
  wire _01639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15075" *)
  wire _01640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15075" *)
  wire _01641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15077" *)
  wire _01642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15077" *)
  wire _01643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15079" *)
  wire _01644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15079" *)
  wire _01645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15081" *)
  wire _01646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15081" *)
  wire _01647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15083" *)
  wire _01648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15083" *)
  wire _01649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15085" *)
  wire _01650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15085" *)
  wire _01651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15087" *)
  wire _01652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15087" *)
  wire _01653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15094" *)
  wire _01654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15102" *)
  wire _01655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15332" *)
  wire _01656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15334" *)
  wire _01657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15336" *)
  wire _01658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15338" *)
  wire _01659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15340" *)
  wire _01660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15342" *)
  wire _01661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15344" *)
  wire _01662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15346" *)
  wire _01663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15348" *)
  wire _01664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15350" *)
  wire _01665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15352" *)
  wire _01666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15354" *)
  wire _01667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15356" *)
  wire _01668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15358" *)
  wire _01669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15360" *)
  wire _01670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15362" *)
  wire _01671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15370" *)
  wire _01672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15370" *)
  wire _01673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15384" *)
  wire _01674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15384" *)
  wire _01675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15397" *)
  wire _01676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15397" *)
  wire _01677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15411" *)
  wire _01678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15411" *)
  wire _01679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15425" *)
  wire _01680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15425" *)
  wire _01681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15439" *)
  wire _01682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15439" *)
  wire _01683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15453" *)
  wire _01684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15453" *)
  wire _01685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15467" *)
  wire _01686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15467" *)
  wire _01687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15481" *)
  wire _01688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15481" *)
  wire _01689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15515" *)
  wire _01690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15515" *)
  wire _01691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15621" *)
  wire _01692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15629" *)
  wire _01693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15637" *)
  wire _01694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15645" *)
  wire _01695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15654" *)
  wire _01696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15664" *)
  wire _01697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15673" *)
  wire _01698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15726" *)
  wire _01699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15736" *)
  wire _01700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15745" *)
  wire _01701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15754" *)
  wire _01702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15764" *)
  wire _01703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15773" *)
  wire _01704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15782" *)
  wire _01705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15792" *)
  wire _01706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15801" *)
  wire _01707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15810" *)
  wire _01708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15820" *)
  wire _01709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15829" *)
  wire _01710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15838" *)
  wire _01711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15848" *)
  wire _01712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15857" *)
  wire _01713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15866" *)
  wire _01714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15876" *)
  wire _01715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15885" *)
  wire _01716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15894" *)
  wire _01717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15904" *)
  wire _01718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15913" *)
  wire _01719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15922" *)
  wire _01720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15932" *)
  wire _01721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15941" *)
  wire _01722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15950" *)
  wire _01723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15960" *)
  wire _01724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15969" *)
  wire _01725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15978" *)
  wire _01726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15988" *)
  wire _01727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15997" *)
  wire _01728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16006" *)
  wire _01729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16016" *)
  wire _01730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16025" *)
  wire _01731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16034" *)
  wire _01732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16044" *)
  wire _01733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16053" *)
  wire _01734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16062" *)
  wire _01735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16072" *)
  wire _01736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16081" *)
  wire _01737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16090" *)
  wire _01738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16100" *)
  wire _01739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16109" *)
  wire _01740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16118" *)
  wire _01741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16128" *)
  wire _01742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16304" *)
  wire _01743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *)
  wire _01744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *)
  wire _01745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16312" *)
  wire _01746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *)
  wire _01747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *)
  wire _01748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16320" *)
  wire _01749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *)
  wire _01750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *)
  wire _01751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16328" *)
  wire _01752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *)
  wire _01753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *)
  wire _01754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16336" *)
  wire _01755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *)
  wire _01756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *)
  wire _01757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16344" *)
  wire _01758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *)
  wire _01759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *)
  wire _01760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16352" *)
  wire _01761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *)
  wire _01762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *)
  wire _01763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16360" *)
  wire _01764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *)
  wire _01765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *)
  wire _01766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16368" *)
  wire _01767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *)
  wire _01768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *)
  wire _01769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16376" *)
  wire _01770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *)
  wire _01771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *)
  wire _01772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16384" *)
  wire _01773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *)
  wire _01774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *)
  wire _01775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16393" *)
  wire _01776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *)
  wire _01777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *)
  wire _01778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16401" *)
  wire _01779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *)
  wire _01780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *)
  wire _01781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16409" *)
  wire _01782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *)
  wire _01783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *)
  wire _01784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16417" *)
  wire _01785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *)
  wire _01786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *)
  wire _01787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16425" *)
  wire _01788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *)
  wire _01789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *)
  wire _01790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16448" *)
  wire _01791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16449" *)
  wire _01792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16494" *)
  wire _01793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16503" *)
  wire _01794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16522" *)
  wire _01795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *)
  wire _01796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *)
  wire _01797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *)
  wire _01798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *)
  wire _01799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *)
  wire _01800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *)
  wire _01801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *)
  wire _01802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *)
  wire _01803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *)
  wire _01804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *)
  wire _01805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *)
  wire _01806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *)
  wire _01807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *)
  wire _01808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16717" *)
  wire _01809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16718" *)
  wire _01810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16718" *)
  wire _01811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16728" *)
  wire _01812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16736" *)
  wire _01813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16737" *)
  wire _01814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16737" *)
  wire _01815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16759" *)
  wire _01816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16760" *)
  wire _01817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16760" *)
  wire _01818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16770" *)
  wire _01819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16771" *)
  wire _01820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16771" *)
  wire _01821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16781" *)
  wire _01822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16781" *)
  wire _01823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16782" *)
  wire _01824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16792" *)
  wire _01825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16800" *)
  wire _01826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16801" *)
  wire _01827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16801" *)
  wire _01828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16831" *)
  wire _01829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16832" *)
  wire _01830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16832" *)
  wire _01831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16842" *)
  wire _01832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16843" *)
  wire _01833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16843" *)
  wire _01834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16853" *)
  wire _01835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16854" *)
  wire _01836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16854" *)
  wire _01837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16876" *)
  wire _01838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16877" *)
  wire _01839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16877" *)
  wire _01840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16887" *)
  wire _01841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16888" *)
  wire _01842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16888" *)
  wire _01843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16898" *)
  wire _01844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16899" *)
  wire _01845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16899" *)
  wire _01846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16909" *)
  wire _01847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16910" *)
  wire _01848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16910" *)
  wire _01849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16920" *)
  wire _01850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16921" *)
  wire _01851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16921" *)
  wire _01852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16931" *)
  wire _01853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16932" *)
  wire _01854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16932" *)
  wire _01855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16942" *)
  wire _01856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16950" *)
  wire _01857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16951" *)
  wire _01858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16951" *)
  wire _01859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16961" *)
  wire _01860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16969" *)
  wire _01861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16978" *)
  wire _01862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16978" *)
  wire _01863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17000" *)
  wire _01864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17009" *)
  wire _01865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17017" *)
  wire _01866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17026" *)
  wire _01867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17026" *)
  wire _01868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17036" *)
  wire _01869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17058" *)
  wire _01870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17068" *)
  wire _01871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17091" *)
  wire _01872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17100" *)
  wire _01873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17122" *)
  wire _01874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17132" *)
  wire _01875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17141" *)
  wire _01876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17150" *)
  wire _01877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17160" *)
  wire _01878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *)
  wire _01879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *)
  wire _01880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *)
  wire _01881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *)
  wire _01882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17220" *)
  wire _01883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17230" *)
  wire _01884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17239" *)
  wire _01885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17248" *)
  wire _01886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17257" *)
  wire _01887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *)
  wire _01888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *)
  wire _01889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *)
  wire _01890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *)
  wire _01891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17276" *)
  wire _01892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17286" *)
  wire _01893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17295" *)
  wire _01894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17304" *)
  wire _01895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17314" *)
  wire _01896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *)
  wire _01897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *)
  wire _01898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *)
  wire _01899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *)
  wire _01900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17344" *)
  wire _01901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17367" *)
  wire _01902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17376" *)
  wire _01903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17386" *)
  wire _01904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *)
  wire _01905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *)
  wire _01906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *)
  wire _01907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *)
  wire _01908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17406" *)
  wire _01909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17415" *)
  wire _01910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17424" *)
  wire _01911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17434" *)
  wire _01912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *)
  wire _01913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *)
  wire _01914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *)
  wire _01915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *)
  wire _01916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17462" *)
  wire _01917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17472" *)
  wire _01918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17482" *)
  wire _01919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17491" *)
  wire _01920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17500" *)
  wire _01921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17522" *)
  wire _01922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17532" *)
  wire _01923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17541" *)
  wire _01924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17550" *)
  wire _01925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17560" *)
  wire _01926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *)
  wire _01927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *)
  wire _01928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *)
  wire _01929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *)
  wire _01930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17580" *)
  wire _01931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17589" *)
  wire _01932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17598" *)
  wire _01933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17608" *)
  wire _01934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *)
  wire _01935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *)
  wire _01936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *)
  wire _01937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *)
  wire _01938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17628" *)
  wire _01939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17637" *)
  wire _01940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17646" *)
  wire _01941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17656" *)
  wire _01942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *)
  wire _01943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *)
  wire _01944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *)
  wire _01945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *)
  wire _01946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17686" *)
  wire _01947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17695" *)
  wire _01948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17704" *)
  wire _01949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17714" *)
  wire _01950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *)
  wire _01951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *)
  wire _01952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *)
  wire _01953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *)
  wire _01954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17734" *)
  wire _01955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17743" *)
  wire _01956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17764" *)
  wire _01957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17773" *)
  wire _01958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17774" *)
  wire _01959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17774" *)
  wire _01960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17782" *)
  wire _01961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *)
  wire _01962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *)
  wire _01963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *)
  wire _01964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *)
  wire _01965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17801" *)
  wire _01966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17810" *)
  wire _01967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17819" *)
  wire _01968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17829" *)
  wire _01969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17838" *)
  wire _01970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *)
  wire _01971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *)
  wire _01972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *)
  wire _01973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *)
  wire _01974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17857" *)
  wire _01975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17866" *)
  wire _01976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17875" *)
  wire _01977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17885" *)
  wire _01978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17894" *)
  wire _01979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *)
  wire _01980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *)
  wire _01981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *)
  wire _01982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *)
  wire _01983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17913" *)
  wire _01984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17922" *)
  wire _01985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17954" *)
  wire _01986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18029" *)
  wire _01987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18030" *)
  wire _01988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18041" *)
  wire _01989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18136" *)
  wire _01990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18149" *)
  wire _01991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18157" *)
  wire _01992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18166" *)
  wire _01993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18166" *)
  wire _01994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18174" *)
  wire _01995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *)
  wire _01996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *)
  wire _01997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18186" *)
  wire _01998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18199" *)
  wire _01999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18283" *)
  wire _02000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18296" *)
  wire _02001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18305" *)
  wire _02002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18340" *)
  wire _02003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18349" *)
  wire _02004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18350" *)
  wire _02005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18361" *)
  wire _02006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18369" *)
  wire _02007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18369" *)
  wire _02008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18381" *)
  wire _02009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18414" *)
  wire _02010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18425" *)
  wire _02011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18438" *)
  wire _02012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18473" *)
  wire _02013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18474" *)
  wire _02014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18485" *)
  wire _02015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18486" *)
  wire _02016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18486" *)
  wire _02017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18495" *)
  wire _02018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18495" *)
  wire _02019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18503" *)
  wire _02020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18512" *)
  wire _02021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18513" *)
  wire _02022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18524" *)
  wire _02023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18532" *)
  wire _02024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18544" *)
  wire _02025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18557" *)
  wire _02026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18567" *)
  wire _02027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18567" *)
  wire _02028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18575" *)
  wire _02029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18575" *)
  wire _02030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18583" *)
  wire _02031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18592" *)
  wire _02032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18593" *)
  wire _02033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18604" *)
  wire _02034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18615" *)
  wire _02035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18628" *)
  wire _02036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18639" *)
  wire _02037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18652" *)
  wire _02038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18663" *)
  wire _02039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18676" *)
  wire _02040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18687" *)
  wire _02041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18703" *)
  wire _02042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18810" *)
  wire _02043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18883" *)
  wire _02044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18883" *)
  wire _02045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18891" *)
  wire _02046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18900" *)
  wire _02047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18900" *)
  wire _02048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18908" *)
  wire _02049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18938" *)
  wire _02050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18939" *)
  wire _02051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18959" *)
  wire _02052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18967" *)
  wire _02053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18987" *)
  wire _02054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18989" *)
  wire _02055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18989" *)
  wire _02056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *)
  wire _02057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *)
  wire _02058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *)
  wire _02059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18998" *)
  wire _02060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18998" *)
  wire _02061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18999" *)
  wire _02062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19000" *)
  wire _02063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19000" *)
  wire _02064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19000" *)
  wire _02065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19008" *)
  wire _02066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19008" *)
  wire _02067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19009" *)
  wire _02068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19009" *)
  wire _02069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19018" *)
  wire _02070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19027" *)
  wire _02071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19027" *)
  wire _02072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19028" *)
  wire _02073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19037" *)
  wire _02074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19037" *)
  wire _02075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19037" *)
  wire _02076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *)
  wire _02077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *)
  wire _02078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *)
  wire _02079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19039" *)
  wire _02080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *)
  wire _02081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *)
  wire _02082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *)
  wire _02083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19041" *)
  wire _02084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19049" *)
  wire _02085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19049" *)
  wire _02086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19050" *)
  wire _02087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19050" *)
  wire _02088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19061" *)
  wire _02089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19061" *)
  wire _02090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19064" *)
  wire _02091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19064" *)
  wire _02092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19072" *)
  wire _02093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19072" *)
  wire _02094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19072" *)
  wire _02095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *)
  wire _02096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *)
  wire _02097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *)
  wire _02098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19074" *)
  wire _02099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19075" *)
  wire _02100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19075" *)
  wire _02101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19075" *)
  wire _02102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19076" *)
  wire _02103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19084" *)
  wire _02104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19084" *)
  wire _02105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19085" *)
  wire _02106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19085" *)
  wire _02107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19094" *)
  wire _02108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19103" *)
  wire _02109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19103" *)
  wire _02110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19104" *)
  wire _02111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19113" *)
  wire _02112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19113" *)
  wire _02113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19113" *)
  wire _02114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *)
  wire _02115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *)
  wire _02116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *)
  wire _02117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *)
  wire _02118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19115" *)
  wire _02119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19116" *)
  wire _02120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19116" *)
  wire _02121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19117" *)
  wire _02122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19117" *)
  wire _02123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19125" *)
  wire _02124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19125" *)
  wire _02125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19126" *)
  wire _02126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19134" *)
  wire _02127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19134" *)
  wire _02128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19134" *)
  wire _02129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *)
  wire _02130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *)
  wire _02131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *)
  wire _02132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19136" *)
  wire _02133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19137" *)
  wire _02134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19137" *)
  wire _02135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19137" *)
  wire _02136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19138" *)
  wire _02137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19146" *)
  wire _02138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19146" *)
  wire _02139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19147" *)
  wire _02140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19147" *)
  wire _02141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19156" *)
  wire _02142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19166" *)
  wire _02143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19166" *)
  wire _02144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19175" *)
  wire _02145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19175" *)
  wire _02146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19175" *)
  wire _02147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *)
  wire _02148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *)
  wire _02149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *)
  wire _02150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *)
  wire _02151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19177" *)
  wire _02152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19178" *)
  wire _02153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19178" *)
  wire _02154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19179" *)
  wire _02155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19179" *)
  wire _02156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19187" *)
  wire _02157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19187" *)
  wire _02158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19188" *)
  wire _02159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19188" *)
  wire _02160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19197" *)
  wire _02161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19206" *)
  wire _02162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19206" *)
  wire _02163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19206" *)
  wire _02164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *)
  wire _02165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *)
  wire _02166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *)
  wire _02167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *)
  wire _02168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19208" *)
  wire _02169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19209" *)
  wire _02170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19209" *)
  wire _02171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19210" *)
  wire _02172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19210" *)
  wire _02173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19218" *)
  wire _02174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19218" *)
  wire _02175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19219" *)
  wire _02176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19219" *)
  wire _02177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19228" *)
  wire _02178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19237" *)
  wire _02179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19237" *)
  wire _02180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19237" *)
  wire _02181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *)
  wire _02182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *)
  wire _02183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *)
  wire _02184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *)
  wire _02185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19239" *)
  wire _02186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19240" *)
  wire _02187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19240" *)
  wire _02188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19241" *)
  wire _02189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19241" *)
  wire _02190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19249" *)
  wire _02191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19249" *)
  wire _02192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19250" *)
  wire _02193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19250" *)
  wire _02194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19258" *)
  wire _02195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19260" *)
  wire _02196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19260" *)
  wire _02197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19268" *)
  wire _02198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19268" *)
  wire _02199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19268" *)
  wire _02200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *)
  wire _02201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *)
  wire _02202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *)
  wire _02203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19270" *)
  wire _02204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19271" *)
  wire _02205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19271" *)
  wire _02206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19271" *)
  wire _02207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19272" *)
  wire _02208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19280" *)
  wire _02209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19280" *)
  wire _02210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19281" *)
  wire _02211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19281" *)
  wire _02212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19290" *)
  wire _02213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19299" *)
  wire _02214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19308" *)
  wire _02215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19308" *)
  wire _02216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19308" *)
  wire _02217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *)
  wire _02218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *)
  wire _02219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *)
  wire _02220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *)
  wire _02221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19310" *)
  wire _02222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19311" *)
  wire _02223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19311" *)
  wire _02224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19312" *)
  wire _02225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19312" *)
  wire _02226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19320" *)
  wire _02227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19320" *)
  wire _02228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19321" *)
  wire _02229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19321" *)
  wire _02230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19329" *)
  wire _02231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19330" *)
  wire _02232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19339" *)
  wire _02233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19339" *)
  wire _02234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19339" *)
  wire _02235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *)
  wire _02236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *)
  wire _02237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *)
  wire _02238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *)
  wire _02239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19341" *)
  wire _02240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19342" *)
  wire _02241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19342" *)
  wire _02242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19343" *)
  wire _02243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19343" *)
  wire _02244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19351" *)
  wire _02245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19351" *)
  wire _02246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19352" *)
  wire _02247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19352" *)
  wire _02248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19361" *)
  wire _02249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19370" *)
  wire _02250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19370" *)
  wire _02251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19370" *)
  wire _02252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *)
  wire _02253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *)
  wire _02254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *)
  wire _02255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *)
  wire _02256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19372" *)
  wire _02257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19373" *)
  wire _02258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19373" *)
  wire _02259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19374" *)
  wire _02260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19374" *)
  wire _02261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19382" *)
  wire _02262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19382" *)
  wire _02263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19383" *)
  wire _02264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19383" *)
  wire _02265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19403" *)
  wire _02266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19403" *)
  wire _02267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19403" *)
  wire _02268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *)
  wire _02269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *)
  wire _02270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *)
  wire _02271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *)
  wire _02272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19405" *)
  wire _02273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19406" *)
  wire _02274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19406" *)
  wire _02275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19407" *)
  wire _02276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19407" *)
  wire _02277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19415" *)
  wire _02278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19415" *)
  wire _02279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19416" *)
  wire _02280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19416" *)
  wire _02281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19424" *)
  wire _02282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19432" *)
  wire _02283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19440" *)
  wire _02284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19440" *)
  wire _02285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19440" *)
  wire _02286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *)
  wire _02287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *)
  wire _02288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *)
  wire _02289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *)
  wire _02290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19442" *)
  wire _02291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19443" *)
  wire _02292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19443" *)
  wire _02293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19444" *)
  wire _02294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19444" *)
  wire _02295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19452" *)
  wire _02296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19452" *)
  wire _02297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19453" *)
  wire _02298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19461" *)
  wire _02299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19461" *)
  wire _02300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19490" *)
  wire _02301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19490" *)
  wire _02302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19490" *)
  wire _02303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *)
  wire _02304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *)
  wire _02305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *)
  wire _02306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *)
  wire _02307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19492" *)
  wire _02308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19493" *)
  wire _02309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19493" *)
  wire _02310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19494" *)
  wire _02311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19494" *)
  wire _02312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19502" *)
  wire _02313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19502" *)
  wire _02314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19503" *)
  wire _02315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19511" *)
  wire _02316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19511" *)
  wire _02317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19511" *)
  wire _02318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *)
  wire _02319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *)
  wire _02320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *)
  wire _02321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *)
  wire _02322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19513" *)
  wire _02323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19514" *)
  wire _02324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19514" *)
  wire _02325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19515" *)
  wire _02326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19515" *)
  wire _02327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19523" *)
  wire _02328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19523" *)
  wire _02329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19524" *)
  wire _02330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19524" *)
  wire _02331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19532" *)
  wire _02332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19540" *)
  wire _02333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19568" *)
  wire _02334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19578" *)
  wire _02335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19578" *)
  wire _02336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19586" *)
  wire _02337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19587" *)
  wire _02338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19607" *)
  wire _02339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19607" *)
  wire _02340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *)
  wire _02341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *)
  wire _02342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *)
  wire _02343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *)
  wire _02344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19609" *)
  wire _02345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19609" *)
  wire _02346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19663" *)
  wire _02347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19663" *)
  wire _02348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19699" *)
  wire _02349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19700" *)
  wire _02350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19805" *)
  wire _02351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19813" *)
  wire _02352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19821" *)
  wire _02353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19829" *)
  wire _02354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19837" *)
  wire _02355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19845" *)
  wire _02356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19853" *)
  wire _02357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19861" *)
  wire _02358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19869" *)
  wire _02359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19877" *)
  wire _02360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19885" *)
  wire _02361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19893" *)
  wire _02362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19901" *)
  wire _02363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19909" *)
  wire _02364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19917" *)
  wire _02365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19925" *)
  wire _02366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19933" *)
  wire _02367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19941" *)
  wire _02368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19949" *)
  wire _02369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19957" *)
  wire _02370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19965" *)
  wire _02371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19973" *)
  wire _02372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19981" *)
  wire _02373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19989" *)
  wire _02374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19997" *)
  wire _02375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20005" *)
  wire _02376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20013" *)
  wire _02377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20021" *)
  wire _02378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20029" *)
  wire _02379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20037" *)
  wire _02380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20045" *)
  wire _02381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20053" *)
  wire _02382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20061" *)
  wire _02383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20069" *)
  wire _02384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20078" *)
  wire _02385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20078" *)
  wire _02386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20078" *)
  wire _02387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *)
  wire _02388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *)
  wire _02389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20088" *)
  wire _02390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20097" *)
  wire _02391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20097" *)
  wire _02392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20097" *)
  wire _02393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20098" *)
  wire _02394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20098" *)
  wire _02395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20107" *)
  wire _02396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20116" *)
  wire _02397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20116" *)
  wire _02398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20116" *)
  wire _02399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20117" *)
  wire _02400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20117" *)
  wire _02401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20126" *)
  wire _02402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20135" *)
  wire _02403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20135" *)
  wire _02404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20135" *)
  wire _02405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20136" *)
  wire _02406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20136" *)
  wire _02407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20145" *)
  wire _02408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20154" *)
  wire _02409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20154" *)
  wire _02410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20154" *)
  wire _02411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20155" *)
  wire _02412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20155" *)
  wire _02413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20164" *)
  wire _02414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20173" *)
  wire _02415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20173" *)
  wire _02416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20173" *)
  wire _02417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20174" *)
  wire _02418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20174" *)
  wire _02419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20183" *)
  wire _02420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20192" *)
  wire _02421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20192" *)
  wire _02422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20192" *)
  wire _02423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20193" *)
  wire _02424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20193" *)
  wire _02425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20202" *)
  wire _02426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20211" *)
  wire _02427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20211" *)
  wire _02428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20211" *)
  wire _02429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20212" *)
  wire _02430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20212" *)
  wire _02431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20221" *)
  wire _02432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20230" *)
  wire _02433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20230" *)
  wire _02434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20230" *)
  wire _02435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20231" *)
  wire _02436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20231" *)
  wire _02437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20240" *)
  wire _02438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20249" *)
  wire _02439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20249" *)
  wire _02440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20249" *)
  wire _02441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20250" *)
  wire _02442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20250" *)
  wire _02443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20259" *)
  wire _02444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20268" *)
  wire _02445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20268" *)
  wire _02446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20268" *)
  wire _02447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20269" *)
  wire _02448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20269" *)
  wire _02449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20278" *)
  wire _02450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20287" *)
  wire _02451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20287" *)
  wire _02452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20287" *)
  wire _02453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20288" *)
  wire _02454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20288" *)
  wire _02455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20297" *)
  wire _02456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20306" *)
  wire _02457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20306" *)
  wire _02458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20306" *)
  wire _02459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20307" *)
  wire _02460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20307" *)
  wire _02461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20316" *)
  wire _02462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20325" *)
  wire _02463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20325" *)
  wire _02464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20325" *)
  wire _02465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20326" *)
  wire _02466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20326" *)
  wire _02467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20335" *)
  wire _02468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20344" *)
  wire _02469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20344" *)
  wire _02470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20344" *)
  wire _02471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20345" *)
  wire _02472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20345" *)
  wire _02473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20354" *)
  wire _02474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20363" *)
  wire _02475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20363" *)
  wire _02476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20363" *)
  wire _02477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20364" *)
  wire _02478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20364" *)
  wire _02479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20375" *)
  wire _02480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20375" *)
  wire _02481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20387" *)
  wire _02482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20387" *)
  wire _02483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20399" *)
  wire _02484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20399" *)
  wire _02485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20411" *)
  wire _02486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20411" *)
  wire _02487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20423" *)
  wire _02488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20423" *)
  wire _02489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20435" *)
  wire _02490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20435" *)
  wire _02491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20447" *)
  wire _02492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20447" *)
  wire _02493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20459" *)
  wire _02494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20459" *)
  wire _02495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20471" *)
  wire _02496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20471" *)
  wire _02497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20483" *)
  wire _02498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20483" *)
  wire _02499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20495" *)
  wire _02500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20495" *)
  wire _02501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20506" *)
  wire _02502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20507" *)
  wire _02503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20518" *)
  wire _02504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20519" *)
  wire _02505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20530" *)
  wire _02506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20531" *)
  wire _02507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20542" *)
  wire _02508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20543" *)
  wire _02509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20554" *)
  wire _02510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20555" *)
  wire _02511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20581" *)
  wire _02512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20583" *)
  wire _02513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20585" *)
  wire _02514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20587" *)
  wire _02515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20589" *)
  wire _02516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20591" *)
  wire _02517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20593" *)
  wire _02518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20595" *)
  wire _02519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20597" *)
  wire _02520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20599" *)
  wire _02521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20601" *)
  wire _02522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20603" *)
  wire _02523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20605" *)
  wire _02524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20607" *)
  wire _02525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20609" *)
  wire _02526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20616" *)
  wire _02527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20625" *)
  wire _02528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20635" *)
  wire _02529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20646" *)
  wire _02530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20656" *)
  wire _02531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20666" *)
  wire _02532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20676" *)
  wire _02533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20701" *)
  wire _02534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20726" *)
  wire _02535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20726" *)
  wire _02536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20737" *)
  wire _02537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20762" *)
  wire _02538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20787" *)
  wire _02539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20787" *)
  wire _02540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20798" *)
  wire _02541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20809" *)
  wire _02542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20819" *)
  wire _02543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20819" *)
  wire _02544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20820" *)
  wire _02545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20820" *)
  wire _02546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *)
  wire _02547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *)
  wire _02548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *)
  wire _02549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *)
  wire _02550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *)
  wire _02551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *)
  wire _02552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *)
  wire _02553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *)
  wire _02554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *)
  wire _02555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *)
  wire _02556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *)
  wire _02557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *)
  wire _02558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20904" *)
  wire _02559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20914" *)
  wire _02560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20914" *)
  wire _02561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *)
  wire _02562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *)
  wire _02563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *)
  wire _02564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *)
  wire _02565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *)
  wire _02566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *)
  wire _02567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *)
  wire _02568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *)
  wire _02569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *)
  wire _02570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20979" *)
  wire _02571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20989" *)
  wire _02572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20989" *)
  wire _02573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *)
  wire _02574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *)
  wire _02575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21007" *)
  wire _02576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *)
  wire _02577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *)
  wire _02578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *)
  wire _02579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *)
  wire _02580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *)
  wire _02581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21045" *)
  wire _02582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21055" *)
  wire _02583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21065" *)
  wire _02584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21065" *)
  wire _02585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21075" *)
  wire _02586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *)
  wire _02587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *)
  wire _02588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21094" *)
  wire _02589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *)
  wire _02590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *)
  wire _02591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *)
  wire _02592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *)
  wire _02593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21122" *)
  wire _02594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21152" *)
  wire _02595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *)
  wire _02596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *)
  wire _02597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21180" *)
  wire _02598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21180" *)
  wire _02599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *)
  wire _02600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *)
  wire _02601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21206" *)
  wire _02602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21207" *)
  wire _02603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21226" *)
  wire _02604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21234" *)
  wire _02605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21234" *)
  wire _02606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21243" *)
  wire _02607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21252" *)
  wire _02608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *)
  wire _02609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *)
  wire _02610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *)
  wire _02611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *)
  wire _02612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *)
  wire _02613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *)
  wire _02614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *)
  wire _02615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *)
  wire _02616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *)
  wire _02617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *)
  wire _02618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *)
  wire _02619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *)
  wire _02620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *)
  wire _02621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *)
  wire _02622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *)
  wire _02623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *)
  wire _02624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21429" *)
  wire _02625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21431" *)
  wire _02626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21433" *)
  wire _02627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21435" *)
  wire _02628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21437" *)
  wire _02629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21439" *)
  wire _02630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21441" *)
  wire _02631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21443" *)
  wire _02632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21445" *)
  wire _02633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21447" *)
  wire _02634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21449" *)
  wire _02635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21451" *)
  wire _02636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21453" *)
  wire _02637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21455" *)
  wire _02638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21457" *)
  wire _02639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21459" *)
  wire _02640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21547" *)
  wire _02641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21574" *)
  wire _02642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21600" *)
  wire _02643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21627" *)
  wire _02644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21654" *)
  wire _02645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21681" *)
  wire _02646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21708" *)
  wire _02647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21735" *)
  wire _02648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21762" *)
  wire _02649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21789" *)
  wire _02650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21816" *)
  wire _02651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21843" *)
  wire _02652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21870" *)
  wire _02653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21920" *)
  wire _02654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21935" *)
  wire _02655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21969" *)
  wire _02656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21969" *)
  wire _02657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *)
  wire _02658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *)
  wire _02659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *)
  wire _02660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22096" *)
  wire _02661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22096" *)
  wire _02662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22125" *)
  wire _02663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22125" *)
  wire _02664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22147" *)
  wire _02665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22147" *)
  wire _02666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22224" *)
  wire _02667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22224" *)
  wire _02668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22301" *)
  wire _02669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22301" *)
  wire _02670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22538" *)
  wire _02671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22541" *)
  wire _02672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22556" *)
  wire _02673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22573" *)
  wire _02674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22575" *)
  wire _02675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22589" *)
  wire _02676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22610" *)
  wire _02677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22629" *)
  wire _02678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22631" *)
  wire _02679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22647" *)
  wire _02680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22648" *)
  wire _02681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22663" *)
  wire _02682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22664" *)
  wire _02683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22697" *)
  wire _02684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22699" *)
  wire _02685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22715" *)
  wire _02686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22717" *)
  wire _02687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22733" *)
  wire _02688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22752" *)
  wire _02689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22757" *)
  wire _02690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22773" *)
  wire _02691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22792" *)
  wire _02692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22797" *)
  wire _02693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22817" *)
  wire _02694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22822" *)
  wire _02695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22887" *)
  wire _02696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22901" *)
  wire _02697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22911" *)
  wire _02698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *)
  wire _02699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22937" *)
  wire _02700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22953" *)
  wire _02701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22958" *)
  wire _02702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22960" *)
  wire _02703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22962" *)
  wire _02704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22971" *)
  wire _02705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22986" *)
  wire _02706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23000" *)
  wire _02707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23022" *)
  wire _02708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23032" *)
  wire _02709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23047" *)
  wire _02710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23061" *)
  wire _02711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23076" *)
  wire _02712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23090" *)
  wire _02713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23094" *)
  wire _02714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *)
  wire _02715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *)
  wire _02716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23140" *)
  wire _02717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23160" *)
  wire _02718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23170" *)
  wire _02719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23180" *)
  wire _02720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23190" *)
  wire _02721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23200" *)
  wire _02722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23364" *)
  wire _02723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23380" *)
  wire _02724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23381" *)
  wire _02725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23393" *)
  wire _02726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *)
  wire _02727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23412" *)
  wire _02728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *)
  wire _02729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23426" *)
  wire _02730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *)
  wire _02731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23435" *)
  wire _02732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *)
  wire _02733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23453" *)
  wire _02734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *)
  wire _02735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23465" *)
  wire _02736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *)
  wire _02737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23481" *)
  wire _02738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *)
  wire _02739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23499" *)
  wire _02740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *)
  wire _02741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23509" *)
  wire _02742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23510" *)
  wire _02743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *)
  wire _02744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23522" *)
  wire _02745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *)
  wire _02746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23530" *)
  wire _02747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23543" *)
  wire _02748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *)
  wire _02749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23550" *)
  wire _02750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23551" *)
  wire _02751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *)
  wire _02752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23556" *)
  wire _02753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23557" *)
  wire _02754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23557" *)
  wire _02755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23562" *)
  wire _02756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23563" *)
  wire _02757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23563" *)
  wire _02758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23571" *)
  wire _02759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23572" *)
  wire _02760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *)
  wire _02761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23580" *)
  wire _02762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23581" *)
  wire _02763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *)
  wire _02764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23589" *)
  wire _02765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *)
  wire _02766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23620" *)
  wire _02767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23625" *)
  wire _02768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23644" *)
  wire _02769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23667" *)
  wire _02770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23690" *)
  wire _02771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23713" *)
  wire _02772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23736" *)
  wire _02773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23738" *)
  wire _02774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23738" *)
  wire _02775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *)
  wire _02776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *)
  wire _02777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *)
  wire _02778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23759" *)
  wire _02779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23782" *)
  wire _02780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23805" *)
  wire _02781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23828" *)
  wire _02782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23851" *)
  wire _02783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23874" *)
  wire _02784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23897" *)
  wire _02785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23920" *)
  wire _02786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23943" *)
  wire _02787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23966" *)
  wire _02788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23989" *)
  wire _02789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24031" *)
  wire _02790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24033" *)
  wire _02791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *)
  wire _02792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24056" *)
  wire _02793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24058" *)
  wire _02794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24063" *)
  wire _02795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24099" *)
  wire _02796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24110" *)
  wire _02797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24119" *)
  wire _02798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24132" *)
  wire _02799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24229" *)
  wire _02800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *)
  wire _02863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _02926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _02989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _02999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _03000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _03001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _03002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _03003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _03004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *)
  wire _03005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _03021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _03037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _03053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _03069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *)
  wire [14:0] _03097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _03125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _03153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24297" *)
  wire [14:0] _03154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24297" *)
  wire [14:0] _03155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24297" *)
  wire [14:0] _03156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *)
  wire [14:0] _03157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *)
  wire [14:0] _03158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *)
  wire [14:0] _03159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *)
  wire [14:0] _03160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *)
  wire [14:0] _03161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *)
  wire [14:0] _03162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *)
  wire [14:0] _03163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *)
  wire [14:0] _03164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *)
  wire [14:0] _03165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *)
  wire [14:0] _03166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *)
  wire [14:0] _03167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *)
  wire [14:0] _03168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *)
  wire [14:0] _03169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *)
  wire [14:0] _03170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *)
  wire [14:0] _03171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *)
  wire [14:0] _03184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _03197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _03210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _03223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _03236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _03249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *)
  wire [14:0] _03262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24334" *)
  wire [15:0] _03263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24335" *)
  wire [15:0] _03264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24336" *)
  wire [15:0] _03265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *)
  wire [3:0] _03281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _03297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _03313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *)
  wire [3:0] _03329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *)
  wire [3:0] _03345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _03361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _03377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _03393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _03409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _03425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *)
  wire [4:0] _03441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _03457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *)
  wire [4:0] _03473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *)
  wire [6:0] _03489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03520_;
  wire [1:0] _03521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24408" *)
  wire [8:0] _03522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24409" *)
  wire [8:0] _03523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24410" *)
  wire [8:0] _03524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24411" *)
  wire [8:0] _03525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *)
  wire [8:0] _03540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _03555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _03570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _03585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _03600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8773" *)
  wire _03601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8773" *)
  wire _03602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8777" *)
  wire _03603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8779" *)
  wire _03604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8779" *)
  wire _03605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8781" *)
  wire _03606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8781" *)
  wire _03607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8783" *)
  wire _03608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8783" *)
  wire _03609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8785" *)
  wire _03610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8785" *)
  wire _03611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8786" *)
  wire _03612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8788" *)
  wire _03613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8788" *)
  wire _03614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8790" *)
  wire _03615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8790" *)
  wire _03616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8792" *)
  wire _03617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8792" *)
  wire _03618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8794" *)
  wire _03619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8794" *)
  wire _03620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8796" *)
  wire _03621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8796" *)
  wire _03622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8800" *)
  wire _03623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8802" *)
  wire _03624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8802" *)
  wire _03625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8805" *)
  wire _03626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8805" *)
  wire _03627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8806" *)
  wire _03628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8807" *)
  wire _03629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8809" *)
  wire _03630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8809" *)
  wire _03631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8822" *)
  wire _03632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8871" *)
  wire _03633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8872" *)
  wire _03634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8872" *)
  wire _03635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8882" *)
  wire _03636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8883" *)
  wire _03637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8883" *)
  wire _03638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8893" *)
  wire _03639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8894" *)
  wire _03640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8895" *)
  wire _03641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8899" *)
  wire _03642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8900" *)
  wire _03643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8901" *)
  wire _03644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8921" *)
  wire _03645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8922" *)
  wire _03646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8939" *)
  wire _03647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8940" *)
  wire _03648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8957" *)
  wire _03649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8958" *)
  wire _03650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8968" *)
  wire _03651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8969" *)
  wire _03652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8976" *)
  wire _03653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8977" *)
  wire _03654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8977" *)
  wire _03655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8984" *)
  wire _03656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8985" *)
  wire _03657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8992" *)
  wire _03658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8993" *)
  wire _03659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9001" *)
  wire _03660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9002" *)
  wire _03661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9014" *)
  wire _03662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9015" *)
  wire _03663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9016" *)
  wire _03664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9032" *)
  wire _03665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9032" *)
  wire _03666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9038" *)
  wire _03667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9038" *)
  wire _03668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9048" *)
  wire _03669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9049" *)
  wire _03670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9051" *)
  wire _03671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9059" *)
  wire _03672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9060" *)
  wire _03673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9091" *)
  wire _03674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9103" *)
  wire _03675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9107" *)
  wire _03676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9121" *)
  wire _03677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9123" *)
  wire _03678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9125" *)
  wire _03679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9129" *)
  wire _03680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9130" *)
  wire _03681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9152" *)
  wire _03682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9154" *)
  wire _03683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9156" *)
  wire _03684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9167" *)
  wire _03685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9172" *)
  wire _03686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9174" *)
  wire _03687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9184" *)
  wire _03688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9186" *)
  wire _03689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9188" *)
  wire _03690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9192" *)
  wire _03691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9202" *)
  wire _03692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *)
  wire _03693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *)
  wire _03694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9209" *)
  wire _03695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9213" *)
  wire _03696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9215" *)
  wire _03697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9217" *)
  wire _03698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9239" *)
  wire _03699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9241" *)
  wire _03700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9243" *)
  wire _03701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9247" *)
  wire _03702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9248" *)
  wire _03703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9263" *)
  wire _03704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9266" *)
  wire _03705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9277" *)
  wire _03706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9279" *)
  wire _03707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9281" *)
  wire _03708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *)
  wire _03709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9292" *)
  wire _03710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9293" *)
  wire _03711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *)
  wire _03712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9295" *)
  wire _03713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9300" *)
  wire _03714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9302" *)
  wire _03715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9304" *)
  wire _03716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9306" *)
  wire _03717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9324" *)
  wire _03718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9329" *)
  wire _03719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9331" *)
  wire _03720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9333" *)
  wire _03721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9346" *)
  wire _03722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9348" *)
  wire _03723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9350" *)
  wire _03724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9354" *)
  wire _03725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9355" *)
  wire _03726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9355" *)
  wire _03727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9367" *)
  wire _03728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9373" *)
  wire _03729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9377" *)
  wire _03730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9379" *)
  wire _03731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9381" *)
  wire _03732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9395" *)
  wire _03733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9397" *)
  wire _03734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9399" *)
  wire _03735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9404" *)
  wire _03736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9404" *)
  wire _03737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9424" *)
  wire _03738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9426" *)
  wire _03739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9428" *)
  wire _03740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9444" *)
  wire _03741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9446" *)
  wire _03742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9448" *)
  wire _03743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9461" *)
  wire _03744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9463" *)
  wire _03745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9465" *)
  wire _03746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9482" *)
  wire _03747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *)
  wire _03748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9507" *)
  wire _03749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9512" *)
  wire _03750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9513" *)
  wire _03751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9513" *)
  wire _03752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9525" *)
  wire _03753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9526" *)
  wire _03754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9533" *)
  wire _03755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9533" *)
  wire _03756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9554" *)
  wire _03757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9554" *)
  wire _03758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9569" *)
  wire _03759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9569" *)
  wire _03760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9569" *)
  wire _03761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9575" *)
  wire _03762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9581" *)
  wire _03763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9582" *)
  wire _03764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9582" *)
  wire _03765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9595" *)
  wire _03766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9595" *)
  wire _03767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9603" *)
  wire _03768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9603" *)
  wire _03769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9603" *)
  wire _03770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9605" *)
  wire _03771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9614" *)
  wire _03772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9614" *)
  wire _03773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9627" *)
  wire _03774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9627" *)
  wire _03775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9640" *)
  wire _03776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9640" *)
  wire _03777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9650" *)
  wire _03778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9656" *)
  wire _03779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9657" *)
  wire _03780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9657" *)
  wire _03781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9664" *)
  wire _03782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9672" *)
  wire _03783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9672" *)
  wire _03784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9682" *)
  wire _03785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9688" *)
  wire _03786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9689" *)
  wire _03787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9689" *)
  wire _03788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9698" *)
  wire _03789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9704" *)
  wire _03790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9705" *)
  wire _03791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9705" *)
  wire _03792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9713" *)
  wire _03793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9716" *)
  wire _03794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9721" *)
  wire _03795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9722" *)
  wire _03796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9722" *)
  wire _03797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9735" *)
  wire _03798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9735" *)
  wire _03799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9749" *)
  wire _03800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9755" *)
  wire _03801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9755" *)
  wire _03802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9764" *)
  wire _03803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9769" *)
  wire _03804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9770" *)
  wire _03805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9770" *)
  wire _03806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9785" *)
  wire _03807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9787" *)
  wire _03808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9789" *)
  wire _03809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9792" *)
  wire _03810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *)
  wire _03811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *)
  wire _03812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *)
  wire _03813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *)
  wire _03814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9832" *)
  wire _03815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9832" *)
  wire _03816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9839" *)
  wire _03817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9840" *)
  wire _03818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9861" *)
  wire _03819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9869" *)
  wire _03820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9879" *)
  wire _03821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9884" *)
  wire _03822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9902" *)
  wire _03823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9918" *)
  wire _03824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9920" *)
  wire _03825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9922" *)
  wire _03826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9924" *)
  wire _03827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9926" *)
  wire _03828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9928" *)
  wire _03829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9930" *)
  wire _03830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9932" *)
  wire _03831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9934" *)
  wire _03832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9936" *)
  wire _03833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9938" *)
  wire _03834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9940" *)
  wire _03835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9942" *)
  wire _03836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9944" *)
  wire _03837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9946" *)
  wire _03838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9948" *)
  wire _03839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9968" *)
  wire _03840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9974" *)
  wire _03841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9980" *)
  wire _03842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9986" *)
  wire _03843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9992" *)
  wire _03844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9998" *)
  wire _03845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *)
  wire [6:0] _03846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10137" *)
  (* unused_bits = "3" *)
  wire [3:0] _03847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10149" *)
  (* unused_bits = "3" *)
  wire [3:0] _03848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10161" *)
  (* unused_bits = "3" *)
  wire [3:0] _03849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10173" *)
  (* unused_bits = "3" *)
  wire [3:0] _03850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10185" *)
  (* unused_bits = "3" *)
  wire [3:0] _03851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10197" *)
  (* unused_bits = "3" *)
  wire [3:0] _03852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10209" *)
  (* unused_bits = "3" *)
  wire [3:0] _03853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10221" *)
  (* unused_bits = "3" *)
  wire [3:0] _03854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10233" *)
  (* unused_bits = "3" *)
  wire [3:0] _03855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10245" *)
  (* unused_bits = "3" *)
  wire [3:0] _03856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10257" *)
  (* unused_bits = "3" *)
  wire [3:0] _03857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10269" *)
  (* unused_bits = "3" *)
  wire [3:0] _03858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10281" *)
  (* unused_bits = "3" *)
  wire [3:0] _03859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10293" *)
  (* unused_bits = "3" *)
  wire [3:0] _03860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10305" *)
  (* unused_bits = "3" *)
  wire [3:0] _03861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10317" *)
  (* unused_bits = "3" *)
  wire [3:0] _03862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _03863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6316" *)
  wire [17:0] _03864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10120" *)
  wire _03865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11529" *)
  wire _03866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11536" *)
  wire _03867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11543" *)
  wire _03868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11550" *)
  wire _03869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11557" *)
  wire _03870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11564" *)
  wire _03871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11571" *)
  wire _03872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11578" *)
  wire _03873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11585" *)
  wire _03874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11592" *)
  wire _03875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11599" *)
  wire _03876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11604" *)
  wire _03877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11606" *)
  wire _03878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11613" *)
  wire _03879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11620" *)
  wire _03880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11627" *)
  wire _03881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11634" *)
  wire _03882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11857" *)
  wire _03883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11859" *)
  wire _03884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11861" *)
  wire _03885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11863" *)
  wire _03886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11865" *)
  wire _03887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11867" *)
  wire _03888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11869" *)
  wire _03889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11871" *)
  wire _03890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11873" *)
  wire _03891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11875" *)
  wire _03892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11877" *)
  wire _03893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11879" *)
  wire _03894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11881" *)
  wire _03895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11883" *)
  wire _03896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11885" *)
  wire _03897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11887" *)
  wire _03898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11933" *)
  wire _03899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11981" *)
  wire _03900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12021" *)
  wire _03901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12069" *)
  wire _03902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12117" *)
  wire _03903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12157" *)
  wire _03904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12197" *)
  wire _03905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12245" *)
  wire _03906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12293" *)
  wire _03907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12333" *)
  wire _03908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12381" *)
  wire _03909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12429" *)
  wire _03910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12469" *)
  wire _03911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12509" *)
  wire _03912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12549" *)
  wire _03913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12589" *)
  wire _03914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12613" *)
  wire _03915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12641" *)
  wire _03916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12669" *)
  wire _03917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12697" *)
  wire _03918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12725" *)
  wire _03919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12753" *)
  wire _03920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12781" *)
  wire _03921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12809" *)
  wire _03922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12837" *)
  wire _03923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12865" *)
  wire _03924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12893" *)
  wire _03925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12921" *)
  wire _03926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12949" *)
  wire _03927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12977" *)
  wire _03928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13005" *)
  wire _03929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13033" *)
  wire _03930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14473" *)
  wire _03931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14682" *)
  wire _03932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14748" *)
  wire _03933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14767" *)
  wire _03934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16303" *)
  wire _03935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16311" *)
  wire _03936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16319" *)
  wire _03937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16327" *)
  wire _03938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16335" *)
  wire _03939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16343" *)
  wire _03940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16351" *)
  wire _03941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16359" *)
  wire _03942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16367" *)
  wire _03943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16375" *)
  wire _03944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16383" *)
  wire _03945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16392" *)
  wire _03946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16400" *)
  wire _03947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16408" *)
  wire _03948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16416" *)
  wire _03949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16424" *)
  wire _03950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *)
  wire _03951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *)
  wire _03952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *)
  wire _03953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *)
  wire _03954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *)
  wire _03955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *)
  wire _03956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *)
  wire _03957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *)
  wire _03958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *)
  wire _03959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *)
  wire _03960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *)
  wire _03961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *)
  wire _03962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *)
  wire _03963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18754" *)
  wire _03964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18759" *)
  wire _03965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18762" *)
  wire _03966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18765" *)
  wire _03967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18768" *)
  wire _03968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18771" *)
  wire _03969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18774" *)
  wire _03970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18777" *)
  wire _03971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18780" *)
  wire _03972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18783" *)
  wire _03973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18786" *)
  wire _03974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18789" *)
  wire _03975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18792" *)
  wire _03976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18795" *)
  wire _03977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18798" *)
  wire _03978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18801" *)
  wire _03979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *)
  wire _03980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23360" *)
  wire _03981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23387" *)
  wire _03982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23406" *)
  wire _03983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23420" *)
  wire _03984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23429" *)
  wire _03985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23447" *)
  wire _03986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23459" *)
  wire _03987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23475" *)
  wire _03988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23493" *)
  wire _03989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23504" *)
  wire _03990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23516" *)
  wire _03991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23537" *)
  wire _03992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23546" *)
  wire _03993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23567" *)
  wire _03994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23576" *)
  wire _03995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23585" *)
  wire _03996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24099" *)
  wire _03997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24110" *)
  wire _03998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24119" *)
  wire _03999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9129" *)
  wire _04000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16437" *)
  wire [48:0] _04001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16439" *)
  wire [48:0] _04002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16441" *)
  wire [48:0] _04003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16496" *)
  wire [48:0] _04004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16515" *)
  wire [48:0] _04005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10064" *)
  wire _04006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10819" *)
  wire _04007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10831" *)
  wire _04008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10846" *)
  wire _04009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10874" *)
  wire _04010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10928" *)
  wire _04011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11410" *)
  wire _04012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11412" *)
  wire _04013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11415" *)
  wire _04014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11418" *)
  wire _04015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11421" *)
  wire _04016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11423" *)
  wire _04017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11425" *)
  wire _04018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11427" *)
  wire _04019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11429" *)
  wire _04020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11432" *)
  wire _04021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11435" *)
  wire _04022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11523" *)
  wire _04023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11524" *)
  wire _04024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11530" *)
  wire _04025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11531" *)
  wire _04026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11537" *)
  wire _04027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11538" *)
  wire _04028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11544" *)
  wire _04029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11545" *)
  wire _04030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11551" *)
  wire _04031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11552" *)
  wire _04032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11558" *)
  wire _04033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11559" *)
  wire _04034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11565" *)
  wire _04035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11566" *)
  wire _04036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11572" *)
  wire _04037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11573" *)
  wire _04038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11579" *)
  wire _04039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11580" *)
  wire _04040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11586" *)
  wire _04041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11587" *)
  wire _04042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11593" *)
  wire _04043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11594" *)
  wire _04044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11605" *)
  wire _04045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11607" *)
  wire _04046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11608" *)
  wire _04047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11614" *)
  wire _04048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11615" *)
  wire _04049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11621" *)
  wire _04050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11622" *)
  wire _04051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11628" *)
  wire _04052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11629" *)
  wire _04053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11759" *)
  wire _04054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11765" *)
  wire _04055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11771" *)
  wire _04056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11777" *)
  wire _04057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11783" *)
  wire _04058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11789" *)
  wire _04059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11795" *)
  wire _04060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11801" *)
  wire _04061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11810" *)
  wire _04062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11816" *)
  wire _04063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11825" *)
  wire _04064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11831" *)
  wire _04065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11837" *)
  wire _04066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11843" *)
  wire _04067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11849" *)
  wire _04068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11855" *)
  wire _04069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11935" *)
  wire _04070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11983" *)
  wire _04071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12023" *)
  wire _04072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12071" *)
  wire _04073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12119" *)
  wire _04074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12159" *)
  wire _04075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12199" *)
  wire _04076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12247" *)
  wire _04077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12295" *)
  wire _04078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12335" *)
  wire _04079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12383" *)
  wire _04080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12431" *)
  wire _04081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12471" *)
  wire _04082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12511" *)
  wire _04083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12551" *)
  wire _04084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12591" *)
  wire _04085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12615" *)
  wire _04086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12643" *)
  wire _04087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12671" *)
  wire _04088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12699" *)
  wire _04089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12727" *)
  wire _04090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12755" *)
  wire _04091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12783" *)
  wire _04092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12811" *)
  wire _04093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12839" *)
  wire _04094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12867" *)
  wire _04095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12895" *)
  wire _04096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12923" *)
  wire _04097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12951" *)
  wire _04098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12979" *)
  wire _04099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13007" *)
  wire _04100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13035" *)
  wire _04101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13527" *)
  wire _04102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13528" *)
  wire _04103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13529" *)
  wire _04104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13543" *)
  wire _04105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13544" *)
  wire _04106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13545" *)
  wire _04107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13559" *)
  wire _04108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13560" *)
  wire _04109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13561" *)
  wire _04110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13575" *)
  wire _04111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13576" *)
  wire _04112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13577" *)
  wire _04113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13591" *)
  wire _04114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13592" *)
  wire _04115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13593" *)
  wire _04116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13607" *)
  wire _04117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13608" *)
  wire _04118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13609" *)
  wire _04119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13623" *)
  wire _04120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13624" *)
  wire _04121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13625" *)
  wire _04122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13639" *)
  wire _04123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13640" *)
  wire _04124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13641" *)
  wire _04125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13655" *)
  wire _04126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13656" *)
  wire _04127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13657" *)
  wire _04128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13671" *)
  wire _04129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13672" *)
  wire _04130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13673" *)
  wire _04131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13687" *)
  wire _04132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13688" *)
  wire _04133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13689" *)
  wire _04134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13703" *)
  wire _04135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13704" *)
  wire _04136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13705" *)
  wire _04137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13719" *)
  wire _04138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13720" *)
  wire _04139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13721" *)
  wire _04140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13735" *)
  wire _04141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13736" *)
  wire _04142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13737" *)
  wire _04143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13751" *)
  wire _04144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13752" *)
  wire _04145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13753" *)
  wire _04146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13767" *)
  wire _04147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13768" *)
  wire _04148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13769" *)
  wire _04149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14501" *)
  wire _04150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14525" *)
  wire _04151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16667" *)
  wire _04152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16669" *)
  wire _04153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16671" *)
  wire _04154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16673" *)
  wire _04155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16675" *)
  wire _04156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16677" *)
  wire _04157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16679" *)
  wire _04158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16681" *)
  wire _04159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16683" *)
  wire _04160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16685" *)
  wire _04161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16687" *)
  wire _04162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16689" *)
  wire _04163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16691" *)
  wire _04164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22924" *)
  wire _04165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23307" *)
  wire _04166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23326" *)
  wire _04167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23629" *)
  wire _04168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24092" *)
  wire _04169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24105" *)
  wire _04170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24114" *)
  wire _04171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8776" *)
  wire _04172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *)
  wire _04173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10000" *)
  wire _04174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10004" *)
  wire _04175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10010" *)
  wire _04176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10016" *)
  wire _04177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10022" *)
  wire _04178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10028" *)
  wire _04179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10034" *)
  wire _04180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10040" *)
  wire _04181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10046" *)
  wire _04182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10052" *)
  wire _04183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10058" *)
  wire _04184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *)
  wire _04185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *)
  wire _04186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10076" *)
  wire _04187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10081" *)
  wire _04188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10104" *)
  wire _04189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10140" *)
  wire [7:0] _04190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10153" *)
  wire [7:0] _04191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10165" *)
  wire [7:0] _04192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10177" *)
  wire [7:0] _04193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10189" *)
  wire [7:0] _04194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10201" *)
  wire [7:0] _04195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10213" *)
  wire [7:0] _04196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10225" *)
  wire [7:0] _04197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10237" *)
  wire [7:0] _04198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10249" *)
  wire [7:0] _04199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10261" *)
  wire [7:0] _04200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10273" *)
  wire [7:0] _04201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10285" *)
  wire [7:0] _04202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10297" *)
  wire [7:0] _04203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10309" *)
  wire [7:0] _04204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10321" *)
  wire [7:0] _04205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10402" *)
  wire _04206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10428" *)
  wire _04207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10454" *)
  wire _04208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10480" *)
  wire _04209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10506" *)
  wire _04210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10532" *)
  wire _04211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10558" *)
  wire _04212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10584" *)
  wire _04213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10610" *)
  wire _04214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10636" *)
  wire _04215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10662" *)
  wire _04216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10688" *)
  wire _04217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10714" *)
  wire _04218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10740" *)
  wire _04219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10766" *)
  wire _04220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10792" *)
  wire _04221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10817" *)
  wire _04222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10829" *)
  wire _04223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10844" *)
  wire _04224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10856" *)
  wire _04225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10872" *)
  wire _04226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10884" *)
  wire _04227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10897" *)
  wire _04228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10907" *)
  wire _04229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10926" *)
  wire _04230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10938" *)
  wire _04231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10948" *)
  wire _04232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10958" *)
  wire _04233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10968" *)
  wire _04234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10978" *)
  wire _04235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10988" *)
  wire _04236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10998" *)
  wire _04237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11006" *)
  wire _04238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11008" *)
  wire _04239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11011" *)
  wire [9:0] _04240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11016" *)
  wire _04241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11018" *)
  wire _04242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11021" *)
  wire [9:0] _04243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11026" *)
  wire _04244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11032" *)
  wire _04245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11035" *)
  wire [9:0] _04246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11039" *)
  wire _04247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11041" *)
  wire _04248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11044" *)
  wire [9:0] _04249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11048" *)
  wire _04250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11054" *)
  wire _04251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11057" *)
  wire [9:0] _04252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11061" *)
  wire _04253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11063" *)
  wire _04254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11066" *)
  wire [9:0] _04255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11070" *)
  wire _04256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11072" *)
  wire _04257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11075" *)
  wire [9:0] _04258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11079" *)
  wire _04259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11085" *)
  wire _04260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11088" *)
  wire [9:0] _04261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11093" *)
  wire _04262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11095" *)
  wire _04263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11098" *)
  wire [9:0] _04264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11102" *)
  wire _04265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11104" *)
  wire _04266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11107" *)
  wire [9:0] _04267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11111" *)
  wire _04268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11113" *)
  wire _04269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11116" *)
  wire [9:0] _04270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11120" *)
  wire _04271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11122" *)
  wire _04272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11125" *)
  wire [9:0] _04273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11129" *)
  wire _04274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11135" *)
  wire _04275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11138" *)
  wire [9:0] _04276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11142" *)
  wire _04277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11144" *)
  wire _04278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11147" *)
  wire [9:0] _04279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11151" *)
  wire _04280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11153" *)
  wire _04281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11156" *)
  wire [9:0] _04282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11160" *)
  wire _04283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11162" *)
  wire _04284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11165" *)
  wire [9:0] _04285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11235" *)
  wire _04286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11260" *)
  wire _04287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11261" *)
  wire _04288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11280" *)
  wire _04289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11281" *)
  wire _04290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11294" *)
  wire _04291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11295" *)
  wire _04292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11308" *)
  wire _04293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11309" *)
  wire _04294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11322" *)
  wire _04295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11323" *)
  wire _04296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11336" *)
  wire _04297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11337" *)
  wire _04298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11350" *)
  wire _04299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11351" *)
  wire _04300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11364" *)
  wire _04301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11365" *)
  wire _04302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11378" *)
  wire _04303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11379" *)
  wire _04304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11392" *)
  wire _04305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11393" *)
  wire _04306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11406" *)
  wire _04307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11407" *)
  wire _04308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11523" *)
  wire _04309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11526" *)
  wire _04310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11530" *)
  wire _04311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11533" *)
  wire _04312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11537" *)
  wire _04313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11540" *)
  wire _04314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11544" *)
  wire _04315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11547" *)
  wire _04316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11551" *)
  wire _04317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11554" *)
  wire _04318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11558" *)
  wire _04319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11561" *)
  wire _04320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11565" *)
  wire _04321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11568" *)
  wire _04322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11572" *)
  wire _04323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11575" *)
  wire _04324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11579" *)
  wire _04325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11582" *)
  wire _04326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11586" *)
  wire _04327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11589" *)
  wire _04328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11593" *)
  wire _04329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11596" *)
  wire _04330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11601" *)
  wire _04331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11607" *)
  wire _04332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11610" *)
  wire _04333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11614" *)
  wire _04334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11617" *)
  wire _04335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11621" *)
  wire _04336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11624" *)
  wire _04337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11628" *)
  wire _04338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11631" *)
  wire _04339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11639" *)
  wire _04340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *)
  wire _04341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *)
  wire _04342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11645" *)
  wire _04343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *)
  wire _04344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *)
  wire _04345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11651" *)
  wire _04346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *)
  wire _04347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *)
  wire _04348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11657" *)
  wire _04349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *)
  wire _04350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *)
  wire _04351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11663" *)
  wire _04352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *)
  wire _04353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *)
  wire _04354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11669" *)
  wire _04355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *)
  wire _04356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *)
  wire _04357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11675" *)
  wire _04358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *)
  wire _04359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *)
  wire _04360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11681" *)
  wire _04361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *)
  wire _04362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *)
  wire _04363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11687" *)
  wire _04364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *)
  wire _04365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *)
  wire _04366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11693" *)
  wire _04367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *)
  wire _04368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *)
  wire _04369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11700" *)
  wire _04370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *)
  wire _04371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *)
  wire _04372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11707" *)
  wire _04373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *)
  wire _04374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *)
  wire _04375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11714" *)
  wire _04376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *)
  wire _04377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *)
  wire _04378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11721" *)
  wire _04379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *)
  wire _04380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *)
  wire _04381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11728" *)
  wire _04382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *)
  wire _04383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *)
  wire _04384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11735" *)
  wire _04385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *)
  wire _04386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *)
  wire _04387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11738" *)
  wire _04388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11928" *)
  wire _04389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11933" *)
  wire _04390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11935" *)
  wire _04391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11976" *)
  wire _04392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11981" *)
  wire _04393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11983" *)
  wire _04394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12016" *)
  wire _04395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12021" *)
  wire _04396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12023" *)
  wire _04397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12064" *)
  wire _04398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12069" *)
  wire _04399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12071" *)
  wire _04400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12112" *)
  wire _04401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12117" *)
  wire _04402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12119" *)
  wire _04403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12152" *)
  wire _04404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12157" *)
  wire _04405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12159" *)
  wire _04406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12192" *)
  wire _04407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12197" *)
  wire _04408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12199" *)
  wire _04409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12240" *)
  wire _04410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12245" *)
  wire _04411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12247" *)
  wire _04412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12288" *)
  wire _04413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12293" *)
  wire _04414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12295" *)
  wire _04415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12328" *)
  wire _04416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12333" *)
  wire _04417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12335" *)
  wire _04418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12376" *)
  wire _04419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12381" *)
  wire _04420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12383" *)
  wire _04421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12424" *)
  wire _04422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12429" *)
  wire _04423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12431" *)
  wire _04424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12464" *)
  wire _04425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12469" *)
  wire _04426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12471" *)
  wire _04427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12504" *)
  wire _04428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12509" *)
  wire _04429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12511" *)
  wire _04430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12544" *)
  wire _04431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12549" *)
  wire _04432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12551" *)
  wire _04433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12584" *)
  wire _04434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12589" *)
  wire _04435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12591" *)
  wire _04436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12608" *)
  wire _04437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12613" *)
  wire _04438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12615" *)
  wire _04439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12636" *)
  wire _04440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12641" *)
  wire _04441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12643" *)
  wire _04442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12664" *)
  wire _04443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12669" *)
  wire _04444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12671" *)
  wire _04445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12692" *)
  wire _04446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12697" *)
  wire _04447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12699" *)
  wire _04448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12720" *)
  wire _04449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12725" *)
  wire _04450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12727" *)
  wire _04451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12748" *)
  wire _04452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12753" *)
  wire _04453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12755" *)
  wire _04454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12776" *)
  wire _04455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12781" *)
  wire _04456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12783" *)
  wire _04457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12804" *)
  wire _04458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12809" *)
  wire _04459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12811" *)
  wire _04460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12832" *)
  wire _04461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12837" *)
  wire _04462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12839" *)
  wire _04463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12860" *)
  wire _04464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12865" *)
  wire _04465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12867" *)
  wire _04466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12888" *)
  wire _04467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12893" *)
  wire _04468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12895" *)
  wire _04469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12916" *)
  wire _04470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12921" *)
  wire _04471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12923" *)
  wire _04472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12944" *)
  wire _04473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12949" *)
  wire _04474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12951" *)
  wire _04475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12972" *)
  wire _04476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12977" *)
  wire _04477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12979" *)
  wire _04478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13000" *)
  wire _04479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13005" *)
  wire _04480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13007" *)
  wire _04481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13028" *)
  wire _04482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13033" *)
  wire _04483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13035" *)
  wire _04484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13041" *)
  wire [3:0] _04485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13050" *)
  wire [3:0] _04486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13059" *)
  wire [3:0] _04487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13068" *)
  wire [3:0] _04488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13077" *)
  wire [3:0] _04489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13086" *)
  wire [3:0] _04490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13095" *)
  wire [3:0] _04491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13104" *)
  wire [3:0] _04492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13113" *)
  wire [3:0] _04493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13122" *)
  wire [3:0] _04494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13131" *)
  wire [3:0] _04495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13140" *)
  wire [3:0] _04496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13149" *)
  wire [3:0] _04497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13158" *)
  wire [3:0] _04498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13167" *)
  wire [3:0] _04499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13176" *)
  wire [3:0] _04500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13195" *)
  wire _04501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13209" *)
  wire _04502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13227" *)
  wire _04503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13240" *)
  wire _04504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13254" *)
  wire _04505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13268" *)
  wire _04506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13282" *)
  wire _04507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13296" *)
  wire _04508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13310" *)
  wire _04509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13324" *)
  wire _04510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13338" *)
  wire _04511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13352" *)
  wire _04512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13366" *)
  wire _04513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13375" *)
  wire _04514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13389" *)
  wire _04515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13403" *)
  wire _04516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13412" *)
  wire _04517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13416" *)
  wire [14:0] _04518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13417" *)
  wire _04519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13421" *)
  wire [14:0] _04520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13422" *)
  wire _04521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13426" *)
  wire [14:0] _04522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13427" *)
  wire _04523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13431" *)
  wire [14:0] _04524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13432" *)
  wire _04525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13436" *)
  wire [14:0] _04526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13437" *)
  wire _04527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13441" *)
  wire [14:0] _04528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13442" *)
  wire _04529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13446" *)
  wire [14:0] _04530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13447" *)
  wire _04531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13451" *)
  wire [14:0] _04532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13452" *)
  wire _04533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13456" *)
  wire [14:0] _04534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13457" *)
  wire _04535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13461" *)
  wire [14:0] _04536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13462" *)
  wire _04537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13466" *)
  wire [14:0] _04538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13467" *)
  wire _04539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13471" *)
  wire [14:0] _04540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13472" *)
  wire _04541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13476" *)
  wire [14:0] _04542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13477" *)
  wire _04543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13481" *)
  wire [14:0] _04544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13482" *)
  wire _04545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13486" *)
  wire [14:0] _04546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13487" *)
  wire _04547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13491" *)
  wire [14:0] _04548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13492" *)
  wire _04549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13790" *)
  wire _04550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13798" *)
  wire _04551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13806" *)
  wire _04552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13814" *)
  wire _04553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13822" *)
  wire _04554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13830" *)
  wire _04555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13838" *)
  wire _04556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13846" *)
  wire _04557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13854" *)
  wire _04558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13862" *)
  wire _04559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13870" *)
  wire _04560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13878" *)
  wire _04561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13886" *)
  wire _04562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13894" *)
  wire _04563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13902" *)
  wire _04564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13910" *)
  wire _04565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14072" *)
  wire _04566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14107" *)
  wire _04567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14111" *)
  wire _04568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14121" *)
  wire _04569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14131" *)
  wire _04570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14136" *)
  wire _04571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14139" *)
  wire _04572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14143" *)
  wire _04573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14145" *)
  wire _04574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14153" *)
  wire _04575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14156" *)
  wire _04576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14174" *)
  wire _04577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14184" *)
  wire _04578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14186" *)
  wire _04579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *)
  wire _04580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14204" *)
  wire _04581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14214" *)
  wire _04582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14225" *)
  wire _04583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14229" *)
  wire _04584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14273" *)
  wire _04585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14278" *)
  wire _04586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14284" *)
  wire _04587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14286" *)
  wire _04588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14288" *)
  wire _04589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14290" *)
  wire _04590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14306" *)
  wire _04591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14317" *)
  wire _04592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14347" *)
  wire _04593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14349" *)
  wire _04594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14354" *)
  wire _04595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14356" *)
  wire _04596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14358" *)
  wire _04597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14364" *)
  wire _04598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14368" *)
  wire _04599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14370" *)
  wire _04600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14374" *)
  wire _04601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14376" *)
  wire _04602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14378" *)
  wire _04603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14382" *)
  wire _04604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14384" *)
  wire _04605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14390" *)
  wire _04606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14392" *)
  wire _04607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14397" *)
  wire _04608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14399" *)
  wire _04609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14401" *)
  wire _04610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14407" *)
  wire _04611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14413" *)
  wire _04612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14415" *)
  wire _04613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14417" *)
  wire _04614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14419" *)
  wire _04615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14423" *)
  wire _04616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14425" *)
  wire _04617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14427" *)
  wire _04618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14437" *)
  wire _04619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14441" *)
  wire _04620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14443" *)
  wire _04621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14445" *)
  wire _04622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14447" *)
  wire _04623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14449" *)
  wire _04624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14453" *)
  wire _04625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14455" *)
  wire _04626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14457" *)
  wire _04627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14459" *)
  wire _04628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14467" *)
  wire _04629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14469" *)
  wire _04630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14471" *)
  wire _04631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14490" *)
  wire _04632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14494" *)
  wire _04633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14500" *)
  wire _04634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14504" *)
  wire _04635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14507" *)
  wire _04636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14513" *)
  wire _04637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14522" *)
  wire _04638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14527" *)
  wire _04639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14540" *)
  wire _04640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14546" *)
  wire _04641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14559" *)
  wire _04642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14566" *)
  wire _04643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14568" *)
  wire _04644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14607" *)
  wire _04645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14624" *)
  wire _04646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14625" *)
  wire _04647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14675" *)
  wire _04648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14684" *)
  wire _04649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14737" *)
  wire _04650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14742" *)
  wire _04651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14750" *)
  wire _04652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14764" *)
  wire _04653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14767" *)
  wire _04654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14788" *)
  wire _04655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14789" *)
  wire _04656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14790" *)
  wire _04657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14791" *)
  wire _04658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14792" *)
  wire _04659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14793" *)
  wire _04660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14794" *)
  wire _04661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14795" *)
  wire _04662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14796" *)
  wire _04663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14797" *)
  wire _04664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14798" *)
  wire _04665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14799" *)
  wire _04666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14800" *)
  wire _04667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14801" *)
  wire _04668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14802" *)
  wire _04669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14803" *)
  wire _04670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14804" *)
  wire _04671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14805" *)
  wire _04672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14806" *)
  wire _04673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14807" *)
  wire _04674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14808" *)
  wire _04675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14809" *)
  wire _04676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14810" *)
  wire _04677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14811" *)
  wire _04678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14812" *)
  wire _04679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14813" *)
  wire _04680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14814" *)
  wire _04681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14815" *)
  wire _04682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14816" *)
  wire _04683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14817" *)
  wire _04684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14818" *)
  wire _04685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14819" *)
  wire _04686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14849" *)
  wire _04687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14854" *)
  wire _04688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14859" *)
  wire _04689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14862" *)
  wire _04690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14881" *)
  wire _04691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14883" *)
  wire _04692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14886" *)
  wire _04693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *)
  wire _04694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14983" *)
  wire _04695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *)
  wire _04696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14990" *)
  wire _04697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14992" *)
  wire _04698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15056" *)
  wire _04699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15057" *)
  wire _04700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15058" *)
  wire _04701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15059" *)
  wire _04702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15060" *)
  wire _04703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15061" *)
  wire _04704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15062" *)
  wire _04705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15063" *)
  wire _04706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15064" *)
  wire _04707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15065" *)
  wire _04708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15066" *)
  wire _04709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15067" *)
  wire _04710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15068" *)
  wire _04711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15069" *)
  wire _04712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15070" *)
  wire _04713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15071" *)
  wire _04714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15072" *)
  wire _04715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15073" *)
  wire _04716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15074" *)
  wire _04717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15075" *)
  wire _04718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15076" *)
  wire _04719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15077" *)
  wire _04720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15078" *)
  wire _04721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15079" *)
  wire _04722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15080" *)
  wire _04723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15081" *)
  wire _04724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15082" *)
  wire _04725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15083" *)
  wire _04726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15084" *)
  wire _04727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15085" *)
  wire _04728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15086" *)
  wire _04729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15087" *)
  wire _04730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15094" *)
  wire _04731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15094" *)
  wire _04732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15369" *)
  wire _04733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15383" *)
  wire _04734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15396" *)
  wire _04735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15410" *)
  wire _04736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15424" *)
  wire _04737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15438" *)
  wire _04738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15452" *)
  wire _04739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15466" *)
  wire _04740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15480" *)
  wire _04741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15622" *)
  wire _04742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15630" *)
  wire _04743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15654" *)
  wire _04744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15664" *)
  wire _04745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15726" *)
  wire _04746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15736" *)
  wire _04747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15754" *)
  wire _04748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15764" *)
  wire _04749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15782" *)
  wire _04750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15792" *)
  wire _04751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15801" *)
  wire _04752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15810" *)
  wire _04753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15820" *)
  wire _04754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15829" *)
  wire _04755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15838" *)
  wire _04756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15848" *)
  wire _04757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15857" *)
  wire _04758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15866" *)
  wire _04759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15876" *)
  wire _04760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15894" *)
  wire _04761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15904" *)
  wire _04762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15922" *)
  wire _04763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15932" *)
  wire _04764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15941" *)
  wire _04765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15950" *)
  wire _04766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15960" *)
  wire _04767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15978" *)
  wire _04768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15988" *)
  wire _04769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16006" *)
  wire _04770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16016" *)
  wire _04771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16025" *)
  wire _04772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16034" *)
  wire _04773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16044" *)
  wire _04774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16062" *)
  wire _04775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16072" *)
  wire _04776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16090" *)
  wire _04777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16100" *)
  wire _04778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16118" *)
  wire _04779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16128" *)
  wire _04780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *)
  wire _04781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *)
  wire _04782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *)
  wire _04783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *)
  wire _04784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *)
  wire _04785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *)
  wire _04786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *)
  wire _04787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *)
  wire _04788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *)
  wire _04789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *)
  wire _04790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *)
  wire _04791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *)
  wire _04792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *)
  wire _04793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *)
  wire _04794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *)
  wire _04795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *)
  wire _04796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *)
  wire _04797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *)
  wire _04798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *)
  wire _04799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *)
  wire _04800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *)
  wire _04801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *)
  wire _04802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *)
  wire _04803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *)
  wire _04804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *)
  wire _04805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *)
  wire _04806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *)
  wire _04807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *)
  wire _04808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *)
  wire _04809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *)
  wire _04810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *)
  wire _04811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *)
  wire _04812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16523" *)
  wire _04813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16667" *)
  wire _04814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *)
  wire _04815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *)
  wire _04816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16669" *)
  wire _04817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *)
  wire _04818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *)
  wire _04819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16671" *)
  wire _04820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *)
  wire _04821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *)
  wire _04822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16673" *)
  wire _04823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *)
  wire _04824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *)
  wire _04825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16675" *)
  wire _04826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *)
  wire _04827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *)
  wire _04828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16677" *)
  wire _04829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *)
  wire _04830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *)
  wire _04831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16679" *)
  wire _04832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *)
  wire _04833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *)
  wire _04834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16681" *)
  wire _04835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *)
  wire _04836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *)
  wire _04837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16683" *)
  wire _04838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *)
  wire _04839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *)
  wire _04840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16685" *)
  wire _04841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *)
  wire _04842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *)
  wire _04843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16687" *)
  wire _04844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *)
  wire _04845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *)
  wire _04846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16689" *)
  wire _04847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *)
  wire _04848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *)
  wire _04849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16691" *)
  wire _04850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *)
  wire _04851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *)
  wire _04852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16792" *)
  wire _04853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16942" *)
  wire _04854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16961" *)
  wire _04855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17000" *)
  wire _04856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17209" *)
  wire _04857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17257" *)
  wire _04858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17265" *)
  wire _04859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17333" *)
  wire _04860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17395" *)
  wire _04861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17443" *)
  wire _04862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17451" *)
  wire _04863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17569" *)
  wire _04864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17617" *)
  wire _04865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17675" *)
  wire _04866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *)
  wire _04867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17723" *)
  wire _04868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17790" *)
  wire _04869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17838" *)
  wire _04870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17846" *)
  wire _04871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17894" *)
  wire _04872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17902" *)
  wire _04873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17955" *)
  wire _04874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18532" *)
  wire _04875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18755" *)
  wire _04876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18760" *)
  wire _04877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18763" *)
  wire _04878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18766" *)
  wire _04879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18769" *)
  wire _04880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18772" *)
  wire _04881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18775" *)
  wire _04882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18778" *)
  wire _04883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18781" *)
  wire _04884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18784" *)
  wire _04885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18787" *)
  wire _04886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18790" *)
  wire _04887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18793" *)
  wire _04888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18796" *)
  wire _04889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18799" *)
  wire _04890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18802" *)
  wire _04891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18882" *)
  wire _04892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18883" *)
  wire _04893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18899" *)
  wire _04894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18900" *)
  wire _04895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18938" *)
  wire _04896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18959" *)
  wire _04897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18988" *)
  wire _04898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18989" *)
  wire _04899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18990" *)
  wire _04900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *)
  wire _04901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18998" *)
  wire _04902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18999" *)
  wire _04903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19028" *)
  wire _04904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *)
  wire _04905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19039" *)
  wire _04906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19060" *)
  wire _04907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19061" *)
  wire _04908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19062" *)
  wire _04909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19063" *)
  wire _04910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19064" *)
  wire _04911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19065" *)
  wire _04912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *)
  wire _04913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19074" *)
  wire _04914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19104" *)
  wire _04915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19115" *)
  wire _04916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19116" *)
  wire _04917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *)
  wire _04918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19166" *)
  wire _04919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19177" *)
  wire _04920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19178" *)
  wire _04921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19197" *)
  wire _04922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19208" *)
  wire _04923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19209" *)
  wire _04924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19228" *)
  wire _04925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19239" *)
  wire _04926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19240" *)
  wire _04927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19259" *)
  wire _04928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19260" *)
  wire _04929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19261" *)
  wire _04930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *)
  wire _04931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19270" *)
  wire _04932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19310" *)
  wire _04933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19311" *)
  wire _04934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19329" *)
  wire _04935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19341" *)
  wire _04936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19342" *)
  wire _04937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19360" *)
  wire _04938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19372" *)
  wire _04939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19373" *)
  wire _04940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19405" *)
  wire _04941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19406" *)
  wire _04942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19424" *)
  wire _04943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19432" *)
  wire _04944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19442" *)
  wire _04945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19443" *)
  wire _04946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19461" *)
  wire _04947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19492" *)
  wire _04948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19493" *)
  wire _04949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19513" *)
  wire _04950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19514" *)
  wire _04951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19576" *)
  wire _04952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19577" *)
  wire _04953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19586" *)
  wire _04954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19805" *)
  wire _04955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20069" *)
  wire _04956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *)
  wire _04957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20088" *)
  wire _04958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20107" *)
  wire _04959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20126" *)
  wire _04960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20145" *)
  wire _04961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20164" *)
  wire _04962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20202" *)
  wire _04963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20221" *)
  wire _04964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20240" *)
  wire _04965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20278" *)
  wire _04966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20297" *)
  wire _04967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20316" *)
  wire _04968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20335" *)
  wire _04969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20354" *)
  wire _04970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20581" *)
  wire _04971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20583" *)
  wire _04972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20585" *)
  wire _04973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20587" *)
  wire _04974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20589" *)
  wire _04975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20591" *)
  wire _04976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20593" *)
  wire _04977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20595" *)
  wire _04978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20597" *)
  wire _04979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20599" *)
  wire _04980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20601" *)
  wire _04981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20603" *)
  wire _04982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20605" *)
  wire _04983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20607" *)
  wire _04984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20609" *)
  wire _04985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *)
  wire _04986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *)
  wire _04987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *)
  wire _04988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *)
  wire _04989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *)
  wire _04990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *)
  wire _04991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *)
  wire _04992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *)
  wire _04993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20903" *)
  wire _04994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20913" *)
  wire _04995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *)
  wire _04996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *)
  wire _04997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *)
  wire _04998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *)
  wire _04999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *)
  wire _05000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *)
  wire _05001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20978" *)
  wire _05002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20988" *)
  wire _05003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *)
  wire _05004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *)
  wire _05005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *)
  wire _05006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *)
  wire _05007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *)
  wire _05008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *)
  wire _05009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *)
  wire _05010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *)
  wire _05011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *)
  wire _05012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *)
  wire _05013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *)
  wire _05014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *)
  wire _05015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *)
  wire _05016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *)
  wire _05017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21152" *)
  wire _05018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *)
  wire _05019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *)
  wire _05020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21179" *)
  wire _05021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *)
  wire _05022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *)
  wire _05023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *)
  wire _05024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *)
  wire _05025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *)
  wire _05026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *)
  wire _05027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *)
  wire _05028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *)
  wire _05029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *)
  wire _05030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *)
  wire _05031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *)
  wire _05032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *)
  wire _05033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *)
  wire _05034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *)
  wire _05035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *)
  wire _05036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *)
  wire _05037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *)
  wire _05038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *)
  wire _05039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21417" *)
  wire _05040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21420" *)
  wire _05041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21423" *)
  wire _05042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21426" *)
  wire _05043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21462" *)
  wire _05044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21467" *)
  wire _05045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21474" *)
  wire _05046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21480" *)
  wire _05047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21485" *)
  wire _05048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21493" *)
  wire _05049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21499" *)
  wire _05050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21504" *)
  wire _05051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21512" *)
  wire _05052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21517" *)
  wire _05053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21522" *)
  wire _05054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21528" *)
  wire _05055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21547" *)
  wire _05056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21574" *)
  wire _05057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21600" *)
  wire _05058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21627" *)
  wire _05059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21654" *)
  wire _05060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21681" *)
  wire _05061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21708" *)
  wire _05062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21735" *)
  wire _05063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21762" *)
  wire _05064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21789" *)
  wire _05065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21816" *)
  wire _05066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21843" *)
  wire _05067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21870" *)
  wire _05068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21920" *)
  wire _05069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21935" *)
  wire _05070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21963" *)
  wire _05071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21967" *)
  wire _05072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21970" *)
  wire _05073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21971" *)
  wire _05074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *)
  wire _05075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21982" *)
  wire _05076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22008" *)
  wire _05077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22031" *)
  wire _05078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22054" *)
  wire _05079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22075" *)
  wire _05080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22104" *)
  wire _05081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22157" *)
  wire _05082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22180" *)
  wire _05083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22201" *)
  wire _05084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22234" *)
  wire _05085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22257" *)
  wire _05086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22278" *)
  wire _05087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22311" *)
  wire _05088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22334" *)
  wire _05089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22357" *)
  wire _05090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22590" *)
  wire _05091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22594" *)
  wire _05092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22597" *)
  wire _05093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22634" *)
  wire _05094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22637" *)
  wire _05095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22650" *)
  wire _05096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22653" *)
  wire _05097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22666" *)
  wire _05098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22669" *)
  wire _05099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22702" *)
  wire _05100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22705" *)
  wire _05101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22720" *)
  wire _05102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22723" *)
  wire _05103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22738" *)
  wire _05104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22741" *)
  wire _05105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22747" *)
  wire _05106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22753" *)
  wire _05107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22758" *)
  wire _05108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22761" *)
  wire _05109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22768" *)
  wire _05110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22781" *)
  wire _05111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22798" *)
  wire _05112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22801" *)
  wire _05113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22807" *)
  wire _05114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22811" *)
  wire _05115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22823" *)
  wire _05116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22826" *)
  wire _05117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22833" *)
  wire _05118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22837" *)
  wire _05119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22879" *)
  wire _05120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22882" *)
  wire _05121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22890" *)
  wire _05122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22895" *)
  wire _05123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22899" *)
  wire _05124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22901" *)
  wire _05125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22909" *)
  wire _05126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22916" *)
  wire _05127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *)
  wire _05128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *)
  wire _05129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *)
  wire _05130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22931" *)
  wire _05131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22935" *)
  wire _05132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22947" *)
  wire _05133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22951" *)
  wire _05134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22957" *)
  wire _05135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22962" *)
  wire _05136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22965" *)
  wire _05137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22969" *)
  wire _05138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22975" *)
  wire _05139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22977" *)
  wire _05140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22989" *)
  wire _05141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22994" *)
  wire _05142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22998" *)
  wire _05143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23016" *)
  wire _05144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23020" *)
  wire _05145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23026" *)
  wire _05146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23030" *)
  wire _05147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23036" *)
  wire _05148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23038" *)
  wire _05149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23050" *)
  wire _05150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23055" *)
  wire _05151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23059" *)
  wire _05152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23065" *)
  wire _05153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23067" *)
  wire _05154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23079" *)
  wire _05155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23084" *)
  wire _05156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23088" *)
  wire _05157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23095" *)
  wire _05158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *)
  wire _05159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *)
  wire _05160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *)
  wire _05161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *)
  wire _05162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *)
  wire _05163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *)
  wire _05164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23113" *)
  wire _05165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23113" *)
  wire _05166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23114" *)
  wire _05167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23117" *)
  wire _05168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23119" *)
  wire _05169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23132" *)
  wire _05170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23134" *)
  wire _05171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23138" *)
  wire _05172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23144" *)
  wire _05173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23146" *)
  wire _05174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23164" *)
  wire _05175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23168" *)
  wire _05176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23174" *)
  wire _05177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23178" *)
  wire _05178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23184" *)
  wire _05179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23188" *)
  wire _05180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23194" *)
  wire _05181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23198" *)
  wire _05182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23308" *)
  wire _05183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23309" *)
  wire _05184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23316" *)
  wire _05185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *)
  wire _05186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *)
  wire _05187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *)
  wire _05188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *)
  wire _05189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *)
  wire _05190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *)
  wire _05191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *)
  wire _05192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *)
  wire _05193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *)
  wire _05194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *)
  wire _05195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *)
  wire _05196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *)
  wire _05197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23360" *)
  wire _05198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *)
  wire _05199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23380" *)
  wire _05200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23380" *)
  wire _05201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23382" *)
  wire _05202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23387" *)
  wire _05203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *)
  wire _05204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *)
  wire _05205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23406" *)
  wire _05206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *)
  wire _05207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *)
  wire _05208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23420" *)
  wire _05209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *)
  wire _05210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *)
  wire _05211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23429" *)
  wire _05212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *)
  wire _05213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *)
  wire _05214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23447" *)
  wire _05215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *)
  wire _05216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *)
  wire _05217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23459" *)
  wire _05218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *)
  wire _05219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *)
  wire _05220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23475" *)
  wire _05221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *)
  wire _05222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *)
  wire _05223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23493" *)
  wire _05224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *)
  wire _05225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *)
  wire _05226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23504" *)
  wire _05227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *)
  wire _05228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *)
  wire _05229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23516" *)
  wire _05230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *)
  wire _05231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *)
  wire _05232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *)
  wire _05233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23530" *)
  wire _05234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23537" *)
  wire _05235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *)
  wire _05236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *)
  wire _05237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *)
  wire _05238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23546" *)
  wire _05239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *)
  wire _05240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *)
  wire _05241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23556" *)
  wire _05242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23562" *)
  wire _05243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23567" *)
  wire _05244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *)
  wire _05245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *)
  wire _05246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23576" *)
  wire _05247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *)
  wire _05248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *)
  wire _05249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23585" *)
  wire _05250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *)
  wire _05251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *)
  wire _05252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23595" *)
  wire _05253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23599" *)
  wire _05254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23620" *)
  wire _05255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23622" *)
  wire _05256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23625" *)
  wire _05257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23650" *)
  wire _05258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23651" *)
  wire _05259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23673" *)
  wire _05260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23674" *)
  wire _05261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23696" *)
  wire _05262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23697" *)
  wire _05263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23719" *)
  wire _05264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23720" *)
  wire _05265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23726" *)
  wire _05266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *)
  wire _05267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23742" *)
  wire _05268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23743" *)
  wire _05269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23765" *)
  wire _05270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23766" *)
  wire _05271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23788" *)
  wire _05272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23789" *)
  wire _05273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23811" *)
  wire _05274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23812" *)
  wire _05275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23834" *)
  wire _05276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23835" *)
  wire _05277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23857" *)
  wire _05278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23858" *)
  wire _05279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23880" *)
  wire _05280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23881" *)
  wire _05281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23903" *)
  wire _05282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23904" *)
  wire _05283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23926" *)
  wire _05284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23927" *)
  wire _05285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23949" *)
  wire _05286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23950" *)
  wire _05287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23972" *)
  wire _05288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23973" *)
  wire _05289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23995" *)
  wire _05290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23996" *)
  wire _05291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *)
  wire _05292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24063" *)
  wire _05293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24123" *)
  wire _05294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24125" *)
  wire _05295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24127" *)
  wire _05296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24132" *)
  wire _05297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24229" *)
  wire _05298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8774" *)
  wire _05299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8799" *)
  wire _05300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8821" *)
  wire _05301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8825" *)
  wire _05302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8830" *)
  wire _05303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8831" *)
  wire _05304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8841" *)
  wire _05305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8845" *)
  wire _05306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8846" *)
  wire _05307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8847" *)
  wire _05308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8848" *)
  wire _05309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8853" *)
  wire _05310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8854" *)
  wire _05311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8855" *)
  wire _05312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8856" *)
  wire _05313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8857" *)
  wire _05314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8858" *)
  wire _05315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8859" *)
  wire _05316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8861" *)
  wire _05317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8871" *)
  wire _05318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8882" *)
  wire _05319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8893" *)
  wire _05320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8947" *)
  wire _05321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8954" *)
  wire _05322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8966" *)
  wire _05323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8976" *)
  wire _05324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8979" *)
  wire _05325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9007" *)
  wire _05326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9011" *)
  wire _05327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9016" *)
  wire _05328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9045" *)
  wire _05329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9051" *)
  wire _05330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9071" *)
  wire _05331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9120" *)
  wire _05332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9125" *)
  wire _05333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9151" *)
  wire _05334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9156" *)
  wire _05335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9167" *)
  wire _05336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9169" *)
  wire _05337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9183" *)
  wire _05338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9188" *)
  wire _05339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9217" *)
  wire _05340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9243" *)
  wire _05341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9264" *)
  wire _05342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9276" *)
  wire _05343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9281" *)
  wire _05344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *)
  wire _05345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *)
  wire _05346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *)
  wire _05347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9301" *)
  wire _05348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9306" *)
  wire _05349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9333" *)
  wire _05350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9345" *)
  wire _05351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9350" *)
  wire _05352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9367" *)
  wire _05353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9381" *)
  wire _05354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9394" *)
  wire _05355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9399" *)
  wire _05356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9423" *)
  wire _05357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9428" *)
  wire _05358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9443" *)
  wire _05359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9448" *)
  wire _05360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9460" *)
  wire _05361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9465" *)
  wire _05362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9479" *)
  wire _05363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9481" *)
  wire _05364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9482" *)
  wire _05365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *)
  wire _05366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *)
  wire _05367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9495" *)
  wire _05368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9533" *)
  wire _05369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9554" *)
  wire _05370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9581" *)
  wire _05371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9595" *)
  wire _05372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9606" *)
  wire _05373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9627" *)
  wire _05374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9640" *)
  wire _05375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9656" *)
  wire _05376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9672" *)
  wire _05377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9688" *)
  wire _05378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9704" *)
  wire _05379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9721" *)
  wire _05380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9735" *)
  wire _05381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9769" *)
  wire _05382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9789" *)
  wire _05383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9838" *)
  wire _05384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9850" *)
  wire _05385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9861" *)
  wire _05386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9864" *)
  wire _05387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9869" *)
  wire _05388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9879" *)
  wire _05389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9884" *)
  wire _05390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9899" *)
  wire _05391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9901" *)
  wire _05392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9902" *)
  wire _05393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9905" *)
  wire _05394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9910" *)
  wire _05395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9913" *)
  wire _05396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9916" *)
  wire _05397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9968" *)
  wire _05398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9974" *)
  wire _05399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9980" *)
  wire _05400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9986" *)
  wire _05401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9992" *)
  wire _05402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9998" *)
  wire _05403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10002" *)
  wire _05404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10002" *)
  wire _05405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10008" *)
  wire _05406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10008" *)
  wire _05407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10014" *)
  wire _05408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10014" *)
  wire _05409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10020" *)
  wire _05410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10020" *)
  wire _05411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10026" *)
  wire _05412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10026" *)
  wire _05413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10032" *)
  wire _05414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10032" *)
  wire _05415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10038" *)
  wire _05416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10038" *)
  wire _05417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10044" *)
  wire _05418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10044" *)
  wire _05419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10050" *)
  wire _05420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10050" *)
  wire _05421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10056" *)
  wire _05422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10056" *)
  wire _05423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *)
  wire _05424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *)
  wire _05425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10064" *)
  wire _05426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10065" *)
  wire _05427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *)
  wire _05428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10106" *)
  wire _05429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10115" *)
  wire _05430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10809" *)
  wire _05431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10817" *)
  wire _05432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10819" *)
  wire _05433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10819" *)
  wire _05434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10821" *)
  wire _05435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10829" *)
  wire _05436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10831" *)
  wire _05437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10831" *)
  wire _05438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10836" *)
  wire _05439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10844" *)
  wire _05440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10846" *)
  wire _05441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10846" *)
  wire _05442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10856" *)
  wire _05443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10872" *)
  wire _05444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10874" *)
  wire _05445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10874" *)
  wire _05446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10884" *)
  wire _05447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10897" *)
  wire _05448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10907" *)
  wire _05449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10918" *)
  wire _05450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10926" *)
  wire _05451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10928" *)
  wire _05452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10928" *)
  wire _05453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10938" *)
  wire _05454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10948" *)
  wire _05455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10958" *)
  wire _05456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10968" *)
  wire _05457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10978" *)
  wire _05458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10988" *)
  wire _05459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10998" *)
  wire _05460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11006" *)
  wire _05461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11008" *)
  wire _05462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11016" *)
  wire _05463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11018" *)
  wire _05464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11026" *)
  wire _05465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11032" *)
  wire _05466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11039" *)
  wire _05467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11041" *)
  wire _05468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11048" *)
  wire _05469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11054" *)
  wire _05470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11061" *)
  wire _05471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11063" *)
  wire _05472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11070" *)
  wire _05473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11072" *)
  wire _05474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11079" *)
  wire _05475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11085" *)
  wire _05476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11093" *)
  wire _05477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11095" *)
  wire _05478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11102" *)
  wire _05479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11104" *)
  wire _05480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11111" *)
  wire _05481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11113" *)
  wire _05482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11120" *)
  wire _05483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11122" *)
  wire _05484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11129" *)
  wire _05485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11135" *)
  wire _05486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11142" *)
  wire _05487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11144" *)
  wire _05488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11151" *)
  wire _05489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11153" *)
  wire _05490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11160" *)
  wire _05491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11162" *)
  wire _05492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11262" *)
  wire _05493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11282" *)
  wire _05494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11296" *)
  wire _05495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11310" *)
  wire _05496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11324" *)
  wire _05497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11338" *)
  wire _05498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11352" *)
  wire _05499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11366" *)
  wire _05500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11380" *)
  wire _05501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11394" *)
  wire _05502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11408" *)
  wire _05503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11410" *)
  wire _05504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11410" *)
  wire _05505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11412" *)
  wire _05506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11413" *)
  wire _05507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11415" *)
  wire _05508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11416" *)
  wire _05509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11418" *)
  wire _05510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11419" *)
  wire _05511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11421" *)
  wire _05512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11421" *)
  wire _05513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11423" *)
  wire _05514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11423" *)
  wire _05515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11425" *)
  wire _05516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11425" *)
  wire _05517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11427" *)
  wire _05518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11427" *)
  wire _05519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11429" *)
  wire _05520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11430" *)
  wire _05521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11432" *)
  wire _05522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11433" *)
  wire _05523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11435" *)
  wire _05524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11436" *)
  wire _05525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11438" *)
  wire _05526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11438" *)
  wire _05527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11439" *)
  wire _05528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11439" *)
  wire _05529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11439" *)
  wire _05530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11440" *)
  wire _05531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11440" *)
  wire _05532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11440" *)
  wire _05533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *)
  wire _05534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *)
  wire _05535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *)
  wire _05536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *)
  wire _05537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11443" *)
  wire _05538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11443" *)
  wire _05539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11444" *)
  wire _05540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11444" *)
  wire _05541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11444" *)
  wire _05542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11445" *)
  wire _05543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11445" *)
  wire _05544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11445" *)
  wire _05545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *)
  wire _05546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *)
  wire _05547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *)
  wire _05548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *)
  wire _05549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11448" *)
  wire _05550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11448" *)
  wire _05551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11449" *)
  wire _05552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11449" *)
  wire _05553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11449" *)
  wire _05554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11450" *)
  wire _05555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11450" *)
  wire _05556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11450" *)
  wire _05557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *)
  wire _05558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *)
  wire _05559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *)
  wire _05560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *)
  wire _05561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11453" *)
  wire _05562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11453" *)
  wire _05563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11454" *)
  wire _05564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11454" *)
  wire _05565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11454" *)
  wire _05566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11455" *)
  wire _05567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11455" *)
  wire _05568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11455" *)
  wire _05569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *)
  wire _05570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *)
  wire _05571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *)
  wire _05572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *)
  wire _05573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11458" *)
  wire _05574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11458" *)
  wire _05575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11459" *)
  wire _05576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11459" *)
  wire _05577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11459" *)
  wire _05578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11460" *)
  wire _05579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11460" *)
  wire _05580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11460" *)
  wire _05581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *)
  wire _05582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *)
  wire _05583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *)
  wire _05584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *)
  wire _05585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11463" *)
  wire _05586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11463" *)
  wire _05587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11464" *)
  wire _05588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11464" *)
  wire _05589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11464" *)
  wire _05590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11465" *)
  wire _05591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11465" *)
  wire _05592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11465" *)
  wire _05593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *)
  wire _05594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *)
  wire _05595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *)
  wire _05596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *)
  wire _05597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11468" *)
  wire _05598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11468" *)
  wire _05599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11469" *)
  wire _05600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11469" *)
  wire _05601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11469" *)
  wire _05602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11470" *)
  wire _05603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11470" *)
  wire _05604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11470" *)
  wire _05605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *)
  wire _05606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *)
  wire _05607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *)
  wire _05608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *)
  wire _05609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11473" *)
  wire _05610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11473" *)
  wire _05611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11474" *)
  wire _05612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11474" *)
  wire _05613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11474" *)
  wire _05614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11475" *)
  wire _05615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11475" *)
  wire _05616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11475" *)
  wire _05617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *)
  wire _05618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *)
  wire _05619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *)
  wire _05620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *)
  wire _05621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11478" *)
  wire _05622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11478" *)
  wire _05623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11479" *)
  wire _05624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11479" *)
  wire _05625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11479" *)
  wire _05626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11480" *)
  wire _05627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11480" *)
  wire _05628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11480" *)
  wire _05629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *)
  wire _05630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *)
  wire _05631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *)
  wire _05632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *)
  wire _05633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11483" *)
  wire _05634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11484" *)
  wire _05635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11484" *)
  wire _05636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11484" *)
  wire _05637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11485" *)
  wire _05638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11485" *)
  wire _05639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11485" *)
  wire _05640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11486" *)
  wire _05641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11486" *)
  wire _05642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11486" *)
  wire _05643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11487" *)
  wire _05644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11487" *)
  wire _05645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11489" *)
  wire _05646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11490" *)
  wire _05647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11490" *)
  wire _05648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11490" *)
  wire _05649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11491" *)
  wire _05650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11491" *)
  wire _05651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11491" *)
  wire _05652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11492" *)
  wire _05653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11492" *)
  wire _05654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11492" *)
  wire _05655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11493" *)
  wire _05656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11493" *)
  wire _05657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11495" *)
  wire _05658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11496" *)
  wire _05659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11496" *)
  wire _05660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11496" *)
  wire _05661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11497" *)
  wire _05662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11497" *)
  wire _05663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11497" *)
  wire _05664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11498" *)
  wire _05665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11498" *)
  wire _05666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11498" *)
  wire _05667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11499" *)
  wire _05668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11499" *)
  wire _05669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11501" *)
  wire _05670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11502" *)
  wire _05671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11502" *)
  wire _05672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11502" *)
  wire _05673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11503" *)
  wire _05674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11503" *)
  wire _05675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11503" *)
  wire _05676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11504" *)
  wire _05677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11504" *)
  wire _05678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11504" *)
  wire _05679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11505" *)
  wire _05680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11505" *)
  wire _05681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11507" *)
  wire _05682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11508" *)
  wire _05683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11508" *)
  wire _05684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11508" *)
  wire _05685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11509" *)
  wire _05686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11509" *)
  wire _05687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11509" *)
  wire _05688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11510" *)
  wire _05689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11510" *)
  wire _05690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11510" *)
  wire _05691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11511" *)
  wire _05692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11511" *)
  wire _05693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11513" *)
  wire _05694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11514" *)
  wire _05695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11514" *)
  wire _05696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11514" *)
  wire _05697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11515" *)
  wire _05698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11515" *)
  wire _05699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11515" *)
  wire _05700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11516" *)
  wire _05701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11516" *)
  wire _05702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11516" *)
  wire _05703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11517" *)
  wire _05704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11517" *)
  wire _05705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11519" *)
  wire _05706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11519" *)
  wire _05707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11520" *)
  wire _05708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11520" *)
  wire _05709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11520" *)
  wire _05710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11521" *)
  wire _05711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11521" *)
  wire _05712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11521" *)
  wire _05713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *)
  wire _05714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *)
  wire _05715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *)
  wire _05716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *)
  wire _05717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11524" *)
  wire _05718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11531" *)
  wire _05719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11538" *)
  wire _05720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11545" *)
  wire _05721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11552" *)
  wire _05722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11559" *)
  wire _05723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11566" *)
  wire _05724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11573" *)
  wire _05725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11580" *)
  wire _05726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11587" *)
  wire _05727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11594" *)
  wire _05728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11608" *)
  wire _05729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11615" *)
  wire _05730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11622" *)
  wire _05731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11629" *)
  wire _05732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *)
  wire _05733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *)
  wire _05734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *)
  wire _05735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *)
  wire _05736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *)
  wire _05737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *)
  wire _05738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *)
  wire _05739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *)
  wire _05740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *)
  wire _05741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *)
  wire _05742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *)
  wire _05743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *)
  wire _05744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *)
  wire _05745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *)
  wire _05746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *)
  wire _05747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *)
  wire _05748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *)
  wire _05749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *)
  wire _05750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *)
  wire _05751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *)
  wire _05752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *)
  wire _05753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *)
  wire _05754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *)
  wire _05755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *)
  wire _05756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *)
  wire _05757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *)
  wire _05758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *)
  wire _05759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *)
  wire _05760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *)
  wire _05761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *)
  wire _05762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *)
  wire _05763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *)
  wire _05764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11898" *)
  wire _05765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11898" *)
  wire _05766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11899" *)
  wire _05767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11899" *)
  wire _05768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11900" *)
  wire _05769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11900" *)
  wire _05770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11901" *)
  wire _05771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11901" *)
  wire _05772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11902" *)
  wire _05773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11902" *)
  wire _05774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11903" *)
  wire _05775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11903" *)
  wire _05776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11904" *)
  wire _05777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11904" *)
  wire _05778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11905" *)
  wire _05779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11905" *)
  wire _05780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11906" *)
  wire _05781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11906" *)
  wire _05782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11907" *)
  wire _05783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11907" *)
  wire _05784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11908" *)
  wire _05785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11908" *)
  wire _05786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11909" *)
  wire _05787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11909" *)
  wire _05788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11910" *)
  wire _05789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11910" *)
  wire _05790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11911" *)
  wire _05791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11911" *)
  wire _05792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11912" *)
  wire _05793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11912" *)
  wire _05794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11913" *)
  wire _05795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11913" *)
  wire _05796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11914" *)
  wire _05797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11914" *)
  wire _05798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11915" *)
  wire _05799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11915" *)
  wire _05800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11916" *)
  wire _05801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11916" *)
  wire _05802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11917" *)
  wire _05803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11917" *)
  wire _05804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11918" *)
  wire _05805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11918" *)
  wire _05806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11919" *)
  wire _05807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11919" *)
  wire _05808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11920" *)
  wire _05809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11920" *)
  wire _05810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11921" *)
  wire _05811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11921" *)
  wire _05812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11922" *)
  wire _05813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11922" *)
  wire _05814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11923" *)
  wire _05815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11923" *)
  wire _05816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11924" *)
  wire _05817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11924" *)
  wire _05818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11925" *)
  wire _05819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11925" *)
  wire _05820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11926" *)
  wire _05821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11926" *)
  wire _05822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11927" *)
  wire _05823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11927" *)
  wire _05824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11928" *)
  wire _05825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11928" *)
  wire _05826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11946" *)
  wire _05827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11946" *)
  wire _05828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11947" *)
  wire _05829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11947" *)
  wire _05830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11948" *)
  wire _05831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11948" *)
  wire _05832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11949" *)
  wire _05833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11949" *)
  wire _05834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11950" *)
  wire _05835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11950" *)
  wire _05836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11951" *)
  wire _05837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11951" *)
  wire _05838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11952" *)
  wire _05839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11952" *)
  wire _05840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11953" *)
  wire _05841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11953" *)
  wire _05842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11954" *)
  wire _05843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11954" *)
  wire _05844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11955" *)
  wire _05845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11955" *)
  wire _05846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11956" *)
  wire _05847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11956" *)
  wire _05848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11957" *)
  wire _05849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11957" *)
  wire _05850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11958" *)
  wire _05851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11958" *)
  wire _05852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11959" *)
  wire _05853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11959" *)
  wire _05854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11960" *)
  wire _05855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11960" *)
  wire _05856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11961" *)
  wire _05857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11961" *)
  wire _05858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11962" *)
  wire _05859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11962" *)
  wire _05860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11963" *)
  wire _05861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11963" *)
  wire _05862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11964" *)
  wire _05863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11964" *)
  wire _05864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11965" *)
  wire _05865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11965" *)
  wire _05866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11966" *)
  wire _05867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11966" *)
  wire _05868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11967" *)
  wire _05869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11967" *)
  wire _05870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11968" *)
  wire _05871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11968" *)
  wire _05872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11969" *)
  wire _05873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11969" *)
  wire _05874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11970" *)
  wire _05875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11970" *)
  wire _05876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11971" *)
  wire _05877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11971" *)
  wire _05878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11972" *)
  wire _05879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11972" *)
  wire _05880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11973" *)
  wire _05881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11973" *)
  wire _05882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11974" *)
  wire _05883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11974" *)
  wire _05884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11975" *)
  wire _05885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11975" *)
  wire _05886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11976" *)
  wire _05887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11976" *)
  wire _05888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11986" *)
  wire _05889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11986" *)
  wire _05890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11987" *)
  wire _05891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11987" *)
  wire _05892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11988" *)
  wire _05893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11988" *)
  wire _05894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11989" *)
  wire _05895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11989" *)
  wire _05896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11990" *)
  wire _05897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11990" *)
  wire _05898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11991" *)
  wire _05899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11991" *)
  wire _05900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11992" *)
  wire _05901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11992" *)
  wire _05902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11993" *)
  wire _05903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11993" *)
  wire _05904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11994" *)
  wire _05905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11994" *)
  wire _05906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11995" *)
  wire _05907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11995" *)
  wire _05908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11996" *)
  wire _05909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11996" *)
  wire _05910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11997" *)
  wire _05911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11997" *)
  wire _05912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11998" *)
  wire _05913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11998" *)
  wire _05914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11999" *)
  wire _05915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11999" *)
  wire _05916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12000" *)
  wire _05917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12000" *)
  wire _05918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12001" *)
  wire _05919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12001" *)
  wire _05920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12002" *)
  wire _05921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12002" *)
  wire _05922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12003" *)
  wire _05923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12003" *)
  wire _05924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12004" *)
  wire _05925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12004" *)
  wire _05926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12005" *)
  wire _05927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12005" *)
  wire _05928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12006" *)
  wire _05929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12006" *)
  wire _05930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12007" *)
  wire _05931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12007" *)
  wire _05932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12008" *)
  wire _05933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12008" *)
  wire _05934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12009" *)
  wire _05935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12009" *)
  wire _05936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12010" *)
  wire _05937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12010" *)
  wire _05938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12011" *)
  wire _05939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12011" *)
  wire _05940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12012" *)
  wire _05941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12012" *)
  wire _05942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12013" *)
  wire _05943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12013" *)
  wire _05944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12014" *)
  wire _05945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12014" *)
  wire _05946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12015" *)
  wire _05947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12015" *)
  wire _05948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12016" *)
  wire _05949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12016" *)
  wire _05950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12034" *)
  wire _05951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12034" *)
  wire _05952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12035" *)
  wire _05953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12035" *)
  wire _05954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12036" *)
  wire _05955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12036" *)
  wire _05956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12037" *)
  wire _05957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12037" *)
  wire _05958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12038" *)
  wire _05959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12038" *)
  wire _05960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12039" *)
  wire _05961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12039" *)
  wire _05962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12040" *)
  wire _05963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12040" *)
  wire _05964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12041" *)
  wire _05965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12041" *)
  wire _05966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12042" *)
  wire _05967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12042" *)
  wire _05968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12043" *)
  wire _05969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12043" *)
  wire _05970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12044" *)
  wire _05971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12044" *)
  wire _05972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12045" *)
  wire _05973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12045" *)
  wire _05974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12046" *)
  wire _05975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12046" *)
  wire _05976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12047" *)
  wire _05977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12047" *)
  wire _05978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12048" *)
  wire _05979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12048" *)
  wire _05980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12049" *)
  wire _05981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12049" *)
  wire _05982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12050" *)
  wire _05983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12050" *)
  wire _05984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12051" *)
  wire _05985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12051" *)
  wire _05986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12052" *)
  wire _05987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12052" *)
  wire _05988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12053" *)
  wire _05989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12053" *)
  wire _05990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12054" *)
  wire _05991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12054" *)
  wire _05992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12055" *)
  wire _05993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12055" *)
  wire _05994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12056" *)
  wire _05995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12056" *)
  wire _05996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12057" *)
  wire _05997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12057" *)
  wire _05998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12058" *)
  wire _05999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12058" *)
  wire _06000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12059" *)
  wire _06001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12059" *)
  wire _06002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12060" *)
  wire _06003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12060" *)
  wire _06004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12061" *)
  wire _06005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12061" *)
  wire _06006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12062" *)
  wire _06007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12062" *)
  wire _06008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12063" *)
  wire _06009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12063" *)
  wire _06010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12064" *)
  wire _06011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12064" *)
  wire _06012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12082" *)
  wire _06013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12082" *)
  wire _06014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12083" *)
  wire _06015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12083" *)
  wire _06016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12084" *)
  wire _06017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12084" *)
  wire _06018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12085" *)
  wire _06019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12085" *)
  wire _06020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12086" *)
  wire _06021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12086" *)
  wire _06022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12087" *)
  wire _06023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12087" *)
  wire _06024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12088" *)
  wire _06025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12088" *)
  wire _06026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12089" *)
  wire _06027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12089" *)
  wire _06028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12090" *)
  wire _06029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12090" *)
  wire _06030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12091" *)
  wire _06031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12091" *)
  wire _06032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12092" *)
  wire _06033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12092" *)
  wire _06034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12093" *)
  wire _06035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12093" *)
  wire _06036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12094" *)
  wire _06037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12094" *)
  wire _06038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12095" *)
  wire _06039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12095" *)
  wire _06040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12096" *)
  wire _06041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12096" *)
  wire _06042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12097" *)
  wire _06043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12097" *)
  wire _06044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12098" *)
  wire _06045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12098" *)
  wire _06046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12099" *)
  wire _06047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12099" *)
  wire _06048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12100" *)
  wire _06049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12100" *)
  wire _06050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12101" *)
  wire _06051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12101" *)
  wire _06052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12102" *)
  wire _06053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12102" *)
  wire _06054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12103" *)
  wire _06055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12103" *)
  wire _06056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12104" *)
  wire _06057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12104" *)
  wire _06058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12105" *)
  wire _06059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12105" *)
  wire _06060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12106" *)
  wire _06061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12106" *)
  wire _06062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12107" *)
  wire _06063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12107" *)
  wire _06064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12108" *)
  wire _06065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12108" *)
  wire _06066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12109" *)
  wire _06067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12109" *)
  wire _06068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12110" *)
  wire _06069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12110" *)
  wire _06070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12111" *)
  wire _06071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12111" *)
  wire _06072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12112" *)
  wire _06073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12112" *)
  wire _06074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12122" *)
  wire _06075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12122" *)
  wire _06076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12123" *)
  wire _06077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12123" *)
  wire _06078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12124" *)
  wire _06079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12124" *)
  wire _06080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12125" *)
  wire _06081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12125" *)
  wire _06082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12126" *)
  wire _06083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12126" *)
  wire _06084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12127" *)
  wire _06085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12127" *)
  wire _06086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12128" *)
  wire _06087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12128" *)
  wire _06088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12129" *)
  wire _06089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12129" *)
  wire _06090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12130" *)
  wire _06091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12130" *)
  wire _06092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12131" *)
  wire _06093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12131" *)
  wire _06094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12132" *)
  wire _06095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12132" *)
  wire _06096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12133" *)
  wire _06097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12133" *)
  wire _06098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12134" *)
  wire _06099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12134" *)
  wire _06100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12135" *)
  wire _06101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12135" *)
  wire _06102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12136" *)
  wire _06103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12136" *)
  wire _06104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12137" *)
  wire _06105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12137" *)
  wire _06106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12138" *)
  wire _06107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12138" *)
  wire _06108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12139" *)
  wire _06109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12139" *)
  wire _06110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12140" *)
  wire _06111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12140" *)
  wire _06112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12141" *)
  wire _06113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12141" *)
  wire _06114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12142" *)
  wire _06115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12142" *)
  wire _06116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12143" *)
  wire _06117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12143" *)
  wire _06118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12144" *)
  wire _06119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12144" *)
  wire _06120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12145" *)
  wire _06121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12145" *)
  wire _06122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12146" *)
  wire _06123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12146" *)
  wire _06124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12147" *)
  wire _06125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12147" *)
  wire _06126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12148" *)
  wire _06127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12148" *)
  wire _06128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12149" *)
  wire _06129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12149" *)
  wire _06130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12150" *)
  wire _06131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12150" *)
  wire _06132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12151" *)
  wire _06133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12151" *)
  wire _06134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12152" *)
  wire _06135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12152" *)
  wire _06136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12162" *)
  wire _06137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12162" *)
  wire _06138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12163" *)
  wire _06139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12163" *)
  wire _06140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12164" *)
  wire _06141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12164" *)
  wire _06142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12165" *)
  wire _06143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12165" *)
  wire _06144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12166" *)
  wire _06145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12166" *)
  wire _06146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12167" *)
  wire _06147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12167" *)
  wire _06148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12168" *)
  wire _06149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12168" *)
  wire _06150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12169" *)
  wire _06151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12169" *)
  wire _06152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12170" *)
  wire _06153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12170" *)
  wire _06154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12171" *)
  wire _06155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12171" *)
  wire _06156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12172" *)
  wire _06157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12172" *)
  wire _06158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12173" *)
  wire _06159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12173" *)
  wire _06160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12174" *)
  wire _06161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12174" *)
  wire _06162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12175" *)
  wire _06163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12175" *)
  wire _06164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12176" *)
  wire _06165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12176" *)
  wire _06166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12177" *)
  wire _06167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12177" *)
  wire _06168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12178" *)
  wire _06169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12178" *)
  wire _06170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12179" *)
  wire _06171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12179" *)
  wire _06172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12180" *)
  wire _06173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12180" *)
  wire _06174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12181" *)
  wire _06175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12181" *)
  wire _06176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12182" *)
  wire _06177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12182" *)
  wire _06178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12183" *)
  wire _06179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12183" *)
  wire _06180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12184" *)
  wire _06181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12184" *)
  wire _06182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12185" *)
  wire _06183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12185" *)
  wire _06184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12186" *)
  wire _06185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12186" *)
  wire _06186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12187" *)
  wire _06187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12187" *)
  wire _06188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12188" *)
  wire _06189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12188" *)
  wire _06190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12189" *)
  wire _06191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12189" *)
  wire _06192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12190" *)
  wire _06193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12190" *)
  wire _06194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12191" *)
  wire _06195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12191" *)
  wire _06196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12192" *)
  wire _06197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12192" *)
  wire _06198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12210" *)
  wire _06199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12210" *)
  wire _06200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12211" *)
  wire _06201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12211" *)
  wire _06202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12212" *)
  wire _06203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12212" *)
  wire _06204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12213" *)
  wire _06205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12213" *)
  wire _06206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12214" *)
  wire _06207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12214" *)
  wire _06208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12215" *)
  wire _06209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12215" *)
  wire _06210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12216" *)
  wire _06211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12216" *)
  wire _06212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12217" *)
  wire _06213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12217" *)
  wire _06214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12218" *)
  wire _06215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12218" *)
  wire _06216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12219" *)
  wire _06217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12219" *)
  wire _06218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12220" *)
  wire _06219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12220" *)
  wire _06220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12221" *)
  wire _06221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12221" *)
  wire _06222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12222" *)
  wire _06223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12222" *)
  wire _06224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12223" *)
  wire _06225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12223" *)
  wire _06226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12224" *)
  wire _06227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12224" *)
  wire _06228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12225" *)
  wire _06229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12225" *)
  wire _06230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12226" *)
  wire _06231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12226" *)
  wire _06232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12227" *)
  wire _06233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12227" *)
  wire _06234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12228" *)
  wire _06235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12228" *)
  wire _06236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12229" *)
  wire _06237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12229" *)
  wire _06238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12230" *)
  wire _06239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12230" *)
  wire _06240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12231" *)
  wire _06241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12231" *)
  wire _06242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12232" *)
  wire _06243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12232" *)
  wire _06244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12233" *)
  wire _06245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12233" *)
  wire _06246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12234" *)
  wire _06247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12234" *)
  wire _06248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12235" *)
  wire _06249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12235" *)
  wire _06250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12236" *)
  wire _06251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12236" *)
  wire _06252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12237" *)
  wire _06253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12237" *)
  wire _06254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12238" *)
  wire _06255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12238" *)
  wire _06256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12239" *)
  wire _06257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12239" *)
  wire _06258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12240" *)
  wire _06259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12240" *)
  wire _06260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12258" *)
  wire _06261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12258" *)
  wire _06262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12259" *)
  wire _06263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12259" *)
  wire _06264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12260" *)
  wire _06265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12260" *)
  wire _06266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12261" *)
  wire _06267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12261" *)
  wire _06268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12262" *)
  wire _06269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12262" *)
  wire _06270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12263" *)
  wire _06271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12263" *)
  wire _06272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12264" *)
  wire _06273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12264" *)
  wire _06274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12265" *)
  wire _06275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12265" *)
  wire _06276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12266" *)
  wire _06277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12266" *)
  wire _06278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12267" *)
  wire _06279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12267" *)
  wire _06280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12268" *)
  wire _06281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12268" *)
  wire _06282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12269" *)
  wire _06283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12269" *)
  wire _06284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12270" *)
  wire _06285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12270" *)
  wire _06286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12271" *)
  wire _06287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12271" *)
  wire _06288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12272" *)
  wire _06289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12272" *)
  wire _06290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12273" *)
  wire _06291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12273" *)
  wire _06292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12274" *)
  wire _06293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12274" *)
  wire _06294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12275" *)
  wire _06295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12275" *)
  wire _06296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12276" *)
  wire _06297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12276" *)
  wire _06298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12277" *)
  wire _06299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12277" *)
  wire _06300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12278" *)
  wire _06301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12278" *)
  wire _06302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12279" *)
  wire _06303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12279" *)
  wire _06304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12280" *)
  wire _06305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12280" *)
  wire _06306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12281" *)
  wire _06307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12281" *)
  wire _06308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12282" *)
  wire _06309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12282" *)
  wire _06310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12283" *)
  wire _06311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12283" *)
  wire _06312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12284" *)
  wire _06313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12284" *)
  wire _06314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12285" *)
  wire _06315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12285" *)
  wire _06316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12286" *)
  wire _06317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12286" *)
  wire _06318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12287" *)
  wire _06319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12287" *)
  wire _06320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12288" *)
  wire _06321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12288" *)
  wire _06322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12298" *)
  wire _06323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12298" *)
  wire _06324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12299" *)
  wire _06325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12299" *)
  wire _06326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12300" *)
  wire _06327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12300" *)
  wire _06328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12301" *)
  wire _06329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12301" *)
  wire _06330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12302" *)
  wire _06331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12302" *)
  wire _06332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12303" *)
  wire _06333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12303" *)
  wire _06334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12304" *)
  wire _06335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12304" *)
  wire _06336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12305" *)
  wire _06337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12305" *)
  wire _06338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12306" *)
  wire _06339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12306" *)
  wire _06340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12307" *)
  wire _06341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12307" *)
  wire _06342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12308" *)
  wire _06343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12308" *)
  wire _06344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12309" *)
  wire _06345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12309" *)
  wire _06346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12310" *)
  wire _06347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12310" *)
  wire _06348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12311" *)
  wire _06349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12311" *)
  wire _06350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12312" *)
  wire _06351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12312" *)
  wire _06352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12313" *)
  wire _06353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12313" *)
  wire _06354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12314" *)
  wire _06355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12314" *)
  wire _06356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12315" *)
  wire _06357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12315" *)
  wire _06358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12316" *)
  wire _06359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12316" *)
  wire _06360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12317" *)
  wire _06361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12317" *)
  wire _06362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12318" *)
  wire _06363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12318" *)
  wire _06364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12319" *)
  wire _06365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12319" *)
  wire _06366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12320" *)
  wire _06367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12320" *)
  wire _06368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12321" *)
  wire _06369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12321" *)
  wire _06370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12322" *)
  wire _06371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12322" *)
  wire _06372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12323" *)
  wire _06373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12323" *)
  wire _06374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12324" *)
  wire _06375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12324" *)
  wire _06376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12325" *)
  wire _06377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12325" *)
  wire _06378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12326" *)
  wire _06379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12326" *)
  wire _06380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12327" *)
  wire _06381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12327" *)
  wire _06382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12328" *)
  wire _06383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12328" *)
  wire _06384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12346" *)
  wire _06385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12346" *)
  wire _06386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12347" *)
  wire _06387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12347" *)
  wire _06388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12348" *)
  wire _06389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12348" *)
  wire _06390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12349" *)
  wire _06391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12349" *)
  wire _06392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12350" *)
  wire _06393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12350" *)
  wire _06394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12351" *)
  wire _06395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12351" *)
  wire _06396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12352" *)
  wire _06397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12352" *)
  wire _06398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12353" *)
  wire _06399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12353" *)
  wire _06400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12354" *)
  wire _06401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12354" *)
  wire _06402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12355" *)
  wire _06403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12355" *)
  wire _06404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12356" *)
  wire _06405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12356" *)
  wire _06406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12357" *)
  wire _06407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12357" *)
  wire _06408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12358" *)
  wire _06409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12358" *)
  wire _06410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12359" *)
  wire _06411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12359" *)
  wire _06412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12360" *)
  wire _06413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12360" *)
  wire _06414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12361" *)
  wire _06415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12361" *)
  wire _06416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12362" *)
  wire _06417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12362" *)
  wire _06418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12363" *)
  wire _06419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12363" *)
  wire _06420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12364" *)
  wire _06421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12364" *)
  wire _06422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12365" *)
  wire _06423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12365" *)
  wire _06424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12366" *)
  wire _06425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12366" *)
  wire _06426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12367" *)
  wire _06427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12367" *)
  wire _06428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12368" *)
  wire _06429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12368" *)
  wire _06430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12369" *)
  wire _06431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12369" *)
  wire _06432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12370" *)
  wire _06433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12370" *)
  wire _06434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12371" *)
  wire _06435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12371" *)
  wire _06436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12372" *)
  wire _06437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12372" *)
  wire _06438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12373" *)
  wire _06439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12373" *)
  wire _06440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12374" *)
  wire _06441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12374" *)
  wire _06442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12375" *)
  wire _06443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12375" *)
  wire _06444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12376" *)
  wire _06445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12376" *)
  wire _06446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12394" *)
  wire _06447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12394" *)
  wire _06448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12395" *)
  wire _06449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12395" *)
  wire _06450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12396" *)
  wire _06451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12396" *)
  wire _06452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12397" *)
  wire _06453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12397" *)
  wire _06454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12398" *)
  wire _06455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12398" *)
  wire _06456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12399" *)
  wire _06457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12399" *)
  wire _06458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12400" *)
  wire _06459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12400" *)
  wire _06460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12401" *)
  wire _06461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12401" *)
  wire _06462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12402" *)
  wire _06463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12402" *)
  wire _06464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12403" *)
  wire _06465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12403" *)
  wire _06466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12404" *)
  wire _06467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12404" *)
  wire _06468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12405" *)
  wire _06469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12405" *)
  wire _06470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12406" *)
  wire _06471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12406" *)
  wire _06472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12407" *)
  wire _06473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12407" *)
  wire _06474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12408" *)
  wire _06475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12408" *)
  wire _06476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12409" *)
  wire _06477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12409" *)
  wire _06478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12410" *)
  wire _06479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12410" *)
  wire _06480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12411" *)
  wire _06481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12411" *)
  wire _06482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12412" *)
  wire _06483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12412" *)
  wire _06484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12413" *)
  wire _06485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12413" *)
  wire _06486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12414" *)
  wire _06487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12414" *)
  wire _06488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12415" *)
  wire _06489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12415" *)
  wire _06490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12416" *)
  wire _06491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12416" *)
  wire _06492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12417" *)
  wire _06493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12417" *)
  wire _06494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12418" *)
  wire _06495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12418" *)
  wire _06496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12419" *)
  wire _06497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12419" *)
  wire _06498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12420" *)
  wire _06499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12420" *)
  wire _06500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12421" *)
  wire _06501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12421" *)
  wire _06502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12422" *)
  wire _06503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12422" *)
  wire _06504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12423" *)
  wire _06505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12423" *)
  wire _06506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12424" *)
  wire _06507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12424" *)
  wire _06508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12434" *)
  wire _06509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12434" *)
  wire _06510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12435" *)
  wire _06511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12435" *)
  wire _06512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12436" *)
  wire _06513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12436" *)
  wire _06514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12437" *)
  wire _06515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12437" *)
  wire _06516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12438" *)
  wire _06517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12438" *)
  wire _06518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12439" *)
  wire _06519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12439" *)
  wire _06520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12440" *)
  wire _06521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12440" *)
  wire _06522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12441" *)
  wire _06523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12441" *)
  wire _06524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12442" *)
  wire _06525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12442" *)
  wire _06526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12443" *)
  wire _06527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12443" *)
  wire _06528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12444" *)
  wire _06529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12444" *)
  wire _06530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12445" *)
  wire _06531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12445" *)
  wire _06532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12446" *)
  wire _06533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12446" *)
  wire _06534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12447" *)
  wire _06535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12447" *)
  wire _06536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12448" *)
  wire _06537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12448" *)
  wire _06538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12449" *)
  wire _06539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12449" *)
  wire _06540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12450" *)
  wire _06541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12450" *)
  wire _06542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12451" *)
  wire _06543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12451" *)
  wire _06544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12452" *)
  wire _06545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12452" *)
  wire _06546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12453" *)
  wire _06547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12453" *)
  wire _06548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12454" *)
  wire _06549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12454" *)
  wire _06550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12455" *)
  wire _06551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12455" *)
  wire _06552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12456" *)
  wire _06553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12456" *)
  wire _06554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12457" *)
  wire _06555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12457" *)
  wire _06556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12458" *)
  wire _06557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12458" *)
  wire _06558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12459" *)
  wire _06559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12459" *)
  wire _06560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12460" *)
  wire _06561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12460" *)
  wire _06562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12461" *)
  wire _06563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12461" *)
  wire _06564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12462" *)
  wire _06565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12462" *)
  wire _06566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12463" *)
  wire _06567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12463" *)
  wire _06568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12464" *)
  wire _06569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12464" *)
  wire _06570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12474" *)
  wire _06571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12474" *)
  wire _06572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12475" *)
  wire _06573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12475" *)
  wire _06574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12476" *)
  wire _06575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12476" *)
  wire _06576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12477" *)
  wire _06577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12477" *)
  wire _06578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12478" *)
  wire _06579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12478" *)
  wire _06580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12479" *)
  wire _06581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12479" *)
  wire _06582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12480" *)
  wire _06583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12480" *)
  wire _06584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12481" *)
  wire _06585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12481" *)
  wire _06586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12482" *)
  wire _06587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12482" *)
  wire _06588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12483" *)
  wire _06589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12483" *)
  wire _06590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12484" *)
  wire _06591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12484" *)
  wire _06592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12485" *)
  wire _06593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12485" *)
  wire _06594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12486" *)
  wire _06595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12486" *)
  wire _06596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12487" *)
  wire _06597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12487" *)
  wire _06598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12488" *)
  wire _06599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12488" *)
  wire _06600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12489" *)
  wire _06601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12489" *)
  wire _06602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12490" *)
  wire _06603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12490" *)
  wire _06604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12491" *)
  wire _06605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12491" *)
  wire _06606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12492" *)
  wire _06607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12492" *)
  wire _06608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12493" *)
  wire _06609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12493" *)
  wire _06610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12494" *)
  wire _06611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12494" *)
  wire _06612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12495" *)
  wire _06613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12495" *)
  wire _06614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12496" *)
  wire _06615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12496" *)
  wire _06616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12497" *)
  wire _06617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12497" *)
  wire _06618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12498" *)
  wire _06619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12498" *)
  wire _06620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12499" *)
  wire _06621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12499" *)
  wire _06622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12500" *)
  wire _06623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12500" *)
  wire _06624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12501" *)
  wire _06625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12501" *)
  wire _06626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12502" *)
  wire _06627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12502" *)
  wire _06628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12503" *)
  wire _06629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12503" *)
  wire _06630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12504" *)
  wire _06631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12504" *)
  wire _06632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12514" *)
  wire _06633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12514" *)
  wire _06634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12515" *)
  wire _06635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12515" *)
  wire _06636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12516" *)
  wire _06637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12516" *)
  wire _06638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12517" *)
  wire _06639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12517" *)
  wire _06640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12518" *)
  wire _06641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12518" *)
  wire _06642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12519" *)
  wire _06643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12519" *)
  wire _06644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12520" *)
  wire _06645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12520" *)
  wire _06646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12521" *)
  wire _06647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12521" *)
  wire _06648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12522" *)
  wire _06649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12522" *)
  wire _06650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12523" *)
  wire _06651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12523" *)
  wire _06652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12524" *)
  wire _06653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12524" *)
  wire _06654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12525" *)
  wire _06655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12525" *)
  wire _06656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12526" *)
  wire _06657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12526" *)
  wire _06658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12527" *)
  wire _06659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12527" *)
  wire _06660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12528" *)
  wire _06661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12528" *)
  wire _06662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12529" *)
  wire _06663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12529" *)
  wire _06664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12530" *)
  wire _06665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12530" *)
  wire _06666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12531" *)
  wire _06667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12531" *)
  wire _06668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12532" *)
  wire _06669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12532" *)
  wire _06670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12533" *)
  wire _06671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12533" *)
  wire _06672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12534" *)
  wire _06673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12534" *)
  wire _06674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12535" *)
  wire _06675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12535" *)
  wire _06676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12536" *)
  wire _06677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12536" *)
  wire _06678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12537" *)
  wire _06679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12537" *)
  wire _06680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12538" *)
  wire _06681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12538" *)
  wire _06682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12539" *)
  wire _06683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12539" *)
  wire _06684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12540" *)
  wire _06685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12540" *)
  wire _06686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12541" *)
  wire _06687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12541" *)
  wire _06688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12542" *)
  wire _06689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12542" *)
  wire _06690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12543" *)
  wire _06691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12543" *)
  wire _06692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12544" *)
  wire _06693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12544" *)
  wire _06694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12554" *)
  wire _06695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12554" *)
  wire _06696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12555" *)
  wire _06697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12555" *)
  wire _06698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12556" *)
  wire _06699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12556" *)
  wire _06700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12557" *)
  wire _06701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12557" *)
  wire _06702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12558" *)
  wire _06703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12558" *)
  wire _06704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12559" *)
  wire _06705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12559" *)
  wire _06706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12560" *)
  wire _06707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12560" *)
  wire _06708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12561" *)
  wire _06709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12561" *)
  wire _06710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12562" *)
  wire _06711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12562" *)
  wire _06712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12563" *)
  wire _06713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12563" *)
  wire _06714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12564" *)
  wire _06715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12564" *)
  wire _06716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12565" *)
  wire _06717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12565" *)
  wire _06718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12566" *)
  wire _06719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12566" *)
  wire _06720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12567" *)
  wire _06721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12567" *)
  wire _06722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12568" *)
  wire _06723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12568" *)
  wire _06724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12569" *)
  wire _06725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12569" *)
  wire _06726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12570" *)
  wire _06727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12570" *)
  wire _06728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12571" *)
  wire _06729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12571" *)
  wire _06730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12572" *)
  wire _06731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12572" *)
  wire _06732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12573" *)
  wire _06733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12573" *)
  wire _06734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12574" *)
  wire _06735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12574" *)
  wire _06736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12575" *)
  wire _06737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12575" *)
  wire _06738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12576" *)
  wire _06739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12576" *)
  wire _06740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12577" *)
  wire _06741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12577" *)
  wire _06742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12578" *)
  wire _06743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12578" *)
  wire _06744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12579" *)
  wire _06745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12579" *)
  wire _06746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12580" *)
  wire _06747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12580" *)
  wire _06748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12581" *)
  wire _06749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12581" *)
  wire _06750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12582" *)
  wire _06751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12582" *)
  wire _06752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12583" *)
  wire _06753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12583" *)
  wire _06754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12584" *)
  wire _06755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12584" *)
  wire _06756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12594" *)
  wire _06757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12594" *)
  wire _06758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12595" *)
  wire _06759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12595" *)
  wire _06760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12596" *)
  wire _06761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12596" *)
  wire _06762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12597" *)
  wire _06763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12597" *)
  wire _06764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12598" *)
  wire _06765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12598" *)
  wire _06766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12599" *)
  wire _06767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12599" *)
  wire _06768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12600" *)
  wire _06769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12600" *)
  wire _06770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12601" *)
  wire _06771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12601" *)
  wire _06772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12602" *)
  wire _06773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12602" *)
  wire _06774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12603" *)
  wire _06775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12603" *)
  wire _06776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12604" *)
  wire _06777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12604" *)
  wire _06778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12605" *)
  wire _06779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12605" *)
  wire _06780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12606" *)
  wire _06781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12606" *)
  wire _06782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12607" *)
  wire _06783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12607" *)
  wire _06784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12608" *)
  wire _06785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12608" *)
  wire _06786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12615" *)
  wire _06787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12622" *)
  wire _06788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12622" *)
  wire _06789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12623" *)
  wire _06790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12623" *)
  wire _06791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12624" *)
  wire _06792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12624" *)
  wire _06793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12625" *)
  wire _06794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12625" *)
  wire _06795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12626" *)
  wire _06796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12626" *)
  wire _06797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12627" *)
  wire _06798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12627" *)
  wire _06799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12628" *)
  wire _06800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12628" *)
  wire _06801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12629" *)
  wire _06802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12629" *)
  wire _06803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12630" *)
  wire _06804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12630" *)
  wire _06805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12631" *)
  wire _06806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12631" *)
  wire _06807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12632" *)
  wire _06808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12632" *)
  wire _06809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12633" *)
  wire _06810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12633" *)
  wire _06811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12634" *)
  wire _06812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12634" *)
  wire _06813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12635" *)
  wire _06814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12635" *)
  wire _06815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12636" *)
  wire _06816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12636" *)
  wire _06817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12643" *)
  wire _06818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12650" *)
  wire _06819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12650" *)
  wire _06820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12651" *)
  wire _06821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12651" *)
  wire _06822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12652" *)
  wire _06823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12652" *)
  wire _06824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12653" *)
  wire _06825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12653" *)
  wire _06826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12654" *)
  wire _06827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12654" *)
  wire _06828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12655" *)
  wire _06829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12655" *)
  wire _06830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12656" *)
  wire _06831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12656" *)
  wire _06832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12657" *)
  wire _06833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12657" *)
  wire _06834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12658" *)
  wire _06835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12658" *)
  wire _06836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12659" *)
  wire _06837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12659" *)
  wire _06838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12660" *)
  wire _06839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12660" *)
  wire _06840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12661" *)
  wire _06841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12661" *)
  wire _06842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12662" *)
  wire _06843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12662" *)
  wire _06844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12663" *)
  wire _06845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12663" *)
  wire _06846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12664" *)
  wire _06847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12664" *)
  wire _06848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12671" *)
  wire _06849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12678" *)
  wire _06850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12678" *)
  wire _06851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12679" *)
  wire _06852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12679" *)
  wire _06853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12680" *)
  wire _06854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12680" *)
  wire _06855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12681" *)
  wire _06856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12681" *)
  wire _06857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12682" *)
  wire _06858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12682" *)
  wire _06859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12683" *)
  wire _06860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12683" *)
  wire _06861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12684" *)
  wire _06862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12684" *)
  wire _06863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12685" *)
  wire _06864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12685" *)
  wire _06865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12686" *)
  wire _06866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12686" *)
  wire _06867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12687" *)
  wire _06868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12687" *)
  wire _06869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12688" *)
  wire _06870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12688" *)
  wire _06871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12689" *)
  wire _06872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12689" *)
  wire _06873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12690" *)
  wire _06874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12690" *)
  wire _06875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12691" *)
  wire _06876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12691" *)
  wire _06877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12692" *)
  wire _06878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12692" *)
  wire _06879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12699" *)
  wire _06880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12706" *)
  wire _06881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12706" *)
  wire _06882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12707" *)
  wire _06883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12707" *)
  wire _06884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12708" *)
  wire _06885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12708" *)
  wire _06886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12709" *)
  wire _06887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12709" *)
  wire _06888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12710" *)
  wire _06889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12710" *)
  wire _06890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12711" *)
  wire _06891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12711" *)
  wire _06892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12712" *)
  wire _06893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12712" *)
  wire _06894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12713" *)
  wire _06895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12713" *)
  wire _06896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12714" *)
  wire _06897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12714" *)
  wire _06898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12715" *)
  wire _06899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12715" *)
  wire _06900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12716" *)
  wire _06901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12716" *)
  wire _06902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12717" *)
  wire _06903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12717" *)
  wire _06904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12718" *)
  wire _06905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12718" *)
  wire _06906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12719" *)
  wire _06907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12719" *)
  wire _06908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12720" *)
  wire _06909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12720" *)
  wire _06910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12727" *)
  wire _06911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12734" *)
  wire _06912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12734" *)
  wire _06913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12735" *)
  wire _06914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12735" *)
  wire _06915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12736" *)
  wire _06916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12736" *)
  wire _06917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12737" *)
  wire _06918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12737" *)
  wire _06919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12738" *)
  wire _06920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12738" *)
  wire _06921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12739" *)
  wire _06922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12739" *)
  wire _06923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12740" *)
  wire _06924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12740" *)
  wire _06925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12741" *)
  wire _06926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12741" *)
  wire _06927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12742" *)
  wire _06928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12742" *)
  wire _06929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12743" *)
  wire _06930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12743" *)
  wire _06931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12744" *)
  wire _06932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12744" *)
  wire _06933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12745" *)
  wire _06934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12745" *)
  wire _06935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12746" *)
  wire _06936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12746" *)
  wire _06937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12747" *)
  wire _06938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12747" *)
  wire _06939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12748" *)
  wire _06940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12748" *)
  wire _06941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12755" *)
  wire _06942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12762" *)
  wire _06943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12762" *)
  wire _06944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12763" *)
  wire _06945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12763" *)
  wire _06946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12764" *)
  wire _06947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12764" *)
  wire _06948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12765" *)
  wire _06949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12765" *)
  wire _06950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12766" *)
  wire _06951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12766" *)
  wire _06952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12767" *)
  wire _06953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12767" *)
  wire _06954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12768" *)
  wire _06955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12768" *)
  wire _06956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12769" *)
  wire _06957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12769" *)
  wire _06958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12770" *)
  wire _06959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12770" *)
  wire _06960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12771" *)
  wire _06961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12771" *)
  wire _06962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12772" *)
  wire _06963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12772" *)
  wire _06964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12773" *)
  wire _06965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12773" *)
  wire _06966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12774" *)
  wire _06967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12774" *)
  wire _06968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12775" *)
  wire _06969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12775" *)
  wire _06970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12776" *)
  wire _06971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12776" *)
  wire _06972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12783" *)
  wire _06973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12790" *)
  wire _06974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12790" *)
  wire _06975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12791" *)
  wire _06976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12791" *)
  wire _06977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12792" *)
  wire _06978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12792" *)
  wire _06979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12793" *)
  wire _06980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12793" *)
  wire _06981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12794" *)
  wire _06982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12794" *)
  wire _06983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12795" *)
  wire _06984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12795" *)
  wire _06985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12796" *)
  wire _06986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12796" *)
  wire _06987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12797" *)
  wire _06988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12797" *)
  wire _06989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12798" *)
  wire _06990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12798" *)
  wire _06991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12799" *)
  wire _06992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12799" *)
  wire _06993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12800" *)
  wire _06994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12800" *)
  wire _06995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12801" *)
  wire _06996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12801" *)
  wire _06997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12802" *)
  wire _06998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12802" *)
  wire _06999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12803" *)
  wire _07000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12803" *)
  wire _07001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12804" *)
  wire _07002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12804" *)
  wire _07003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12811" *)
  wire _07004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12818" *)
  wire _07005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12818" *)
  wire _07006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12819" *)
  wire _07007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12819" *)
  wire _07008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12820" *)
  wire _07009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12820" *)
  wire _07010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12821" *)
  wire _07011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12821" *)
  wire _07012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12822" *)
  wire _07013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12822" *)
  wire _07014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12823" *)
  wire _07015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12823" *)
  wire _07016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12824" *)
  wire _07017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12824" *)
  wire _07018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12825" *)
  wire _07019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12825" *)
  wire _07020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12826" *)
  wire _07021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12826" *)
  wire _07022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12827" *)
  wire _07023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12827" *)
  wire _07024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12828" *)
  wire _07025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12828" *)
  wire _07026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12829" *)
  wire _07027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12829" *)
  wire _07028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12830" *)
  wire _07029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12830" *)
  wire _07030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12831" *)
  wire _07031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12831" *)
  wire _07032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12832" *)
  wire _07033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12832" *)
  wire _07034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12839" *)
  wire _07035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12846" *)
  wire _07036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12846" *)
  wire _07037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12847" *)
  wire _07038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12847" *)
  wire _07039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12848" *)
  wire _07040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12848" *)
  wire _07041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12849" *)
  wire _07042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12849" *)
  wire _07043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12850" *)
  wire _07044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12850" *)
  wire _07045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12851" *)
  wire _07046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12851" *)
  wire _07047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12852" *)
  wire _07048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12852" *)
  wire _07049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12853" *)
  wire _07050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12853" *)
  wire _07051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12854" *)
  wire _07052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12854" *)
  wire _07053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12855" *)
  wire _07054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12855" *)
  wire _07055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12856" *)
  wire _07056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12856" *)
  wire _07057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12857" *)
  wire _07058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12857" *)
  wire _07059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12858" *)
  wire _07060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12858" *)
  wire _07061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12859" *)
  wire _07062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12859" *)
  wire _07063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12860" *)
  wire _07064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12860" *)
  wire _07065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12867" *)
  wire _07066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12874" *)
  wire _07067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12874" *)
  wire _07068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12875" *)
  wire _07069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12875" *)
  wire _07070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12876" *)
  wire _07071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12876" *)
  wire _07072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12877" *)
  wire _07073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12877" *)
  wire _07074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12878" *)
  wire _07075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12878" *)
  wire _07076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12879" *)
  wire _07077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12879" *)
  wire _07078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12880" *)
  wire _07079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12880" *)
  wire _07080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12881" *)
  wire _07081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12881" *)
  wire _07082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12882" *)
  wire _07083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12882" *)
  wire _07084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12883" *)
  wire _07085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12883" *)
  wire _07086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12884" *)
  wire _07087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12884" *)
  wire _07088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12885" *)
  wire _07089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12885" *)
  wire _07090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12886" *)
  wire _07091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12886" *)
  wire _07092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12887" *)
  wire _07093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12887" *)
  wire _07094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12888" *)
  wire _07095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12888" *)
  wire _07096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12895" *)
  wire _07097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12902" *)
  wire _07098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12902" *)
  wire _07099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12903" *)
  wire _07100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12903" *)
  wire _07101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12904" *)
  wire _07102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12904" *)
  wire _07103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12905" *)
  wire _07104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12905" *)
  wire _07105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12906" *)
  wire _07106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12906" *)
  wire _07107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12907" *)
  wire _07108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12907" *)
  wire _07109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12908" *)
  wire _07110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12908" *)
  wire _07111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12909" *)
  wire _07112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12909" *)
  wire _07113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12910" *)
  wire _07114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12910" *)
  wire _07115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12911" *)
  wire _07116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12911" *)
  wire _07117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12912" *)
  wire _07118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12912" *)
  wire _07119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12913" *)
  wire _07120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12913" *)
  wire _07121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12914" *)
  wire _07122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12914" *)
  wire _07123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12915" *)
  wire _07124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12915" *)
  wire _07125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12916" *)
  wire _07126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12916" *)
  wire _07127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12923" *)
  wire _07128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12930" *)
  wire _07129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12930" *)
  wire _07130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12931" *)
  wire _07131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12931" *)
  wire _07132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12932" *)
  wire _07133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12932" *)
  wire _07134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12933" *)
  wire _07135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12933" *)
  wire _07136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12934" *)
  wire _07137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12934" *)
  wire _07138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12935" *)
  wire _07139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12935" *)
  wire _07140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12936" *)
  wire _07141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12936" *)
  wire _07142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12937" *)
  wire _07143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12937" *)
  wire _07144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12938" *)
  wire _07145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12938" *)
  wire _07146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12939" *)
  wire _07147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12939" *)
  wire _07148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12940" *)
  wire _07149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12940" *)
  wire _07150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12941" *)
  wire _07151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12941" *)
  wire _07152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12942" *)
  wire _07153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12942" *)
  wire _07154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12943" *)
  wire _07155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12943" *)
  wire _07156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12944" *)
  wire _07157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12944" *)
  wire _07158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12951" *)
  wire _07159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12958" *)
  wire _07160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12958" *)
  wire _07161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12959" *)
  wire _07162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12959" *)
  wire _07163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12960" *)
  wire _07164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12960" *)
  wire _07165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12961" *)
  wire _07166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12961" *)
  wire _07167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12962" *)
  wire _07168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12962" *)
  wire _07169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12963" *)
  wire _07170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12963" *)
  wire _07171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12964" *)
  wire _07172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12964" *)
  wire _07173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12965" *)
  wire _07174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12965" *)
  wire _07175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12966" *)
  wire _07176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12966" *)
  wire _07177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12967" *)
  wire _07178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12967" *)
  wire _07179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12968" *)
  wire _07180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12968" *)
  wire _07181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12969" *)
  wire _07182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12969" *)
  wire _07183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12970" *)
  wire _07184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12970" *)
  wire _07185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12971" *)
  wire _07186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12971" *)
  wire _07187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12972" *)
  wire _07188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12972" *)
  wire _07189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12979" *)
  wire _07190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12986" *)
  wire _07191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12986" *)
  wire _07192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12987" *)
  wire _07193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12987" *)
  wire _07194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12988" *)
  wire _07195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12988" *)
  wire _07196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12989" *)
  wire _07197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12989" *)
  wire _07198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12990" *)
  wire _07199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12990" *)
  wire _07200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12991" *)
  wire _07201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12991" *)
  wire _07202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12992" *)
  wire _07203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12992" *)
  wire _07204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12993" *)
  wire _07205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12993" *)
  wire _07206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12994" *)
  wire _07207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12994" *)
  wire _07208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12995" *)
  wire _07209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12995" *)
  wire _07210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12996" *)
  wire _07211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12996" *)
  wire _07212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12997" *)
  wire _07213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12997" *)
  wire _07214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12998" *)
  wire _07215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12998" *)
  wire _07216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12999" *)
  wire _07217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12999" *)
  wire _07218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13000" *)
  wire _07219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13000" *)
  wire _07220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13007" *)
  wire _07221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13014" *)
  wire _07222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13014" *)
  wire _07223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13015" *)
  wire _07224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13015" *)
  wire _07225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13016" *)
  wire _07226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13016" *)
  wire _07227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13017" *)
  wire _07228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13017" *)
  wire _07229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13018" *)
  wire _07230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13018" *)
  wire _07231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13019" *)
  wire _07232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13019" *)
  wire _07233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13020" *)
  wire _07234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13020" *)
  wire _07235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13021" *)
  wire _07236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13021" *)
  wire _07237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13022" *)
  wire _07238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13022" *)
  wire _07239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13023" *)
  wire _07240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13023" *)
  wire _07241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13024" *)
  wire _07242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13024" *)
  wire _07243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13025" *)
  wire _07244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13025" *)
  wire _07245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13026" *)
  wire _07246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13026" *)
  wire _07247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13027" *)
  wire _07248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13027" *)
  wire _07249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13028" *)
  wire _07250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13028" *)
  wire _07251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13035" *)
  wire _07252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13047" *)
  wire _07253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13047" *)
  wire _07254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13048" *)
  wire _07255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13048" *)
  wire _07256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13048" *)
  wire _07257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13056" *)
  wire _07258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13056" *)
  wire _07259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13057" *)
  wire _07260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13057" *)
  wire _07261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13057" *)
  wire _07262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13065" *)
  wire _07263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13065" *)
  wire _07264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13066" *)
  wire _07265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13066" *)
  wire _07266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13066" *)
  wire _07267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13074" *)
  wire _07268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13074" *)
  wire _07269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13075" *)
  wire _07270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13075" *)
  wire _07271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13075" *)
  wire _07272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13083" *)
  wire _07273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13083" *)
  wire _07274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13084" *)
  wire _07275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13084" *)
  wire _07276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13084" *)
  wire _07277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13092" *)
  wire _07278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13092" *)
  wire _07279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13093" *)
  wire _07280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13093" *)
  wire _07281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13093" *)
  wire _07282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13101" *)
  wire _07283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13101" *)
  wire _07284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13102" *)
  wire _07285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13102" *)
  wire _07286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13102" *)
  wire _07287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13110" *)
  wire _07288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13110" *)
  wire _07289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13111" *)
  wire _07290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13111" *)
  wire _07291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13111" *)
  wire _07292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13119" *)
  wire _07293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13119" *)
  wire _07294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13120" *)
  wire _07295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13120" *)
  wire _07296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13120" *)
  wire _07297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13128" *)
  wire _07298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13128" *)
  wire _07299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13129" *)
  wire _07300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13129" *)
  wire _07301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13129" *)
  wire _07302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13137" *)
  wire _07303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13137" *)
  wire _07304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13138" *)
  wire _07305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13138" *)
  wire _07306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13138" *)
  wire _07307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13146" *)
  wire _07308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13146" *)
  wire _07309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13147" *)
  wire _07310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13147" *)
  wire _07311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13147" *)
  wire _07312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13155" *)
  wire _07313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13155" *)
  wire _07314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13156" *)
  wire _07315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13156" *)
  wire _07316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13156" *)
  wire _07317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13164" *)
  wire _07318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13164" *)
  wire _07319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13165" *)
  wire _07320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13165" *)
  wire _07321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13165" *)
  wire _07322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13173" *)
  wire _07323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13173" *)
  wire _07324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13174" *)
  wire _07325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13174" *)
  wire _07326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13174" *)
  wire _07327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13182" *)
  wire _07328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13182" *)
  wire _07329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13183" *)
  wire _07330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13183" *)
  wire _07331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13183" *)
  wire _07332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13193" *)
  wire _07333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13207" *)
  wire _07334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13214" *)
  wire _07335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13214" *)
  wire _07336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13225" *)
  wire _07337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13238" *)
  wire _07338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13252" *)
  wire _07339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13266" *)
  wire _07340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13280" *)
  wire _07341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13294" *)
  wire _07342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13308" *)
  wire _07343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13322" *)
  wire _07344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13336" *)
  wire _07345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13350" *)
  wire _07346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13364" *)
  wire _07347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13373" *)
  wire _07348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13387" *)
  wire _07349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13401" *)
  wire _07350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13528" *)
  wire _07351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13530" *)
  wire _07352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13530" *)
  wire _07353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13544" *)
  wire _07354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13546" *)
  wire _07355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13546" *)
  wire _07356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13560" *)
  wire _07357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13562" *)
  wire _07358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13562" *)
  wire _07359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13576" *)
  wire _07360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13578" *)
  wire _07361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13578" *)
  wire _07362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13592" *)
  wire _07363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13594" *)
  wire _07364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13594" *)
  wire _07365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13608" *)
  wire _07366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13610" *)
  wire _07367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13610" *)
  wire _07368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13624" *)
  wire _07369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13626" *)
  wire _07370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13626" *)
  wire _07371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13640" *)
  wire _07372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13642" *)
  wire _07373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13642" *)
  wire _07374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13656" *)
  wire _07375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13658" *)
  wire _07376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13658" *)
  wire _07377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13672" *)
  wire _07378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13674" *)
  wire _07379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13674" *)
  wire _07380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13688" *)
  wire _07381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13690" *)
  wire _07382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13690" *)
  wire _07383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13704" *)
  wire _07384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13706" *)
  wire _07385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13706" *)
  wire _07386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13720" *)
  wire _07387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13722" *)
  wire _07388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13722" *)
  wire _07389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13736" *)
  wire _07390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13738" *)
  wire _07391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13738" *)
  wire _07392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13752" *)
  wire _07393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13754" *)
  wire _07394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13754" *)
  wire _07395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13768" *)
  wire _07396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13770" *)
  wire _07397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13770" *)
  wire _07398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13976" *)
  wire _07399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13978" *)
  wire _07400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13980" *)
  wire _07401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13982" *)
  wire _07402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13984" *)
  wire _07403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13986" *)
  wire _07404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13988" *)
  wire _07405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13990" *)
  wire _07406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13992" *)
  wire _07407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13994" *)
  wire _07408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13996" *)
  wire _07409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13998" *)
  wire _07410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14000" *)
  wire _07411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14002" *)
  wire _07412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14004" *)
  wire _07413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14006" *)
  wire _07414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14071" *)
  wire _07415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14071" *)
  wire _07416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14110" *)
  wire _07417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14113" *)
  wire _07418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14113" *)
  wire _07419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14121" *)
  wire _07420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14125" *)
  wire _07421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14131" *)
  wire _07422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14134" *)
  wire _07423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14136" *)
  wire _07424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14139" *)
  wire _07425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14143" *)
  wire _07426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14151" *)
  wire _07427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14153" *)
  wire _07428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14157" *)
  wire _07429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14159" *)
  wire _07430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14162" *)
  wire _07431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14164" *)
  wire _07432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14167" *)
  wire _07433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14167" *)
  wire _07434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14171" *)
  wire _07435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14184" *)
  wire _07436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14186" *)
  wire _07437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *)
  wire _07438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *)
  wire _07439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14190" *)
  wire _07440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14191" *)
  wire _07441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14191" *)
  wire _07442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14195" *)
  wire _07443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14197" *)
  wire _07444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14204" *)
  wire _07445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14204" *)
  wire _07446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14206" *)
  wire _07447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14212" *)
  wire _07448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14225" *)
  wire _07449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14226" *)
  wire _07450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14226" *)
  wire _07451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14227" *)
  wire _07452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14227" *)
  wire _07453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14229" *)
  wire _07454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14234" *)
  wire _07455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14236" *)
  wire _07456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14239" *)
  wire _07457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14242" *)
  wire _07458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14242" *)
  wire _07459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14252" *)
  wire _07460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14254" *)
  wire _07461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14258" *)
  wire _07462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14258" *)
  wire _07463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14267" *)
  wire _07464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14269" *)
  wire _07465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14273" *)
  wire _07466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14276" *)
  wire _07467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14276" *)
  wire _07468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14278" *)
  wire _07469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14284" *)
  wire _07470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14286" *)
  wire _07471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14288" *)
  wire _07472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14290" *)
  wire _07473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14293" *)
  wire _07474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14295" *)
  wire _07475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14299" *)
  wire _07476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14303" *)
  wire _07477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14305" *)
  wire _07478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14305" *)
  wire _07479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14309" *)
  wire _07480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14309" *)
  wire _07481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14320" *)
  wire _07482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14322" *)
  wire _07483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14323" *)
  wire _07484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14323" *)
  wire _07485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14326" *)
  wire _07486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14326" *)
  wire _07487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14337" *)
  wire _07488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14340" *)
  wire _07489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14343" *)
  wire _07490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14343" *)
  wire _07491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14347" *)
  wire _07492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14349" *)
  wire _07493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14354" *)
  wire _07494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14356" *)
  wire _07495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14358" *)
  wire _07496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14361" *)
  wire _07497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14363" *)
  wire _07498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14363" *)
  wire _07499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14368" *)
  wire _07500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14370" *)
  wire _07501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14374" *)
  wire _07502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14376" *)
  wire _07503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14378" *)
  wire _07504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14382" *)
  wire _07505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14384" *)
  wire _07506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14387" *)
  wire _07507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14390" *)
  wire _07508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14392" *)
  wire _07509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14397" *)
  wire _07510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14399" *)
  wire _07511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14401" *)
  wire _07512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14404" *)
  wire _07513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14407" *)
  wire _07514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14409" *)
  wire _07515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14413" *)
  wire _07516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14415" *)
  wire _07517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14417" *)
  wire _07518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14419" *)
  wire _07519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14423" *)
  wire _07520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14425" *)
  wire _07521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14427" *)
  wire _07522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14430" *)
  wire _07523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14433" *)
  wire _07524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14435" *)
  wire _07525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14437" *)
  wire _07526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14441" *)
  wire _07527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14443" *)
  wire _07528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14445" *)
  wire _07529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14447" *)
  wire _07530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14449" *)
  wire _07531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14453" *)
  wire _07532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14455" *)
  wire _07533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14457" *)
  wire _07534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14459" *)
  wire _07535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14462" *)
  wire _07536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14465" *)
  wire _07537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14467" *)
  wire _07538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14469" *)
  wire _07539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14471" *)
  wire _07540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14485" *)
  wire _07541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14488" *)
  wire _07542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14490" *)
  wire _07543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14498" *)
  wire _07544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14500" *)
  wire _07545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14501" *)
  wire _07546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14502" *)
  wire _07547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14505" *)
  wire _07548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14507" *)
  wire _07549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14509" *)
  wire _07550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14509" *)
  wire _07551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14522" *)
  wire _07552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14527" *)
  wire _07553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14528" *)
  wire _07554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14534" *)
  wire _07555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14535" *)
  wire _07556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14535" *)
  wire _07557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14540" *)
  wire _07558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14542" *)
  wire _07559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14542" *)
  wire _07560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14557" *)
  wire _07561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14559" *)
  wire _07562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14564" *)
  wire _07563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14566" *)
  wire _07564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14568" *)
  wire _07565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14608" *)
  wire _07566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14612" *)
  wire _07567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14614" *)
  wire _07568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14615" *)
  wire _07569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14624" *)
  wire _07570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14633" *)
  wire _07571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14633" *)
  wire _07572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14633" *)
  wire _07573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14636" *)
  wire _07574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14636" *)
  wire _07575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14636" *)
  wire _07576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14639" *)
  wire _07577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14639" *)
  wire _07578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14639" *)
  wire _07579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14642" *)
  wire _07580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14642" *)
  wire _07581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14642" *)
  wire _07582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14645" *)
  wire _07583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14645" *)
  wire _07584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14645" *)
  wire _07585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14648" *)
  wire _07586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14648" *)
  wire _07587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14648" *)
  wire _07588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14651" *)
  wire _07589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14651" *)
  wire _07590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14651" *)
  wire _07591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14654" *)
  wire _07592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14654" *)
  wire _07593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14654" *)
  wire _07594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14659" *)
  wire _07595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14659" *)
  wire _07596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14662" *)
  wire _07597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14662" *)
  wire _07598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14662" *)
  wire _07599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14665" *)
  wire _07600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14665" *)
  wire _07601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14665" *)
  wire _07602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14668" *)
  wire _07603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14668" *)
  wire _07604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14668" *)
  wire _07605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14671" *)
  wire _07606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14671" *)
  wire _07607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14671" *)
  wire _07608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14674" *)
  wire _07609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14674" *)
  wire _07610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14674" *)
  wire _07611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14698" *)
  wire _07612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14724" *)
  wire _07613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14733" *)
  wire _07614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14746" *)
  wire _07615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14754" *)
  wire _07616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14764" *)
  wire _07617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14777" *)
  wire _07618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14781" *)
  wire _07619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14783" *)
  wire _07620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14785" *)
  wire _07621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14786" *)
  wire _07622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14789" *)
  wire _07623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14791" *)
  wire _07624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14793" *)
  wire _07625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14795" *)
  wire _07626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14797" *)
  wire _07627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14799" *)
  wire _07628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14801" *)
  wire _07629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14803" *)
  wire _07630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14805" *)
  wire _07631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14807" *)
  wire _07632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14809" *)
  wire _07633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14811" *)
  wire _07634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14813" *)
  wire _07635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14815" *)
  wire _07636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14817" *)
  wire _07637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14819" *)
  wire _07638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14828" *)
  wire _07639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14832" *)
  wire _07640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14835" *)
  wire _07641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14841" *)
  wire _07642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14850" *)
  wire _07643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14860" *)
  wire _07644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14860" *)
  wire _07645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14879" *)
  wire _07646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14884" *)
  wire _07647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14884" *)
  wire _07648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14969" *)
  wire _07649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14970" *)
  wire _07650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *)
  wire _07651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *)
  wire _07652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *)
  wire _07653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14983" *)
  wire _07654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *)
  wire _07655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *)
  wire _07656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *)
  wire _07657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14985" *)
  wire _07658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14989" *)
  wire _07659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14990" *)
  wire _07660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14999" *)
  wire _07661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15003" *)
  wire _07662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15009" *)
  wire _07663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15015" *)
  wire _07664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15020" *)
  wire _07665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15027" *)
  wire _07666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15032" *)
  wire _07667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15041" *)
  wire _07668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15045" *)
  wire _07669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15051" *)
  wire _07670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15369" *)
  wire _07671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15369" *)
  wire _07672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15383" *)
  wire _07673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15383" *)
  wire _07674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15396" *)
  wire _07675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15396" *)
  wire _07676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15410" *)
  wire _07677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15410" *)
  wire _07678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15424" *)
  wire _07679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15424" *)
  wire _07680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15438" *)
  wire _07681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15438" *)
  wire _07682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15452" *)
  wire _07683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15452" *)
  wire _07684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15466" *)
  wire _07685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15466" *)
  wire _07686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15480" *)
  wire _07687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15480" *)
  wire _07688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15514" *)
  wire _07689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15514" *)
  wire _07690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15621" *)
  wire _07691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15629" *)
  wire _07692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16448" *)
  wire _07693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16448" *)
  wire _07694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16522" *)
  wire _07695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *)
  wire _07696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *)
  wire _07697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *)
  wire _07698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *)
  wire _07699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *)
  wire _07700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *)
  wire _07701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *)
  wire _07702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *)
  wire _07703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *)
  wire _07704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *)
  wire _07705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *)
  wire _07706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *)
  wire _07707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *)
  wire _07708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16717" *)
  wire _07709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16736" *)
  wire _07710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16759" *)
  wire _07711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16770" *)
  wire _07712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16781" *)
  wire _07713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16800" *)
  wire _07714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16831" *)
  wire _07715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16842" *)
  wire _07716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16853" *)
  wire _07717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16876" *)
  wire _07718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16887" *)
  wire _07719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16898" *)
  wire _07720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16909" *)
  wire _07721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16920" *)
  wire _07722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16931" *)
  wire _07723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16950" *)
  wire _07724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *)
  wire _07725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17257" *)
  wire _07726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *)
  wire _07727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *)
  wire _07728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *)
  wire _07729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17443" *)
  wire _07730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *)
  wire _07731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *)
  wire _07732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *)
  wire _07733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *)
  wire _07734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *)
  wire _07735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17782" *)
  wire _07736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *)
  wire _07737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17838" *)
  wire _07738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *)
  wire _07739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17894" *)
  wire _07740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *)
  wire _07741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17954" *)
  wire _07742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18029" *)
  wire _07743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18029" *)
  wire _07744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18136" *)
  wire _07745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18136" *)
  wire _07746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *)
  wire _07747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *)
  wire _07748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18186" *)
  wire _07749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18186" *)
  wire _07750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18283" *)
  wire _07751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18283" *)
  wire _07752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18305" *)
  wire _07753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18305" *)
  wire _07754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18349" *)
  wire _07755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18349" *)
  wire _07756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18369" *)
  wire _07757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18381" *)
  wire _07758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18381" *)
  wire _07759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18425" *)
  wire _07760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18425" *)
  wire _07761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18473" *)
  wire _07762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18473" *)
  wire _07763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18486" *)
  wire _07764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18494" *)
  wire _07765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18494" *)
  wire _07766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18512" *)
  wire _07767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18512" *)
  wire _07768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18544" *)
  wire _07769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18544" *)
  wire _07770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18575" *)
  wire _07771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18592" *)
  wire _07772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18592" *)
  wire _07773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18615" *)
  wire _07774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18615" *)
  wire _07775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18639" *)
  wire _07776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18639" *)
  wire _07777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18663" *)
  wire _07778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18663" *)
  wire _07779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18687" *)
  wire _07780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18687" *)
  wire _07781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18703" *)
  wire _07782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18703" *)
  wire _07783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18755" *)
  wire _07784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18760" *)
  wire _07785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18763" *)
  wire _07786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18766" *)
  wire _07787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18769" *)
  wire _07788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18772" *)
  wire _07789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18775" *)
  wire _07790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18778" *)
  wire _07791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18781" *)
  wire _07792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18784" *)
  wire _07793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18787" *)
  wire _07794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18790" *)
  wire _07795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18793" *)
  wire _07796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18796" *)
  wire _07797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18799" *)
  wire _07798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18802" *)
  wire _07799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18882" *)
  wire _07800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18899" *)
  wire _07801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18959" *)
  wire _07802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18990" *)
  wire _07803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19027" *)
  wire _07804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19062" *)
  wire _07805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19065" *)
  wire _07806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19103" *)
  wire _07807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19261" *)
  wire _07808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19576" *)
  wire _07809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19577" *)
  wire _07810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19577" *)
  wire _07811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19586" *)
  wire _07812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19609" *)
  wire _07813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19663" *)
  wire _07814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *)
  wire _07815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20098" *)
  wire _07816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20117" *)
  wire _07817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20136" *)
  wire _07818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20155" *)
  wire _07819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20174" *)
  wire _07820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20193" *)
  wire _07821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20212" *)
  wire _07822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20231" *)
  wire _07823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20250" *)
  wire _07824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20269" *)
  wire _07825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20288" *)
  wire _07826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20307" *)
  wire _07827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20326" *)
  wire _07828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20345" *)
  wire _07829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20364" *)
  wire _07830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20374" *)
  wire _07831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20374" *)
  wire _07832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20386" *)
  wire _07833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20386" *)
  wire _07834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20398" *)
  wire _07835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20398" *)
  wire _07836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20410" *)
  wire _07837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20410" *)
  wire _07838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20422" *)
  wire _07839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20422" *)
  wire _07840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20434" *)
  wire _07841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20434" *)
  wire _07842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20446" *)
  wire _07843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20446" *)
  wire _07844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20458" *)
  wire _07845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20458" *)
  wire _07846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20470" *)
  wire _07847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20470" *)
  wire _07848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20482" *)
  wire _07849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20482" *)
  wire _07850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20494" *)
  wire _07851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20494" *)
  wire _07852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20506" *)
  wire _07853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20506" *)
  wire _07854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20518" *)
  wire _07855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20518" *)
  wire _07856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20530" *)
  wire _07857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20530" *)
  wire _07858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20542" *)
  wire _07859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20542" *)
  wire _07860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20554" *)
  wire _07861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20554" *)
  wire _07862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20581" *)
  wire _07863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20583" *)
  wire _07864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20585" *)
  wire _07865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20587" *)
  wire _07866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20589" *)
  wire _07867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20591" *)
  wire _07868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20593" *)
  wire _07869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20595" *)
  wire _07870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20597" *)
  wire _07871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20599" *)
  wire _07872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20601" *)
  wire _07873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20603" *)
  wire _07874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20605" *)
  wire _07875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20607" *)
  wire _07876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20609" *)
  wire _07877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20819" *)
  wire _07878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20830" *)
  wire _07879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20830" *)
  wire _07880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *)
  wire _07881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *)
  wire _07882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *)
  wire _07883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *)
  wire _07884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20848" *)
  wire _07885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20848" *)
  wire _07886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *)
  wire _07887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *)
  wire _07888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20857" *)
  wire _07889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *)
  wire _07890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *)
  wire _07891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20866" *)
  wire _07892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20866" *)
  wire _07893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *)
  wire _07894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *)
  wire _07895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20875" *)
  wire _07896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *)
  wire _07897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *)
  wire _07898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20884" *)
  wire _07899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20884" *)
  wire _07900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *)
  wire _07901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *)
  wire _07902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *)
  wire _07903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20902" *)
  wire _07904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20902" *)
  wire _07905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20903" *)
  wire _07906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20903" *)
  wire _07907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20912" *)
  wire _07908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20913" *)
  wire _07909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20913" *)
  wire _07910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20922" *)
  wire _07911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20922" *)
  wire _07912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *)
  wire _07913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *)
  wire _07914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *)
  wire _07915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20940" *)
  wire _07916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20940" *)
  wire _07917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *)
  wire _07918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *)
  wire _07919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *)
  wire _07920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20958" *)
  wire _07921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20958" *)
  wire _07922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20959" *)
  wire _07923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20959" *)
  wire _07924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20959" *)
  wire _07925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *)
  wire _07926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *)
  wire _07927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20968" *)
  wire _07928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *)
  wire _07929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *)
  wire _07930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20977" *)
  wire _07931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20977" *)
  wire _07932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20978" *)
  wire _07933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20978" *)
  wire _07934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20987" *)
  wire _07935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20988" *)
  wire _07936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20988" *)
  wire _07937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20997" *)
  wire _07938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20997" *)
  wire _07939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *)
  wire _07940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *)
  wire _07941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *)
  wire _07942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *)
  wire _07943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *)
  wire _07944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21015" *)
  wire _07945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21015" *)
  wire _07946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *)
  wire _07947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *)
  wire _07948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *)
  wire _07949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21033" *)
  wire _07950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21033" *)
  wire _07951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21034" *)
  wire _07952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21034" *)
  wire _07953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *)
  wire _07954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *)
  wire _07955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *)
  wire _07956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *)
  wire _07957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *)
  wire _07958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *)
  wire _07959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21053" *)
  wire _07960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *)
  wire _07961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *)
  wire _07962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *)
  wire _07963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *)
  wire _07964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *)
  wire _07965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *)
  wire _07966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *)
  wire _07967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *)
  wire _07968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21073" *)
  wire _07969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21073" *)
  wire _07970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *)
  wire _07971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *)
  wire _07972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *)
  wire _07973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *)
  wire _07974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *)
  wire _07975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *)
  wire _07976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21092" *)
  wire _07977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21092" *)
  wire _07978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *)
  wire _07979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *)
  wire _07980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *)
  wire _07981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *)
  wire _07982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *)
  wire _07983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21102" *)
  wire _07984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *)
  wire _07985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *)
  wire _07986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21111" *)
  wire _07987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21111" *)
  wire _07988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *)
  wire _07989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *)
  wire _07990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *)
  wire _07991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21120" *)
  wire _07992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *)
  wire _07993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *)
  wire _07994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *)
  wire _07995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21179" *)
  wire _07996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21179" *)
  wire _07997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21260" *)
  wire _07998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21261" *)
  wire _07999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21261" *)
  wire _08000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *)
  wire _08001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *)
  wire _08002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21271" *)
  wire _08003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21271" *)
  wire _08004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *)
  wire _08005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *)
  wire _08006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21281" *)
  wire _08007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21281" *)
  wire _08008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *)
  wire _08009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *)
  wire _08010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21291" *)
  wire _08011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21291" *)
  wire _08012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *)
  wire _08013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *)
  wire _08014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21301" *)
  wire _08015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21301" *)
  wire _08016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *)
  wire _08017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *)
  wire _08018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21311" *)
  wire _08019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21311" *)
  wire _08020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *)
  wire _08021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *)
  wire _08022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21321" *)
  wire _08023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21321" *)
  wire _08024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *)
  wire _08025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *)
  wire _08026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21331" *)
  wire _08027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21331" *)
  wire _08028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *)
  wire _08029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *)
  wire _08030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21341" *)
  wire _08031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21341" *)
  wire _08032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *)
  wire _08033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *)
  wire _08034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21351" *)
  wire _08035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21351" *)
  wire _08036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *)
  wire _08037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *)
  wire _08038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21361" *)
  wire _08039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21361" *)
  wire _08040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *)
  wire _08041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *)
  wire _08042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21371" *)
  wire _08043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21371" *)
  wire _08044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *)
  wire _08045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *)
  wire _08046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21381" *)
  wire _08047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21381" *)
  wire _08048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *)
  wire _08049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *)
  wire _08050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21391" *)
  wire _08051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21391" *)
  wire _08052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *)
  wire _08053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *)
  wire _08054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21401" *)
  wire _08055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21401" *)
  wire _08056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *)
  wire _08057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *)
  wire _08058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21411" *)
  wire _08059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21411" *)
  wire _08060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *)
  wire _08061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *)
  wire _08062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21960" *)
  wire _08063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *)
  wire _08064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *)
  wire _08065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *)
  wire _08066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21964" *)
  wire _08067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21965" *)
  wire _08068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21965" *)
  wire _08069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21970" *)
  wire _08070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21971" *)
  wire _08071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21982" *)
  wire _08072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21982" *)
  wire _08073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21986" *)
  wire _08074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21987" *)
  wire _08075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21992" *)
  wire _08076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21992" *)
  wire _08077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21993" *)
  wire _08078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22001" *)
  wire _08079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22001" *)
  wire _08080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22002" *)
  wire _08081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22005" *)
  wire _08082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22006" *)
  wire _08083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22006" *)
  wire _08084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22006" *)
  wire _08085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22009" *)
  wire _08086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22010" *)
  wire _08087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22010" *)
  wire _08088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22013" *)
  wire _08089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22017" *)
  wire _08090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22017" *)
  wire _08091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22018" *)
  wire _08092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22024" *)
  wire _08093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22024" *)
  wire _08094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22025" *)
  wire _08095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22028" *)
  wire _08096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22029" *)
  wire _08097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22029" *)
  wire _08098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22029" *)
  wire _08099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22032" *)
  wire _08100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22033" *)
  wire _08101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22033" *)
  wire _08102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22036" *)
  wire _08103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22040" *)
  wire _08104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22040" *)
  wire _08105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22041" *)
  wire _08106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22047" *)
  wire _08107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22047" *)
  wire _08108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22048" *)
  wire _08109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22051" *)
  wire _08110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22052" *)
  wire _08111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22052" *)
  wire _08112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22052" *)
  wire _08113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22055" *)
  wire _08114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22056" *)
  wire _08115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22056" *)
  wire _08116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22059" *)
  wire _08117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22063" *)
  wire _08118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22063" *)
  wire _08119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22064" *)
  wire _08120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22070" *)
  wire _08121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22070" *)
  wire _08122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22071" *)
  wire _08123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22075" *)
  wire _08124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22076" *)
  wire _08125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22076" *)
  wire _08126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22079" *)
  wire _08127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22080" *)
  wire _08128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22081" *)
  wire _08129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22081" *)
  wire _08130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22083" *)
  wire _08131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22083" *)
  wire _08132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22087" *)
  wire _08133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22087" *)
  wire _08134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22090" *)
  wire _08135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22091" *)
  wire _08136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22091" *)
  wire _08137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22100" *)
  wire _08138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22100" *)
  wire _08139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22104" *)
  wire _08140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22105" *)
  wire _08141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22105" *)
  wire _08142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22108" *)
  wire _08143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22109" *)
  wire _08144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22110" *)
  wire _08145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22110" *)
  wire _08146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22112" *)
  wire _08147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22112" *)
  wire _08148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22116" *)
  wire _08149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22116" *)
  wire _08150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22119" *)
  wire _08151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22120" *)
  wire _08152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22120" *)
  wire _08153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22129" *)
  wire _08154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22129" *)
  wire _08155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22133" *)
  wire _08156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22133" *)
  wire _08157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22134" *)
  wire _08158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22135" *)
  wire _08159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22135" *)
  wire _08160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22137" *)
  wire _08161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22137" *)
  wire _08162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22141" *)
  wire _08163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22142" *)
  wire _08164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22142" *)
  wire _08165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22151" *)
  wire _08166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22154" *)
  wire _08167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22155" *)
  wire _08168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22155" *)
  wire _08169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22155" *)
  wire _08170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22158" *)
  wire _08171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22159" *)
  wire _08172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22159" *)
  wire _08173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22162" *)
  wire _08174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22166" *)
  wire _08175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22166" *)
  wire _08176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22167" *)
  wire _08177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22173" *)
  wire _08178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22173" *)
  wire _08179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22174" *)
  wire _08180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22177" *)
  wire _08181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22178" *)
  wire _08182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22178" *)
  wire _08183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22178" *)
  wire _08184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22181" *)
  wire _08185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22182" *)
  wire _08186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22182" *)
  wire _08187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22185" *)
  wire _08188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22189" *)
  wire _08189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22189" *)
  wire _08190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22190" *)
  wire _08191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22196" *)
  wire _08192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22196" *)
  wire _08193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22197" *)
  wire _08194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22201" *)
  wire _08195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22202" *)
  wire _08196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22202" *)
  wire _08197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22206" *)
  wire _08198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22207" *)
  wire _08199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22208" *)
  wire _08200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22208" *)
  wire _08201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22210" *)
  wire _08202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22210" *)
  wire _08203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22214" *)
  wire _08204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22214" *)
  wire _08205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22218" *)
  wire _08206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22219" *)
  wire _08207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22219" *)
  wire _08208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22228" *)
  wire _08209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22228" *)
  wire _08210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22231" *)
  wire _08211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22232" *)
  wire _08212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22232" *)
  wire _08213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22232" *)
  wire _08214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22235" *)
  wire _08215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22236" *)
  wire _08216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22236" *)
  wire _08217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22239" *)
  wire _08218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22243" *)
  wire _08219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22243" *)
  wire _08220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22244" *)
  wire _08221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22250" *)
  wire _08222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22250" *)
  wire _08223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22251" *)
  wire _08224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22254" *)
  wire _08225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22255" *)
  wire _08226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22255" *)
  wire _08227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22255" *)
  wire _08228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22258" *)
  wire _08229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22259" *)
  wire _08230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22259" *)
  wire _08231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22262" *)
  wire _08232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22266" *)
  wire _08233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22266" *)
  wire _08234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22267" *)
  wire _08235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22273" *)
  wire _08236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22273" *)
  wire _08237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22274" *)
  wire _08238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22278" *)
  wire _08239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22279" *)
  wire _08240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22279" *)
  wire _08241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22283" *)
  wire _08242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22284" *)
  wire _08243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22285" *)
  wire _08244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22285" *)
  wire _08245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22287" *)
  wire _08246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22287" *)
  wire _08247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22291" *)
  wire _08248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22291" *)
  wire _08249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22295" *)
  wire _08250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22296" *)
  wire _08251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22296" *)
  wire _08252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22305" *)
  wire _08253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22305" *)
  wire _08254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22308" *)
  wire _08255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22309" *)
  wire _08256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22309" *)
  wire _08257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22309" *)
  wire _08258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22312" *)
  wire _08259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22313" *)
  wire _08260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22313" *)
  wire _08261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22316" *)
  wire _08262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22320" *)
  wire _08263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22320" *)
  wire _08264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22321" *)
  wire _08265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22327" *)
  wire _08266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22327" *)
  wire _08267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22328" *)
  wire _08268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22331" *)
  wire _08269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22332" *)
  wire _08270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22332" *)
  wire _08271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22332" *)
  wire _08272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22335" *)
  wire _08273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22336" *)
  wire _08274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22336" *)
  wire _08275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22339" *)
  wire _08276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22343" *)
  wire _08277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22343" *)
  wire _08278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22344" *)
  wire _08279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22350" *)
  wire _08280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22350" *)
  wire _08281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22351" *)
  wire _08282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22354" *)
  wire _08283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22355" *)
  wire _08284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22355" *)
  wire _08285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22355" *)
  wire _08286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22358" *)
  wire _08287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22359" *)
  wire _08288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22359" *)
  wire _08289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22362" *)
  wire _08290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22366" *)
  wire _08291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22366" *)
  wire _08292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22367" *)
  wire _08293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22373" *)
  wire _08294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22373" *)
  wire _08295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22374" *)
  wire _08296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22486" *)
  wire _08297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22486" *)
  wire _08298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22486" *)
  wire _08299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22543" *)
  wire _08300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22550" *)
  wire _08301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22552" *)
  wire _08302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22553" *)
  wire _08303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22579" *)
  wire _08304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22586" *)
  wire _08305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22586" *)
  wire _08306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22590" *)
  wire _08307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22594" *)
  wire _08308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22597" *)
  wire _08309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22615" *)
  wire _08310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22620" *)
  wire _08311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22625" *)
  wire _08312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22634" *)
  wire _08313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22637" *)
  wire _08314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22650" *)
  wire _08315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22653" *)
  wire _08316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22666" *)
  wire _08317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22669" *)
  wire _08318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22702" *)
  wire _08319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22705" *)
  wire _08320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22720" *)
  wire _08321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22723" *)
  wire _08322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22738" *)
  wire _08323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22741" *)
  wire _08324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22747" *)
  wire _08325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22753" *)
  wire _08326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22758" *)
  wire _08327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22758" *)
  wire _08328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22761" *)
  wire _08329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22765" *)
  wire _08330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22768" *)
  wire _08331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22781" *)
  wire _08332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22798" *)
  wire _08333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22798" *)
  wire _08334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22801" *)
  wire _08335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22807" *)
  wire _08336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22811" *)
  wire _08337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22823" *)
  wire _08338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22823" *)
  wire _08339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22826" *)
  wire _08340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22830" *)
  wire _08341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22833" *)
  wire _08342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22837" *)
  wire _08343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22879" *)
  wire _08344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22880" *)
  wire _08345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22880" *)
  wire _08346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22880" *)
  wire _08347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22883" *)
  wire _08348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22883" *)
  wire _08349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22887" *)
  wire _08350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22893" *)
  wire _08351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22896" *)
  wire _08352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22896" *)
  wire _08353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22899" *)
  wire _08354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22899" *)
  wire _08355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22906" *)
  wire _08356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22906" *)
  wire _08357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22909" *)
  wire _08358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22909" *)
  wire _08359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22916" *)
  wire _08360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *)
  wire _08361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *)
  wire _08362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22923" *)
  wire _08363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22923" *)
  wire _08364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22925" *)
  wire _08365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22925" *)
  wire _08366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22927" *)
  wire _08367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22929" *)
  wire _08368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22932" *)
  wire _08369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22932" *)
  wire _08370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22935" *)
  wire _08371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22935" *)
  wire _08372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22948" *)
  wire _08373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22948" *)
  wire _08374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22951" *)
  wire _08375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22951" *)
  wire _08376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22966" *)
  wire _08377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22966" *)
  wire _08378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22969" *)
  wire _08379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22969" *)
  wire _08380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22976" *)
  wire _08381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22976" *)
  wire _08382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22976" *)
  wire _08383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22977" *)
  wire _08384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22978" *)
  wire _08385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22978" *)
  wire _08386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22978" *)
  wire _08387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22982" *)
  wire _08388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22982" *)
  wire _08389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22986" *)
  wire _08390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22992" *)
  wire _08391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22995" *)
  wire _08392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22995" *)
  wire _08393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22998" *)
  wire _08394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22998" *)
  wire _08395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *)
  wire _08396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *)
  wire _08397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *)
  wire _08398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *)
  wire _08399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23009" *)
  wire _08400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23009" *)
  wire _08401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23010" *)
  wire _08402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23017" *)
  wire _08403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23017" *)
  wire _08404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23020" *)
  wire _08405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23020" *)
  wire _08406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23027" *)
  wire _08407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23027" *)
  wire _08408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23030" *)
  wire _08409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23030" *)
  wire _08410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23037" *)
  wire _08411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23037" *)
  wire _08412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23037" *)
  wire _08413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23038" *)
  wire _08414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23039" *)
  wire _08415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23039" *)
  wire _08416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23039" *)
  wire _08417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23043" *)
  wire _08418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23043" *)
  wire _08419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23047" *)
  wire _08420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23053" *)
  wire _08421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23056" *)
  wire _08422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23056" *)
  wire _08423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23059" *)
  wire _08424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23059" *)
  wire _08425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23066" *)
  wire _08426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23066" *)
  wire _08427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23066" *)
  wire _08428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23067" *)
  wire _08429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23068" *)
  wire _08430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23068" *)
  wire _08431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23068" *)
  wire _08432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23072" *)
  wire _08433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23072" *)
  wire _08434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23076" *)
  wire _08435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23082" *)
  wire _08436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23085" *)
  wire _08437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23085" *)
  wire _08438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23088" *)
  wire _08439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23088" *)
  wire _08440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *)
  wire _08441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *)
  wire _08442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *)
  wire _08443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *)
  wire _08444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *)
  wire _08445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *)
  wire _08446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *)
  wire _08447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *)
  wire _08448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23113" *)
  wire _08449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23114" *)
  wire _08450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23117" *)
  wire _08451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23118" *)
  wire _08452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23122" *)
  wire _08453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *)
  wire _08454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *)
  wire _08455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *)
  wire _08456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *)
  wire _08457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23129" *)
  wire _08458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23135" *)
  wire _08459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23135" *)
  wire _08460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23138" *)
  wire _08461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23138" *)
  wire _08462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23145" *)
  wire _08463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23145" *)
  wire _08464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23145" *)
  wire _08465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23146" *)
  wire _08466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23147" *)
  wire _08467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23147" *)
  wire _08468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23147" *)
  wire _08469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23151" *)
  wire _08470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23151" *)
  wire _08471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23153" *)
  wire _08472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23153" *)
  wire _08473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23160" *)
  wire _08474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23162" *)
  wire _08475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23165" *)
  wire _08476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23165" *)
  wire _08477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23168" *)
  wire _08478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23168" *)
  wire _08479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23175" *)
  wire _08480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23175" *)
  wire _08481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23178" *)
  wire _08482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23178" *)
  wire _08483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23185" *)
  wire _08484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23185" *)
  wire _08485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23188" *)
  wire _08486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23188" *)
  wire _08487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23195" *)
  wire _08488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23195" *)
  wire _08489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23198" *)
  wire _08490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23198" *)
  wire _08491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23300" *)
  wire _08492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23302" *)
  wire _08493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23302" *)
  wire _08494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23304" *)
  wire _08495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23306" *)
  wire _08496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23307" *)
  wire _08497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23307" *)
  wire _08498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23308" *)
  wire _08499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23309" *)
  wire _08500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23309" *)
  wire _08501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23316" *)
  wire _08502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23322" *)
  wire _08503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *)
  wire _08504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *)
  wire _08505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *)
  wire _08506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *)
  wire _08507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *)
  wire _08508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *)
  wire _08509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *)
  wire _08510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *)
  wire _08511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *)
  wire _08512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *)
  wire _08513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *)
  wire _08514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *)
  wire _08515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *)
  wire _08516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *)
  wire _08517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *)
  wire _08518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *)
  wire _08519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *)
  wire _08520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *)
  wire _08521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *)
  wire _08522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *)
  wire _08523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *)
  wire _08524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *)
  wire _08525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *)
  wire _08526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *)
  wire _08527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23356" *)
  wire _08528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23356" *)
  wire _08529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23356" *)
  wire _08530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *)
  wire _08531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *)
  wire _08532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *)
  wire _08533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *)
  wire _08534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23365" *)
  wire _08535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *)
  wire _08536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *)
  wire _08537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *)
  wire _08538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23369" *)
  wire _08539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23369" *)
  wire _08540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23371" *)
  wire _08541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23371" *)
  wire _08542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23381" *)
  wire _08543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23382" *)
  wire _08544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23391" *)
  wire _08545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23391" *)
  wire _08546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23392" *)
  wire _08547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *)
  wire _08548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *)
  wire _08549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23410" *)
  wire _08550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23410" *)
  wire _08551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23411" *)
  wire _08552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *)
  wire _08553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *)
  wire _08554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23424" *)
  wire _08555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23424" *)
  wire _08556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23425" *)
  wire _08557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23425" *)
  wire _08558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *)
  wire _08559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *)
  wire _08560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23433" *)
  wire _08561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23433" *)
  wire _08562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23434" *)
  wire _08563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *)
  wire _08564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *)
  wire _08565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23439" *)
  wire _08566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23439" *)
  wire _08567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23441" *)
  wire _08568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23441" *)
  wire _08569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23451" *)
  wire _08570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23451" *)
  wire _08571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23452" *)
  wire _08572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23452" *)
  wire _08573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *)
  wire _08574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *)
  wire _08575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23463" *)
  wire _08576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23463" *)
  wire _08577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23464" *)
  wire _08578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23464" *)
  wire _08579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *)
  wire _08580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *)
  wire _08581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23479" *)
  wire _08582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23479" *)
  wire _08583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23480" *)
  wire _08584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23480" *)
  wire _08585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *)
  wire _08586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *)
  wire _08587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23490" *)
  wire _08588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23490" *)
  wire _08589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23491" *)
  wire _08590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23491" *)
  wire _08591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23496" *)
  wire _08592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23497" *)
  wire _08593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23498" *)
  wire _08594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *)
  wire _08595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *)
  wire _08596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23508" *)
  wire _08597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23509" *)
  wire _08598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *)
  wire _08599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *)
  wire _08600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23520" *)
  wire _08601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23521" *)
  wire _08602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *)
  wire _08603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *)
  wire _08604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23530" *)
  wire _08605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23541" *)
  wire _08606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23542" *)
  wire _08607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *)
  wire _08608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *)
  wire _08609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23552" *)
  wire _08610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *)
  wire _08611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *)
  wire _08612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *)
  wire _08613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23556" *)
  wire _08614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23562" *)
  wire _08615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23573" *)
  wire _08616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *)
  wire _08617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *)
  wire _08618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *)
  wire _08619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23582" *)
  wire _08620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *)
  wire _08621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *)
  wire _08622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *)
  wire _08623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23591" *)
  wire _08624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23591" *)
  wire _08625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *)
  wire _08626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *)
  wire _08627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *)
  wire _08628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23595" *)
  wire _08629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23599" *)
  wire _08630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23602" *)
  wire _08631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23606" *)
  wire _08632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23620" *)
  wire _08633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23622" *)
  wire _08634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23625" *)
  wire _08635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23636" *)
  wire _08636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23639" *)
  wire _08637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23640" *)
  wire _08638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23640" *)
  wire _08639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23641" *)
  wire _08640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23642" *)
  wire _08641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23642" *)
  wire _08642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23645" *)
  wire _08643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23646" *)
  wire _08644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23646" *)
  wire _08645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23647" *)
  wire _08646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23647" *)
  wire _08647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23647" *)
  wire _08648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23651" *)
  wire _08649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23651" *)
  wire _08650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23652" *)
  wire _08651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23653" *)
  wire _08652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23653" *)
  wire _08653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23659" *)
  wire _08654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23662" *)
  wire _08655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23663" *)
  wire _08656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23663" *)
  wire _08657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23664" *)
  wire _08658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23665" *)
  wire _08659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23665" *)
  wire _08660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23668" *)
  wire _08661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23669" *)
  wire _08662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23669" *)
  wire _08663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23670" *)
  wire _08664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23670" *)
  wire _08665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23670" *)
  wire _08666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23674" *)
  wire _08667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23674" *)
  wire _08668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23675" *)
  wire _08669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23676" *)
  wire _08670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23676" *)
  wire _08671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23682" *)
  wire _08672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23685" *)
  wire _08673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23686" *)
  wire _08674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23686" *)
  wire _08675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23687" *)
  wire _08676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23688" *)
  wire _08677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23688" *)
  wire _08678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23691" *)
  wire _08679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23692" *)
  wire _08680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23692" *)
  wire _08681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23693" *)
  wire _08682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23693" *)
  wire _08683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23693" *)
  wire _08684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23697" *)
  wire _08685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23697" *)
  wire _08686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23698" *)
  wire _08687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23699" *)
  wire _08688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23699" *)
  wire _08689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23705" *)
  wire _08690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23708" *)
  wire _08691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23709" *)
  wire _08692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23709" *)
  wire _08693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23710" *)
  wire _08694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23711" *)
  wire _08695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23711" *)
  wire _08696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23714" *)
  wire _08697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23715" *)
  wire _08698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23715" *)
  wire _08699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23716" *)
  wire _08700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23716" *)
  wire _08701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23716" *)
  wire _08702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23720" *)
  wire _08703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23720" *)
  wire _08704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23721" *)
  wire _08705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23722" *)
  wire _08706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23722" *)
  wire _08707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23727" *)
  wire _08708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23727" *)
  wire _08709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23728" *)
  wire _08710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23728" *)
  wire _08711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23728" *)
  wire _08712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23729" *)
  wire _08713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23730" *)
  wire _08714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23731" *)
  wire _08715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23732" *)
  wire _08716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23733" *)
  wire _08717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23734" *)
  wire _08718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23734" *)
  wire _08719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *)
  wire _08720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23743" *)
  wire _08721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23744" *)
  wire _08722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23745" *)
  wire _08723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23745" *)
  wire _08724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23751" *)
  wire _08725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23751" *)
  wire _08726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23751" *)
  wire _08727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23754" *)
  wire _08728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23755" *)
  wire _08729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23755" *)
  wire _08730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23756" *)
  wire _08731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23757" *)
  wire _08732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23757" *)
  wire _08733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23760" *)
  wire _08734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23761" *)
  wire _08735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23761" *)
  wire _08736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23762" *)
  wire _08737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23762" *)
  wire _08738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23762" *)
  wire _08739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23766" *)
  wire _08740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23766" *)
  wire _08741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23767" *)
  wire _08742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23768" *)
  wire _08743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23768" *)
  wire _08744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23774" *)
  wire _08745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23774" *)
  wire _08746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23774" *)
  wire _08747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23777" *)
  wire _08748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23778" *)
  wire _08749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23778" *)
  wire _08750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23779" *)
  wire _08751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23780" *)
  wire _08752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23780" *)
  wire _08753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23783" *)
  wire _08754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23784" *)
  wire _08755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23784" *)
  wire _08756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23785" *)
  wire _08757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23785" *)
  wire _08758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23785" *)
  wire _08759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23789" *)
  wire _08760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23789" *)
  wire _08761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23790" *)
  wire _08762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23791" *)
  wire _08763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23791" *)
  wire _08764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23797" *)
  wire _08765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23800" *)
  wire _08766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23801" *)
  wire _08767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23801" *)
  wire _08768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23802" *)
  wire _08769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23803" *)
  wire _08770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23803" *)
  wire _08771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23806" *)
  wire _08772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23807" *)
  wire _08773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23807" *)
  wire _08774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23808" *)
  wire _08775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23808" *)
  wire _08776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23808" *)
  wire _08777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23812" *)
  wire _08778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23812" *)
  wire _08779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23813" *)
  wire _08780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23814" *)
  wire _08781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23814" *)
  wire _08782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23820" *)
  wire _08783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23823" *)
  wire _08784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23824" *)
  wire _08785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23824" *)
  wire _08786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23825" *)
  wire _08787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23826" *)
  wire _08788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23826" *)
  wire _08789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23829" *)
  wire _08790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23830" *)
  wire _08791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23830" *)
  wire _08792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23831" *)
  wire _08793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23831" *)
  wire _08794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23831" *)
  wire _08795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23835" *)
  wire _08796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23835" *)
  wire _08797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23836" *)
  wire _08798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23837" *)
  wire _08799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23837" *)
  wire _08800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23843" *)
  wire _08801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23843" *)
  wire _08802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23843" *)
  wire _08803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23846" *)
  wire _08804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23847" *)
  wire _08805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23847" *)
  wire _08806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23848" *)
  wire _08807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23849" *)
  wire _08808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23849" *)
  wire _08809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23852" *)
  wire _08810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23853" *)
  wire _08811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23853" *)
  wire _08812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23854" *)
  wire _08813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23854" *)
  wire _08814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23854" *)
  wire _08815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23858" *)
  wire _08816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23858" *)
  wire _08817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23859" *)
  wire _08818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23860" *)
  wire _08819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23860" *)
  wire _08820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23866" *)
  wire _08821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23869" *)
  wire _08822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23870" *)
  wire _08823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23870" *)
  wire _08824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23871" *)
  wire _08825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23872" *)
  wire _08826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23872" *)
  wire _08827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23875" *)
  wire _08828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23876" *)
  wire _08829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23876" *)
  wire _08830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23877" *)
  wire _08831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23877" *)
  wire _08832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23877" *)
  wire _08833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23881" *)
  wire _08834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23881" *)
  wire _08835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23882" *)
  wire _08836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23883" *)
  wire _08837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23883" *)
  wire _08838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23889" *)
  wire _08839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23892" *)
  wire _08840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23893" *)
  wire _08841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23893" *)
  wire _08842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23894" *)
  wire _08843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23895" *)
  wire _08844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23895" *)
  wire _08845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23898" *)
  wire _08846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23899" *)
  wire _08847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23899" *)
  wire _08848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23900" *)
  wire _08849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23900" *)
  wire _08850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23900" *)
  wire _08851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23904" *)
  wire _08852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23904" *)
  wire _08853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23905" *)
  wire _08854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23906" *)
  wire _08855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23906" *)
  wire _08856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23912" *)
  wire _08857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23912" *)
  wire _08858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23912" *)
  wire _08859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23915" *)
  wire _08860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23916" *)
  wire _08861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23916" *)
  wire _08862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23917" *)
  wire _08863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23918" *)
  wire _08864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23918" *)
  wire _08865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23921" *)
  wire _08866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23922" *)
  wire _08867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23922" *)
  wire _08868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23923" *)
  wire _08869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23923" *)
  wire _08870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23923" *)
  wire _08871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23927" *)
  wire _08872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23927" *)
  wire _08873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23928" *)
  wire _08874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23929" *)
  wire _08875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23929" *)
  wire _08876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23935" *)
  wire _08877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23938" *)
  wire _08878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23939" *)
  wire _08879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23939" *)
  wire _08880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23940" *)
  wire _08881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23941" *)
  wire _08882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23941" *)
  wire _08883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23944" *)
  wire _08884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23945" *)
  wire _08885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23945" *)
  wire _08886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23946" *)
  wire _08887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23946" *)
  wire _08888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23946" *)
  wire _08889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23950" *)
  wire _08890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23950" *)
  wire _08891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23951" *)
  wire _08892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23952" *)
  wire _08893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23952" *)
  wire _08894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23958" *)
  wire _08895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23961" *)
  wire _08896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23962" *)
  wire _08897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23962" *)
  wire _08898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23963" *)
  wire _08899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23964" *)
  wire _08900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23964" *)
  wire _08901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23967" *)
  wire _08902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23968" *)
  wire _08903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23968" *)
  wire _08904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23969" *)
  wire _08905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23969" *)
  wire _08906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23969" *)
  wire _08907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23973" *)
  wire _08908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23973" *)
  wire _08909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23974" *)
  wire _08910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23975" *)
  wire _08911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23975" *)
  wire _08912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23981" *)
  wire _08913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23984" *)
  wire _08914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23985" *)
  wire _08915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23985" *)
  wire _08916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23986" *)
  wire _08917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23987" *)
  wire _08918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23987" *)
  wire _08919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23990" *)
  wire _08920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23991" *)
  wire _08921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23991" *)
  wire _08922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23992" *)
  wire _08923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23992" *)
  wire _08924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23992" *)
  wire _08925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23996" *)
  wire _08926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23996" *)
  wire _08927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23997" *)
  wire _08928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23998" *)
  wire _08929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23998" *)
  wire _08930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24003" *)
  wire _08931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24003" *)
  wire _08932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24008" *)
  wire _08933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24008" *)
  wire _08934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24013" *)
  wire _08935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24013" *)
  wire _08936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24018" *)
  wire _08937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24018" *)
  wire _08938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24023" *)
  wire _08939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24023" *)
  wire _08940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24028" *)
  wire _08941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24028" *)
  wire _08942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24035" *)
  wire _08943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24035" *)
  wire _08944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *)
  wire _08945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *)
  wire _08946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24043" *)
  wire _08947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24043" *)
  wire _08948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24048" *)
  wire _08949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24048" *)
  wire _08950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24053" *)
  wire _08951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24053" *)
  wire _08952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24060" *)
  wire _08953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24060" *)
  wire _08954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24063" *)
  wire _08955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24068" *)
  wire _08956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24068" *)
  wire _08957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24073" *)
  wire _08958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24073" *)
  wire _08959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24078" *)
  wire _08960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24078" *)
  wire _08961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24083" *)
  wire _08962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24083" *)
  wire _08963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24088" *)
  wire _08964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _08999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *)
  wire _09027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *)
  wire _09058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *)
  wire _09074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *)
  wire _09090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *)
  wire _09106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *)
  wire _09122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *)
  wire [14:0] _09150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *)
  wire [14:0] _09166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *)
  wire [14:0] _09167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *)
  wire [14:0] _09168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *)
  wire [14:0] _09169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *)
  wire [14:0] _09170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *)
  wire [14:0] _09171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *)
  wire [14:0] _09172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *)
  wire [14:0] _09173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *)
  wire [14:0] _09174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *)
  wire [14:0] _09175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *)
  wire [14:0] _09176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *)
  wire [14:0] _09177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *)
  wire [14:0] _09178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *)
  wire [14:0] _09179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *)
  wire [14:0] _09192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *)
  wire [14:0] _09205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *)
  wire [14:0] _09218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *)
  wire [14:0] _09231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *)
  wire [14:0] _09244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24335" *)
  wire [15:0] _09245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *)
  wire [3:0] _09261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *)
  wire [3:0] _09277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *)
  wire [3:0] _09293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *)
  wire [3:0] _09309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *)
  wire [3:0] _09325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *)
  wire [3:0] _09341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *)
  wire [3:0] _09357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *)
  wire [4:0] _09373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *)
  wire [6:0] _09388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24409" *)
  wire [8:0] _09389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24410" *)
  wire [8:0] _09390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24411" *)
  wire [8:0] _09391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *)
  wire [8:0] _09406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *)
  wire [8:0] _09421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *)
  wire [8:0] _09436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *)
  wire [8:0] _09451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8776" *)
  wire _09452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8799" *)
  wire _09453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8799" *)
  wire _09454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8807" *)
  wire _09455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8809" *)
  wire _09456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8818" *)
  wire _09457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8836" *)
  wire _09458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8837" *)
  wire _09459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8861" *)
  wire _09460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8872" *)
  wire _09461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8879" *)
  wire _09462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8883" *)
  wire _09463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8888" *)
  wire _09464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8894" *)
  wire _09465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8897" *)
  wire _09466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8898" *)
  wire _09467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8913" *)
  wire _09468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8923" *)
  wire _09469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8932" *)
  wire _09470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8947" *)
  wire _09471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8954" *)
  wire _09472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8964" *)
  wire _09473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8966" *)
  wire _09474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8977" *)
  wire _09475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8979" *)
  wire _09476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9007" *)
  wire _09477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9011" *)
  wire _09478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9025" *)
  wire _09479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9029" *)
  wire _09480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9045" *)
  wire _09481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9061" *)
  wire _09482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9071" *)
  wire _09483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9073" *)
  wire _09484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9081" *)
  wire _09485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9081" *)
  wire _09486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9082" *)
  wire _09487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9087" *)
  wire _09488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9087" *)
  wire _09489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9090" *)
  wire _09490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9090" *)
  wire _09491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9090" *)
  wire _09492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9096" *)
  wire _09493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9096" *)
  wire _09494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9099" *)
  wire _09495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9099" *)
  wire _09496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9099" *)
  wire _09497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9128" *)
  wire _09498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9133" *)
  wire _09499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9133" *)
  wire _09500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9167" *)
  wire _09501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9169" *)
  wire _09502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9173" *)
  wire _09503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9173" *)
  wire _09504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9175" *)
  wire _09505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9175" *)
  wire _09506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9176" *)
  wire _09507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9176" *)
  wire _09508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9178" *)
  wire _09509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9191" *)
  wire _09510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *)
  wire _09511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *)
  wire _09512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9227" *)
  wire _09513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9228" *)
  wire _09514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9228" *)
  wire _09515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9229" *)
  wire _09516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9229" *)
  wire _09517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9231" *)
  wire _09518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9231" *)
  wire _09519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9234" *)
  wire _09520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9234" *)
  wire _09521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9246" *)
  wire _09522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9266" *)
  wire _09523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9267" *)
  wire _09524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9270" *)
  wire _09525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9271" *)
  wire _09526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9271" *)
  wire _09527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *)
  wire _09528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *)
  wire _09529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *)
  wire _09530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *)
  wire _09531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9310" *)
  wire _09532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9312" *)
  wire _09533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9353" *)
  wire _09534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9364" *)
  wire _09535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9402" *)
  wire _09536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9481" *)
  wire _09537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9484" *)
  wire _09538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9489" *)
  wire _09539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *)
  wire _09540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *)
  wire _09541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9495" *)
  wire _09542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9497" *)
  wire _09543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9497" *)
  wire _09544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9501" *)
  wire _09545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9501" *)
  wire _09546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9501" *)
  wire _09547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9522" *)
  wire _09548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9540" *)
  wire _09549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9540" *)
  wire _09550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *)
  wire _09551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *)
  wire _09552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *)
  wire _09553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *)
  wire _09554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9543" *)
  wire _09555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9543" *)
  wire _09556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9544" *)
  wire _09557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9544" *)
  wire _09558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9562" *)
  wire _09559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9564" *)
  wire _09560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9568" *)
  wire _09561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9606" *)
  wire _09562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9647" *)
  wire _09563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9679" *)
  wire _09564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9714" *)
  wire _09565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9749" *)
  wire _09566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9852" *)
  wire _09567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9852" *)
  wire _09568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9854" *)
  wire _09569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9858" *)
  wire _09570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9861" *)
  wire _09571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9864" *)
  wire _09572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9869" *)
  wire _09573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9875" *)
  wire _09574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9879" *)
  wire _09575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9881" *)
  wire _09576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9884" *)
  wire _09577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9891" *)
  wire _09578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9891" *)
  wire _09579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9966" *)
  wire _09580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9966" *)
  wire _09581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9972" *)
  wire _09582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9972" *)
  wire _09583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9978" *)
  wire _09584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9978" *)
  wire _09585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9984" *)
  wire _09586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9984" *)
  wire _09587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9990" *)
  wire _09588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9990" *)
  wire _09589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9996" *)
  wire _09590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9996" *)
  wire _09591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4123" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4134" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4145" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4156" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4166" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4179" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4024" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4035" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4046" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4057" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4068" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4079" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4090" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4101" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4112" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4012" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3383" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3384" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3385" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3386" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3387" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3388" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3374" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3375" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3376" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3377" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3378" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3379" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3380" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3381" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3382" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2716" *)
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4986" *)
  wire FpFloatToInt_16U_5U_10U_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5063" *)
  wire FpFloatToInt_16U_5U_10U_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5131" *)
  wire FpFloatToInt_16U_5U_10U_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5167" *)
  wire FpFloatToInt_16U_5U_10U_and_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5188" *)
  wire FpFloatToInt_16U_5U_10U_and_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5469" *)
  wire FpFloatToInt_16U_5U_10U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5174" *)
  wire FpFloatToInt_16U_5U_10U_and_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5139" *)
  wire FpFloatToInt_16U_5U_10U_and_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5085" *)
  wire FpFloatToInt_16U_5U_10U_and_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5008" *)
  wire FpFloatToInt_16U_5U_10U_and_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4957" *)
  wire FpFloatToInt_16U_5U_10U_and_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4903" *)
  wire FpFloatToInt_16U_5U_10U_and_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5468" *)
  wire FpFloatToInt_16U_5U_10U_and_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4857" *)
  wire FpFloatToInt_16U_5U_10U_and_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4858" *)
  wire FpFloatToInt_16U_5U_10U_and_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4878" *)
  wire FpFloatToInt_16U_5U_10U_and_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4879" *)
  wire FpFloatToInt_16U_5U_10U_and_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4895" *)
  wire FpFloatToInt_16U_5U_10U_and_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4896" *)
  wire FpFloatToInt_16U_5U_10U_and_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4940" *)
  wire FpFloatToInt_16U_5U_10U_and_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4859" *)
  wire FpFloatToInt_16U_5U_10U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4941" *)
  wire FpFloatToInt_16U_5U_10U_and_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4984" *)
  wire FpFloatToInt_16U_5U_10U_and_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4985" *)
  wire FpFloatToInt_16U_5U_10U_and_42_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5061" *)
  wire FpFloatToInt_16U_5U_10U_and_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5062" *)
  wire FpFloatToInt_16U_5U_10U_and_44_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5129" *)
  wire FpFloatToInt_16U_5U_10U_and_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5130" *)
  wire FpFloatToInt_16U_5U_10U_and_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5165" *)
  wire FpFloatToInt_16U_5U_10U_and_47_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5166" *)
  wire FpFloatToInt_16U_5U_10U_and_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5186" *)
  wire FpFloatToInt_16U_5U_10U_and_49_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5187" *)
  wire FpFloatToInt_16U_5U_10U_and_50_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5172" *)
  wire FpFloatToInt_16U_5U_10U_and_51_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5173" *)
  wire FpFloatToInt_16U_5U_10U_and_52_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5137" *)
  wire FpFloatToInt_16U_5U_10U_and_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5138" *)
  wire FpFloatToInt_16U_5U_10U_and_54_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5083" *)
  wire FpFloatToInt_16U_5U_10U_and_55_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5084" *)
  wire FpFloatToInt_16U_5U_10U_and_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5006" *)
  wire FpFloatToInt_16U_5U_10U_and_57_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5007" *)
  wire FpFloatToInt_16U_5U_10U_and_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4955" *)
  wire FpFloatToInt_16U_5U_10U_and_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4880" *)
  wire FpFloatToInt_16U_5U_10U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4956" *)
  wire FpFloatToInt_16U_5U_10U_and_60_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4901" *)
  wire FpFloatToInt_16U_5U_10U_and_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4902" *)
  wire FpFloatToInt_16U_5U_10U_and_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4897" *)
  wire FpFloatToInt_16U_5U_10U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4942" *)
  wire FpFloatToInt_16U_5U_10U_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5467" *)
  wire FpFloatToInt_16U_5U_10U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3242" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3245" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3248" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3251" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3254" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3257" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2713" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3218" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3221" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3224" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3227" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3230" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3233" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3236" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3239" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3260" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4048" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4059" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4070" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4081" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4092" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4103" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4114" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4014" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4125" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4136" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4147" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4158" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4168" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_44_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4181" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_47_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4026" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4037" *)
  wire FpFloatToInt_16U_5U_10U_else_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3460" *)
  wire FpFloatToInt_16U_5U_10U_if_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3241" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3244" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3247" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3250" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3253" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3256" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2715" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3217" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3220" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3223" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3226" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3229" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3232" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3235" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3238" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3259" *)
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1607" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3058" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1606" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3061" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1605" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3055" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1604" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3049" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1603" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3045" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1602" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3043" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1616" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3024" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1615" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3025" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1614" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3028" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1613" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3031" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1612" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3036" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1611" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3040" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1610" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3044" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1609" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3048" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1608" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3052" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1601" *)
  reg FpFloatToInt_16U_5U_10U_internal_int_0_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3037" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_0_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3153" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3156" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3159" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3162" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3165" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3168" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2712" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3129" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3132" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3135" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3138" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3141" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3144" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3147" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3150" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3171" *)
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2504" *)
  wire FpFloatToInt_16U_5U_10U_internal_int_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4167" *)
  wire FpFloatToInt_16U_5U_10U_mux_102_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4180" *)
  wire FpFloatToInt_16U_5U_10U_mux_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4025" *)
  wire FpFloatToInt_16U_5U_10U_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4036" *)
  wire FpFloatToInt_16U_5U_10U_mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4047" *)
  wire FpFloatToInt_16U_5U_10U_mux_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4058" *)
  wire FpFloatToInt_16U_5U_10U_mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4069" *)
  wire FpFloatToInt_16U_5U_10U_mux_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4080" *)
  wire FpFloatToInt_16U_5U_10U_mux_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4013" *)
  wire FpFloatToInt_16U_5U_10U_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4091" *)
  wire FpFloatToInt_16U_5U_10U_mux_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4102" *)
  wire FpFloatToInt_16U_5U_10U_mux_60_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4113" *)
  wire FpFloatToInt_16U_5U_10U_mux_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4124" *)
  wire FpFloatToInt_16U_5U_10U_mux_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4135" *)
  wire FpFloatToInt_16U_5U_10U_mux_81_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4146" *)
  wire FpFloatToInt_16U_5U_10U_mux_88_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4157" *)
  wire FpFloatToInt_16U_5U_10U_mux_95_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1670" *)
  reg [14:0] FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3034" *)
  wire FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3035" *)
  wire FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5470" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5189" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5175" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5168" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5140" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5132" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5086" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5064" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5009" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4987" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4958" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4943" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4904" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4898" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4881" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4860" *)
  wire FpFloatToInt_16U_5U_10U_o_int_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2623" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2624" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2625" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2626" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2627" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2628" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2615" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2616" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2617" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2618" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2619" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2620" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2621" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2622" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5466" *)
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3738" *)
  wire FpFloatToInt_16U_5U_10U_shift_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3523" *)
  wire FpFloatToInt_16U_5U_10U_shift_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3739" *)
  wire FpFloatToInt_16U_5U_10U_shift_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5249" *)
  wire FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2696" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2697" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2698" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2699" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5473" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2700" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5161" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2701" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2702" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2703" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2704" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2705" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2706" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2707" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4853" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4720" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1970" *)
  reg [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5266" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5136" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5160" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5171" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5185" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5472" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4852" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4877" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4900" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4939" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4954" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4983" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5060" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5082" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5128" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1861" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1869" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1877" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1885" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1893" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1901" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1791" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1800" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1807" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1815" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1821" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1829" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1837" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1845" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1853" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1909" *)
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1790" *)
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1799" *)
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1806" *)
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1852" *)
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3455" *)
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3456" *)
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_15_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3457" *)
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_22_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3453" *)
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2610" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3360" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3362" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3364" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3366" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3368" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3370" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3342" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3344" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3346" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3348" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3350" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3352" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3354" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3356" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3358" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3372" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2598" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2599" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2600" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2601" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2602" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2603" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2604" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2605" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2612" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2614" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2596" *)
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2717" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_int_mant_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2708" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_int_mant_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2710" *)
  wire [16:0] FpIntToFloat_17U_5U_10U_else_int_mant_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6216" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5301" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6225" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6231" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5233" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6237" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5355" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6243" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6249" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6255" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6261" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6267" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6273" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6279" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5252" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5274" *)
  wire FpIntToFloat_17U_5U_10U_else_mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1389" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1394" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1453" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1461" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1471" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1478" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1486" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1493" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1400" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1406" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1413" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1419" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1427" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1434" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1439" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1445" *)
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3533" *)
  wire FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3477" *)
  wire FpIntToFloat_17U_5U_10U_if_and_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3775" *)
  wire FpIntToFloat_17U_5U_10U_if_and_18_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3778" *)
  wire FpIntToFloat_17U_5U_10U_if_and_22_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3776" *)
  wire FpIntToFloat_17U_5U_10U_if_and_27_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3532" *)
  wire FpIntToFloat_17U_5U_10U_if_and_31_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3501" *)
  wire FpIntToFloat_17U_5U_10U_if_and_33_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3781" *)
  wire FpIntToFloat_17U_5U_10U_if_and_36_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3728" *)
  wire FpIntToFloat_17U_5U_10U_if_nor_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3753" *)
  wire FpIntToFloat_17U_5U_10U_if_nor_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3069" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1447" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1862" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3070" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1455" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1870" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3071" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1463" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1878" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3072" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1473" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1886" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1480" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3073" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1894" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3074" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1488" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1902" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1792" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1801" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1808" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3065" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1408" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1816" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1822" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3066" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1421" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1830" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3067" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1429" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1838" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3068" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1436" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1846" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1854" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3760" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3520" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2532" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_and_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3720" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_and_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3783" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_and_23_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3774" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_and_26_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3780" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_and_28_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2530" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3075" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1495" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1910" *)
  reg FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3522" *)
  wire FpIntToFloat_17U_5U_10U_is_inf_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5383" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5371" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5361" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5347" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5332" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5447" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5321" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5305" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5294" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5278" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5261" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5240" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5439" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5430" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5410" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5402" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2884" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2887" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2890" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2893" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2896" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2869" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2899" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2902" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2905" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2908" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2911" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2914" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2872" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2875" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2878" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2881" *)
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5320" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5304" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5293" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5277" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5260" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5239" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5438" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5429" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5409" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5401" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5382" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5370" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5360" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5346" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5331" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5446" *)
  wire FpIntToFloat_17U_5U_10U_o_expo_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3203" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3205" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3207" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3209" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3211" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3213" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3185" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3187" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3189" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3191" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3193" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3195" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3197" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3199" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3201" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3215" *)
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3307" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3312" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3317" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3322" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3327" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3332" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3262" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3267" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3272" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3277" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3282" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3287" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3292" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3297" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3302" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3337" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3308" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3313" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3318" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3323" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3328" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3333" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3263" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3268" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3273" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3278" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3283" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3288" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3293" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3298" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3303" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1745" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1751" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1757" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1763" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1769" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1775" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1692" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1698" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1704" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1710" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1716" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1721" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1727" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1733" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1739" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1781" *)
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3338" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3310" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3315" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3320" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3325" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3330" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3335" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3265" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3270" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3275" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3280" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3285" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3290" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3295" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3300" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3305" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3340" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3311" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3316" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3321" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3326" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3331" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3336" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3266" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3271" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3276" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3281" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3286" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3291" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3296" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3301" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3306" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3341" *)
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2376" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2372" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2368" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2364" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2360" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2356" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2412" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2408" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2404" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2400" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2396" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2392" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2388" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2384" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2380" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2352" *)
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3309" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3314" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3319" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3324" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3329" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3334" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3264" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3269" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3274" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3279" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3284" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3289" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3294" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3299" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3304" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3339" *)
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3178" *)
  wire FpMantRNE_17U_11U_else_carry_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3179" *)
  wire FpMantRNE_17U_11U_else_carry_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3180" *)
  wire FpMantRNE_17U_11U_else_carry_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3181" *)
  wire FpMantRNE_17U_11U_else_carry_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3182" *)
  wire FpMantRNE_17U_11U_else_carry_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3183" *)
  wire FpMantRNE_17U_11U_else_carry_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2718" *)
  wire FpMantRNE_17U_11U_else_carry_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2709" *)
  wire FpMantRNE_17U_11U_else_carry_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3172" *)
  wire FpMantRNE_17U_11U_else_carry_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3173" *)
  wire FpMantRNE_17U_11U_else_carry_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3174" *)
  wire FpMantRNE_17U_11U_else_carry_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3175" *)
  wire FpMantRNE_17U_11U_else_carry_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3176" *)
  wire FpMantRNE_17U_11U_else_carry_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3177" *)
  wire FpMantRNE_17U_11U_else_carry_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2711" *)
  wire FpMantRNE_17U_11U_else_carry_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3184" *)
  wire FpMantRNE_17U_11U_else_carry_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6223" *)
  wire FpMantRNE_17U_11U_else_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6229" *)
  wire FpMantRNE_17U_11U_else_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6235" *)
  wire FpMantRNE_17U_11U_else_mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5353" *)
  wire FpMantRNE_17U_11U_else_mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6241" *)
  wire FpMantRNE_17U_11U_else_mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5231" *)
  wire FpMantRNE_17U_11U_else_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6247" *)
  wire FpMantRNE_17U_11U_else_mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6253" *)
  wire FpMantRNE_17U_11U_else_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6259" *)
  wire FpMantRNE_17U_11U_else_mux_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6265" *)
  wire FpMantRNE_17U_11U_else_mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6271" *)
  wire FpMantRNE_17U_11U_else_mux_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6277" *)
  wire FpMantRNE_17U_11U_else_mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5250" *)
  wire FpMantRNE_17U_11U_else_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5272" *)
  wire FpMantRNE_17U_11U_else_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6214" *)
  wire FpMantRNE_17U_11U_else_mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5299" *)
  wire FpMantRNE_17U_11U_else_mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1747" *)
  reg FpMantRNE_24U_11U_else_carry_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3085" *)
  wire FpMantRNE_24U_11U_else_carry_10_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1753" *)
  reg FpMantRNE_24U_11U_else_carry_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3086" *)
  wire FpMantRNE_24U_11U_else_carry_11_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1759" *)
  reg FpMantRNE_24U_11U_else_carry_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3087" *)
  wire FpMantRNE_24U_11U_else_carry_12_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1765" *)
  reg FpMantRNE_24U_11U_else_carry_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3088" *)
  wire FpMantRNE_24U_11U_else_carry_13_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1771" *)
  reg FpMantRNE_24U_11U_else_carry_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3089" *)
  wire FpMantRNE_24U_11U_else_carry_14_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1777" *)
  reg FpMantRNE_24U_11U_else_carry_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3090" *)
  wire FpMantRNE_24U_11U_else_carry_15_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1694" *)
  reg FpMantRNE_24U_11U_else_carry_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3076" *)
  wire FpMantRNE_24U_11U_else_carry_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1700" *)
  reg FpMantRNE_24U_11U_else_carry_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3077" *)
  wire FpMantRNE_24U_11U_else_carry_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1706" *)
  reg FpMantRNE_24U_11U_else_carry_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3078" *)
  wire FpMantRNE_24U_11U_else_carry_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1712" *)
  reg FpMantRNE_24U_11U_else_carry_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3079" *)
  wire FpMantRNE_24U_11U_else_carry_4_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1718" *)
  reg FpMantRNE_24U_11U_else_carry_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3080" *)
  wire FpMantRNE_24U_11U_else_carry_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1723" *)
  reg FpMantRNE_24U_11U_else_carry_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3081" *)
  wire FpMantRNE_24U_11U_else_carry_6_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1729" *)
  reg FpMantRNE_24U_11U_else_carry_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3082" *)
  wire FpMantRNE_24U_11U_else_carry_7_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1735" *)
  reg FpMantRNE_24U_11U_else_carry_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3083" *)
  wire FpMantRNE_24U_11U_else_carry_8_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1741" *)
  reg FpMantRNE_24U_11U_else_carry_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3084" *)
  wire FpMantRNE_24U_11U_else_carry_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1783" *)
  reg FpMantRNE_24U_11U_else_carry_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3091" *)
  wire FpMantRNE_24U_11U_else_carry_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5748" *)
  wire FpMantRNE_24U_11U_else_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5741" *)
  wire FpMantRNE_24U_11U_else_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5736" *)
  wire FpMantRNE_24U_11U_else_mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5731" *)
  wire FpMantRNE_24U_11U_else_mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5726" *)
  wire FpMantRNE_24U_11U_else_mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5773" *)
  wire FpMantRNE_24U_11U_else_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5719" *)
  wire FpMantRNE_24U_11U_else_mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5714" *)
  wire FpMantRNE_24U_11U_else_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5709" *)
  wire FpMantRNE_24U_11U_else_mux_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5704" *)
  wire FpMantRNE_24U_11U_else_mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5699" *)
  wire FpMantRNE_24U_11U_else_mux_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5694" *)
  wire FpMantRNE_24U_11U_else_mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5768" *)
  wire FpMantRNE_24U_11U_else_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5763" *)
  wire FpMantRNE_24U_11U_else_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5758" *)
  wire FpMantRNE_24U_11U_else_mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5753" *)
  wire FpMantRNE_24U_11U_else_mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6086" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6095" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6104" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6113" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6122" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6131" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6005" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6014" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6023" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6032" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6041" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6050" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6059" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6068" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6077" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5996" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2275" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2271" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2267" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2263" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2259" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2255" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2311" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2307" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2303" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2299" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2295" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2291" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2287" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2283" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2279" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2315" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2297" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2293" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2289" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2285" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2281" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2317" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2277" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2273" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2269" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2265" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2261" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2257" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2313" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5997" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5998" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6006" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6007" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6015" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6016" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6024" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6025" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6033" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6034" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6042" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6043" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6051" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2309" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6052" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6060" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6061" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6069" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6070" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6078" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6079" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6087" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6088" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6096" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6097" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6105" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6106" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6114" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6115" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6123" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6124" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6132" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6133" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2305" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2301" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2240" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2239" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2238" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2237" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2236" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2235" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2249" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2248" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2247" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2246" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2245" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2244" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2243" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2242" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2241" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2250" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6280" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6281" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6282" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6283" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6284" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6285" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6286" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6287" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6288" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6289" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6290" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_42_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6291" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6292" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_44_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6293" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6294" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6295" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_47_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1738" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2957" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1744" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2959" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1750" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2961" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1756" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2963" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1762" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2965" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1768" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2967" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1774" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2969" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1780" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2971" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1691" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2941" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1697" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2943" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1703" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2945" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1709" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2947" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1715" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2949" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1720" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2951" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1726" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2953" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1732" *)
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2955" *)
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6073" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6082" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6091" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6001" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6100" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6109" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_157_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6118" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_169_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6127" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5992" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6010" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6019" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6028" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_49_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6037" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6046" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6055" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_85_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6064" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_97_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1654" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2067" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1651" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2070" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1648" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2073" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1645" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2076" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1642" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2079" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1639" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2082" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1682" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2037" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1679" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2042" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1676" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2045" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1673" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2048" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1669" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2051" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1666" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2055" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1663" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2058" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1660" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2061" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1657" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2064" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1636" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2085" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2996" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2997" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2998" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2999" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3000" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3001" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2987" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2988" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2989" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2990" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2991" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2992" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2993" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2994" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2995" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2986" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6040" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6049" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6058" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6067" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6076" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6085" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6094" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6103" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6112" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6121" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6004" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6130" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_30_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6013" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6022" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6031" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5995" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6081" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6090" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6099" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6108" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6117" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6126" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6000" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6009" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6018" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6027" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6036" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6045" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6054" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6063" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6072" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5991" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3449" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2280" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2276" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2272" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2268" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2264" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2260" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2316" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2312" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2308" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2304" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2300" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2296" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2292" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2288" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2284" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2256" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1947" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1950" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1953" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1956" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1959" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1964" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1916" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1921" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1924" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1927" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1932" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1935" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1938" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1941" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1944" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1911" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2375" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2278" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2132" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2131" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1652" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2371" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2274" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2134" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2133" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1649" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2367" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2270" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2136" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2135" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1646" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2363" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2266" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2138" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2137" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1643" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2359" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2262" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2140" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2139" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1640" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2354" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2258" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2142" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2141" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1637" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2410" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2314" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2114" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2113" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1680" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2406" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2310" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2116" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2115" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1677" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2403" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2306" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2118" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2117" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1674" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2399" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2302" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2120" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2119" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1671" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2395" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2298" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2122" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2121" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1667" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2391" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2294" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2124" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2123" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1664" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2387" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2290" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2126" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2125" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1661" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2383" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2286" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2128" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2127" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1658" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2379" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2282" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2130" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2129" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1655" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2351" *)
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2254" *)
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2144" *)
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2143" *)
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1634" *)
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2374" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1574" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2370" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1569" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2366" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1573" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2362" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1570" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2358" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1571" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2355" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1572" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2411" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1562" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2407" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1565" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2402" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1582" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2398" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1566" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2394" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1579" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2390" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1578" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2386" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1567" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2382" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1568" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2378" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1575" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2350" *)
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_5_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1617" *)
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3514" *)
  wire IntMulExt_33U_16U_49U_and_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3709" *)
  wire IntMulExt_33U_16U_49U_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1855" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_10_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1863" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_11_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1871" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_12_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1879" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_13_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1887" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_14_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1895" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_15_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1786" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1793" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1802" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1809" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_4_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2974" *)
  wire IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1817" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1823" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_6_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1831" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_7_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1839" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_8_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1847" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1903" *)
  reg [48:0] IntMulExt_33U_16U_49U_return_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2012" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2010" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2008" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1982" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1983" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1984" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3092" *)
  wire IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2005" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2003" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2030" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2031" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2028" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2026" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2024" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2022" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2020" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2018" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2016" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2014" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2033" *)
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2850" *)
  wire IntSaturation_17U_16U_and_11_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2847" *)
  wire IntSaturation_17U_16U_and_13_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2844" *)
  wire IntSaturation_17U_16U_and_15_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2841" *)
  wire IntSaturation_17U_16U_and_17_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2838" *)
  wire IntSaturation_17U_16U_and_19_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2865" *)
  wire IntSaturation_17U_16U_and_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2835" *)
  wire IntSaturation_17U_16U_and_21_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2832" *)
  wire IntSaturation_17U_16U_and_23_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2829" *)
  wire IntSaturation_17U_16U_and_25_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2826" *)
  wire IntSaturation_17U_16U_and_27_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2823" *)
  wire IntSaturation_17U_16U_and_29_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2820" *)
  wire IntSaturation_17U_16U_and_31_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3479" *)
  wire IntSaturation_17U_16U_and_33_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2862" *)
  wire IntSaturation_17U_16U_and_3_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2859" *)
  wire IntSaturation_17U_16U_and_5_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2856" *)
  wire IntSaturation_17U_16U_and_7_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2853" *)
  wire IntSaturation_17U_16U_and_9_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1624" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1623" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1622" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1621" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1620" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1619" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1633" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1632" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1631" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1630" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1629" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1628" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1627" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1626" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1625" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1618" *)
  reg [14:0] IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2849" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2852" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2855" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2858" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2861" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2864" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2822" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2825" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2828" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2831" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2834" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2837" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2840" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2843" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2846" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2819" *)
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2851" *)
  wire IntSaturation_17U_16U_o_and_11_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2848" *)
  wire IntSaturation_17U_16U_o_and_13_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2845" *)
  wire IntSaturation_17U_16U_o_and_15_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2842" *)
  wire IntSaturation_17U_16U_o_and_17_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2839" *)
  wire IntSaturation_17U_16U_o_and_19_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2866" *)
  wire IntSaturation_17U_16U_o_and_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2836" *)
  wire IntSaturation_17U_16U_o_and_21_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2833" *)
  wire IntSaturation_17U_16U_o_and_23_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2830" *)
  wire IntSaturation_17U_16U_o_and_25_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2827" *)
  wire IntSaturation_17U_16U_o_and_27_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2824" *)
  wire IntSaturation_17U_16U_o_and_29_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2821" *)
  wire IntSaturation_17U_16U_o_and_31_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2863" *)
  wire IntSaturation_17U_16U_o_and_3_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2860" *)
  wire IntSaturation_17U_16U_o_and_5_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2857" *)
  wire IntSaturation_17U_16U_o_and_7_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2854" *)
  wire IntSaturation_17U_16U_o_and_9_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6482" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6486" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6490" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6492" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6496" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6500" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6446" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6450" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6454" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6458" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6462" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6466" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6470" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6474" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6478" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6442" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4128" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4139" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4150" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6207" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4171" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4177" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4029" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4040" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4051" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4062" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4073" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4084" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4095" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4106" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4117" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4017" *)
  wire IntSaturation_17U_8U_IntSaturation_17U_8U_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6463" *)
  wire IntSaturation_17U_8U_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6467" *)
  wire IntSaturation_17U_8U_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6471" *)
  wire IntSaturation_17U_8U_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6475" *)
  wire IntSaturation_17U_8U_and_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6479" *)
  wire IntSaturation_17U_8U_and_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6443" *)
  wire IntSaturation_17U_8U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6483" *)
  wire IntSaturation_17U_8U_and_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6487" *)
  wire IntSaturation_17U_8U_and_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6491" *)
  wire IntSaturation_17U_8U_and_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6493" *)
  wire IntSaturation_17U_8U_and_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6497" *)
  wire IntSaturation_17U_8U_and_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6501" *)
  wire IntSaturation_17U_8U_and_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6447" *)
  wire IntSaturation_17U_8U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6451" *)
  wire IntSaturation_17U_8U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6455" *)
  wire IntSaturation_17U_8U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6459" *)
  wire IntSaturation_17U_8U_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3204" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3206" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3208" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3210" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3212" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3214" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3186" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3188" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3190" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3192" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3194" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3196" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3198" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3200" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3202" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3216" *)
  wire [6:0] IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1859" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2978" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1867" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2980" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1875" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2979" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1883" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2984" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1891" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2981" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1899" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2983" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1788" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3002" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1797" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3004" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1804" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3006" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1813" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2973" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1819" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3009" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1827" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2975" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1835" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2977" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1843" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2976" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1849" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3014" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1907" *)
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2982" *)
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_sva_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3519" *)
  wire IntShiftRightSat_49U_6U_17U_if_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3516" *)
  wire IntShiftRightSat_49U_6U_17U_if_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1438" *)
  reg IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3107" *)
  wire IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1443" *)
  reg IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3100" *)
  wire IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1451" *)
  reg IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3102" *)
  wire IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1459" *)
  reg IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3101" *)
  wire IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1469" *)
  reg IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3106" *)
  wire IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1476" *)
  reg IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3103" *)
  wire IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1484" *)
  reg IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3105" *)
  wire IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1388" *)
  reg IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3108" *)
  wire IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1393" *)
  reg IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3093" *)
  wire IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1399" *)
  reg IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3095" *)
  wire IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1404" *)
  reg IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3094" *)
  wire IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1411" *)
  reg IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3099" *)
  wire IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1417" *)
  reg IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3096" *)
  wire IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1425" *)
  reg IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3098" *)
  wire IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1432" *)
  reg IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3097" *)
  wire IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1491" *)
  reg IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3104" *)
  wire IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1592" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3016" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1521" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1522" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_11_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3017" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1590" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1591" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_12_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3018" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1526" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1527" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_13_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3019" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1588" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_14_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1589" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_14_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3020" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1536" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1537" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_15_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3021" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1504" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3003" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1599" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1600" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3005" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1560" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1561" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3007" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1597" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1598" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_4_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3008" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1555" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_5_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1556" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_5_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3010" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1595" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1596" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_6_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3011" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1513" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1514" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_7_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3012" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1593" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1594" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_8_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3013" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1547" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_9_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1548" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_9_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3015" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1585" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1586" *)
  reg IntShiftRightSat_49U_6U_17U_o_0_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3022" *)
  wire IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1441" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1856" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2420" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1449" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1864" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2419" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1457" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1872" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2418" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1467" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1880" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2417" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1474" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1888" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2416" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1482" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1896" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2415" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1387" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1787" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2429" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1391" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1794" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2428" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1398" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1803" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2427" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1402" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1810" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2426" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1410" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1818" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2425" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1415" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1824" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2424" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1423" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1832" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2423" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1430" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1840" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2422" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1437" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1848" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2421" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1489" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1904" *)
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2414" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1442" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1857" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_10_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1858" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_10_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2324" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1450" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1865" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_11_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1866" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_11_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2323" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1458" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1873" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_12_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1874" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_12_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2322" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1468" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1881" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_13_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1882" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_13_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2321" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1475" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1889" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_14_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1890" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_14_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2320" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1483" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1897" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_15_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1898" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_15_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2319" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1563" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1564" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2333" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1392" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1795" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1796" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2332" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1583" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1584" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2331" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1403" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1811" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_4_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1812" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_4_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2330" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1580" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_5_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1581" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_5_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2329" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1416" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1825" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_6_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1826" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_6_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2328" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1424" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1833" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1834" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_7_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2327" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1431" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1841" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1842" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_8_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2326" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1576" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_9_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1577" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_9_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2325" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1490" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1905" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1906" *)
  reg IntShiftRightSat_49U_6U_17U_o_16_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2318" *)
  wire IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2629" *)
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3454" *)
  wire IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3480" *)
  wire IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3465" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_103_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3481" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_107_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3482" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_108_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3483" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_109_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3484" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_111_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3485" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_112_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3486" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_114_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3478" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_115_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3749" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_90_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2520" *)
  wire IntShiftRightSat_49U_6U_17U_o_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3765" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_15_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3751" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3511" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3727" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3510" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_and_18_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3779" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_and_22_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3752" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_and_25_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3509" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5521" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5524" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5530" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5515" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5509" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5512" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5503" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5465" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5500" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5506" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5539" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5518" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_30_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5542" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5533" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5536" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5527" *)
  wire IntShiftRightSat_49U_6U_17U_oelse_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3116" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3118" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3117" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3122" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3119" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3121" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3124" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3109" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3111" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3110" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3115" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3112" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3114" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3113" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3123" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3120" *)
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2340" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2339" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2338" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2337" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2336" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2335" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2349" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2348" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2347" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2346" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2345" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2344" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2343" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2342" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2341" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2334" *)
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2442" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2440" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2438" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2436" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2434" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2432" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2460" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2458" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2456" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2454" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2452" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2450" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2448" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2446" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2444" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2430" *)
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3151" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3154" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3157" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3160" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3163" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3166" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3125" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3127" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3130" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3133" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3136" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3139" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3142" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3145" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3148" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3169" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3152" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3155" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3158" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3161" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3164" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3167" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3126" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3128" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3131" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3134" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3137" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3140" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3143" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3146" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3149" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3170" *)
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1963" *)
  reg IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5803" *)
  wire IsNaN_5U_10U_IsNaN_5U_10U_nand_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1920" *)
  reg IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5795" *)
  wire IsNaN_5U_10U_IsNaN_5U_10U_nand_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1915" *)
  reg IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5784" *)
  wire IsNaN_5U_10U_IsNaN_5U_10U_nand_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2508" *)
  wire IsNaN_5U_10U_aelse_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2516" *)
  wire IsNaN_5U_10U_aelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3462" *)
  wire IsNaN_5U_10U_aelse_or_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3461" *)
  wire IsNaN_5U_10U_aelse_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1541" *)
  reg IsNaN_5U_10U_land_10_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1542" *)
  reg IsNaN_5U_10U_land_10_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1518" *)
  reg IsNaN_5U_10U_land_11_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1519" *)
  reg IsNaN_5U_10U_land_11_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1538" *)
  reg IsNaN_5U_10U_land_12_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1539" *)
  reg IsNaN_5U_10U_land_12_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1523" *)
  reg IsNaN_5U_10U_land_13_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1524" *)
  reg IsNaN_5U_10U_land_13_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1528" *)
  reg IsNaN_5U_10U_land_14_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1529" *)
  reg IsNaN_5U_10U_land_14_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1534" *)
  reg IsNaN_5U_10U_land_15_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2251" *)
  wire IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1502" *)
  reg IsNaN_5U_10U_land_1_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2253" *)
  wire IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1505" *)
  reg IsNaN_5U_10U_land_2_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2252" *)
  wire IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1557" *)
  reg IsNaN_5U_10U_land_3_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1558" *)
  reg IsNaN_5U_10U_land_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1507" *)
  reg IsNaN_5U_10U_land_4_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1508" *)
  reg IsNaN_5U_10U_land_4_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1552" *)
  reg IsNaN_5U_10U_land_5_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1553" *)
  reg IsNaN_5U_10U_land_5_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1549" *)
  reg IsNaN_5U_10U_land_6_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1550" *)
  reg IsNaN_5U_10U_land_6_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1510" *)
  reg IsNaN_5U_10U_land_7_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1511" *)
  reg IsNaN_5U_10U_land_7_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1515" *)
  reg IsNaN_5U_10U_land_8_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1516" *)
  reg IsNaN_5U_10U_land_8_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1544" *)
  reg IsNaN_5U_10U_land_9_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1545" *)
  reg IsNaN_5U_10U_land_9_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1531" *)
  reg IsNaN_5U_10U_land_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1532" *)
  reg IsNaN_5U_10U_land_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1962" *)
  reg IsNaN_5U_10U_nor_14_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5799" *)
  wire IsNaN_5U_10U_nor_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1919" *)
  reg IsNaN_5U_10U_nor_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5791" *)
  wire IsNaN_5U_10U_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1914" *)
  reg IsNaN_5U_10U_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5778" *)
  wire IsNaN_5U_10U_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1929" *)
  reg IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:982" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:964" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:961" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:958" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:955" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:952" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:949" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:992" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:989" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:986" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:979" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:976" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:973" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:970" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:967" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:995" *)
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1749" *)
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1755" *)
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1761" *)
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1767" *)
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1773" *)
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1779" *)
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1696" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1702" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1708" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1714" *)
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1725" *)
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1731" *)
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1737" *)
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1743" *)
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1785" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1928" *)
  reg IsNaN_8U_23U_nor_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:983" *)
  wire IsNaN_8U_23U_nor_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3977" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3984" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3990" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3997" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4004" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4009" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3931" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3934" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3940" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3943" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3949" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3955" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3962" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3965" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3971" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3925" *)
  wire SetToInf_5U_10U_SetToInf_5U_10U_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5088" *)
  wire and_1004_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2781" *)
  wire and_1009_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2782" *)
  wire and_1011_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5133" *)
  wire and_1013_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3736" *)
  wire and_1021_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5141" *)
  wire and_1023_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5142" *)
  wire and_1027_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3496" *)
  wire and_1038_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3497" *)
  wire and_1039_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3737" *)
  wire and_1059_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2477" *)
  wire and_1069_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2783" *)
  wire and_1077_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2729" *)
  wire and_1078_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2476" *)
  wire and_1080_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2475" *)
  wire and_1084_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2785" *)
  wire and_1091_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2474" *)
  wire and_1093_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2473" *)
  wire and_1097_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2789" *)
  wire and_1104_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2472" *)
  wire and_1106_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2471" *)
  wire and_1115_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2470" *)
  wire and_1119_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2469" *)
  wire and_1123_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2468" *)
  wire and_1132_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2467" *)
  wire and_1141_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2466" *)
  wire and_1145_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2465" *)
  wire and_1155_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2464" *)
  wire and_1159_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2463" *)
  wire and_1172_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2462" *)
  wire and_1176_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5477" *)
  wire and_1179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2800" *)
  wire and_1213_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2801" *)
  wire and_1247_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3757" *)
  wire and_1249_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2802" *)
  wire and_1250_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2803" *)
  wire and_1321_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2804" *)
  wire and_1325_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2805" *)
  wire and_1329_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4422" *)
  wire and_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2806" *)
  wire and_1333_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2807" *)
  wire and_1337_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2808" *)
  wire and_1341_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2809" *)
  wire and_1345_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2810" *)
  wire and_1349_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2811" *)
  wire and_1353_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2812" *)
  wire and_1357_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2813" *)
  wire and_1361_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2814" *)
  wire and_1365_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2815" *)
  wire and_1369_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4803" *)
  wire and_136_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2816" *)
  wire and_1373_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2817" *)
  wire and_1377_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2818" *)
  wire and_1381_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2867" *)
  wire and_1385_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2728" *)
  wire and_1386_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4448" *)
  wire and_143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4449" *)
  wire and_145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2868" *)
  wire and_1467_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4462" *)
  wire and_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6608" *)
  wire and_152_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6610" *)
  wire and_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4479" *)
  wire and_156_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4480" *)
  wire and_160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4486" *)
  wire and_161_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4492" *)
  wire and_164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4493" *)
  wire and_166_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6621" *)
  wire and_167_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4517" *)
  wire and_168_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4521" *)
  wire and_171_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4527" *)
  wire and_172_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4543" *)
  wire and_173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3767" *)
  wire and_174_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6634" *)
  wire and_176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3587" *)
  wire and_178_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4567" *)
  wire and_179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4568" *)
  wire and_180_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6640" *)
  wire and_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4585" *)
  wire and_182_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4586" *)
  wire and_183_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6648" *)
  wire and_184_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4599" *)
  wire and_185_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4616" *)
  wire and_194_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4621" *)
  wire and_195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4641" *)
  wire and_199_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4660" *)
  wire and_203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4661" *)
  wire and_205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4685" *)
  wire and_210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4686" *)
  wire and_212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3585" *)
  wire and_2136_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4709" *)
  wire and_213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6824" *)
  wire and_2145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6822" *)
  wire and_2146_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6820" *)
  wire and_2147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6818" *)
  wire and_2148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5145" *)
  wire and_2149_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6816" *)
  wire and_2150_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5105" *)
  wire and_2151_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6814" *)
  wire and_2152_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5025" *)
  wire and_2153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4991" *)
  wire and_2154_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6812" *)
  wire and_2155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4917" *)
  wire and_2156_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6810" *)
  wire and_2157_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6808" *)
  wire and_2158_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4710" *)
  wire and_215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5777" *)
  wire and_2160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5745" *)
  wire and_2161_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5723" *)
  wire and_2162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4740" *)
  wire and_216_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2529" *)
  wire and_2186_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5068" *)
  wire and_2189_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4741" *)
  wire and_218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5055" *)
  wire and_2190_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4848" *)
  wire and_2191_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2570" *)
  wire and_2194_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4771" *)
  wire and_2196_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2569" *)
  wire and_2199_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4768" *)
  wire and_219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4743" *)
  wire and_2201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6699" *)
  wire and_2202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4712" *)
  wire and_2203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2568" *)
  wire and_2206_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6686" *)
  wire and_2208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6680" *)
  wire and_2209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6676" *)
  wire and_2210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4663" *)
  wire and_2213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6669" *)
  wire and_2214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4643" *)
  wire and_2217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6661" *)
  wire and_2218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4769" *)
  wire and_221_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4623" *)
  wire and_2221_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4545" *)
  wire and_2229_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2565" *)
  wire and_2230_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4474" *)
  wire and_2233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4467" *)
  wire and_2234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2562" *)
  wire and_2237_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2554" *)
  wire and_2239_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5453" *)
  wire and_223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4198" *)
  wire and_2240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4200" *)
  wire and_2242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5722" *)
  wire and_2243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3755" *)
  wire and_2246_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6738" *)
  wire and_2247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3530" *)
  wire and_2257_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3768" *)
  wire and_2259_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4536" *)
  wire and_2265_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3518" *)
  wire and_2275_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4821" *)
  wire and_227_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4824" *)
  wire and_228_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4835" *)
  wire and_229_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4838" *)
  wire and_230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3742" *)
  wire and_2317_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4871" *)
  wire and_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4874" *)
  wire and_234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4869" *)
  wire and_2357_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4889" *)
  wire and_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2720" *)
  wire and_2360_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2735" *)
  wire and_2365_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2736" *)
  wire and_2369_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4892" *)
  wire and_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4908" *)
  wire and_2371_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3719" *)
  wire and_2372_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4910" *)
  wire and_237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3747" *)
  wire and_2380_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2741" *)
  wire and_2388_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3772" *)
  wire and_2389_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4913" *)
  wire and_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3773" *)
  wire and_2393_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4989" *)
  wire and_2395_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3494" *)
  wire and_2396_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3495" *)
  wire and_2402_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4933" *)
  wire and_240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4936" *)
  wire and_241_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2742" *)
  wire and_2422_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4967" *)
  wire and_242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4970" *)
  wire and_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4976" *)
  wire and_244_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4979" *)
  wire and_245_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5016" *)
  wire and_247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4737" *)
  wire and_2487_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5019" *)
  wire and_248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5041" *)
  wire and_250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5044" *)
  wire and_251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5096" *)
  wire and_252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5099" *)
  wire and_253_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5122" *)
  wire and_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5125" *)
  wire and_256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5147" *)
  wire and_257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5150" *)
  wire and_258_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5154" *)
  wire and_259_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5157" *)
  wire and_260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5177" *)
  wire and_261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5180" *)
  wire and_262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5460" *)
  wire and_271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5449" *)
  wire and_2780_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5441" *)
  wire and_2782_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5432" *)
  wire and_2784_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5412" *)
  wire and_2786_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5404" *)
  wire and_2788_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5387" *)
  wire and_2789_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5385" *)
  wire and_2791_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5373" *)
  wire and_2793_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5363" *)
  wire and_2795_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5349" *)
  wire and_2797_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5334" *)
  wire and_2799_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5323" *)
  wire and_2801_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5307" *)
  wire and_2803_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5296" *)
  wire and_2805_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5280" *)
  wire and_2807_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5263" *)
  wire and_2809_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5242" *)
  wire and_2811_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3513" *)
  wire and_283_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4610" *)
  wire and_2856_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4456" *)
  wire and_2857_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5462" *)
  wire and_295_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3586" *)
  wire and_3024_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3766" *)
  wire and_3063_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6799" *)
  wire and_306_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4005" *)
  wire and_3104_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4008" *)
  wire and_3105_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4000" *)
  wire and_3109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3993" *)
  wire and_3110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3996" *)
  wire and_3112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3987" *)
  wire and_3115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3978" *)
  wire and_3116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3981" *)
  wire and_3118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3974" *)
  wire and_3121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3968" *)
  wire and_3124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3956" *)
  wire and_3128_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3959" *)
  wire and_3130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3952" *)
  wire and_3133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3946" *)
  wire and_3136_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3935" *)
  wire and_3140_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3928" *)
  wire and_3148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5392" *)
  wire and_3372_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5406" *)
  wire and_3373_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2734" *)
  wire and_550_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2743" *)
  wire and_637_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2744" *)
  wire and_639_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2745" *)
  wire and_641_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2746" *)
  wire and_643_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2747" *)
  wire and_646_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2748" *)
  wire and_648_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2749" *)
  wire and_650_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2750" *)
  wire and_652_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2751" *)
  wire and_654_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2752" *)
  wire and_656_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2753" *)
  wire and_658_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2754" *)
  wire and_660_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2755" *)
  wire and_662_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2756" *)
  wire and_664_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2757" *)
  wire and_666_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2758" *)
  wire and_668_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3502" *)
  wire and_676_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2759" *)
  wire and_685_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4508" *)
  wire and_696_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4509" *)
  wire and_699_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2760" *)
  wire and_704_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4528" *)
  wire and_711_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4529" *)
  wire and_714_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2761" *)
  wire and_719_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4559" *)
  wire and_726_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4560" *)
  wire and_729_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2762" *)
  wire and_734_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4581" *)
  wire and_741_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4582" *)
  wire and_744_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2763" *)
  wire and_749_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4600" *)
  wire and_756_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4601" *)
  wire and_759_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2764" *)
  wire and_766_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4637" *)
  wire and_780_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4638" *)
  wire and_783_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2765" *)
  wire and_787_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4656" *)
  wire and_794_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4657" *)
  wire and_797_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2766" *)
  wire and_801_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4677" *)
  wire and_808_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4678" *)
  wire and_811_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2767" *)
  wire and_816_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4703" *)
  wire and_823_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4704" *)
  wire and_826_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2768" *)
  wire and_830_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4730" *)
  wire and_840_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4731" *)
  wire and_843_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2769" *)
  wire and_849_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4757" *)
  wire and_856_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4758" *)
  wire and_859_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2770" *)
  wire and_866_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4786" *)
  wire and_873_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4787" *)
  wire and_876_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2771" *)
  wire and_881_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2772" *)
  wire and_896_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2773" *)
  wire and_900_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5471" *)
  wire and_908_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4861" *)
  wire and_916_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4862" *)
  wire and_921_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4905" *)
  wire and_945_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4906" *)
  wire and_949_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2774" *)
  wire and_954_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2775" *)
  wire and_956_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2776" *)
  wire and_957_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4959" *)
  wire and_961_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4960" *)
  wire and_966_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3493" *)
  wire and_976_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3506" *)
  wire and_978_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2777" *)
  wire and_984_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2778" *)
  wire and_986_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2779" *)
  wire and_987_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2780" *)
  wire and_989_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4189" *)
  wire and_98_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5087" *)
  wire and_999_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1368" *)
  wire and_dcpl_1003;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1242" *)
  wire and_dcpl_102;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1243" *)
  wire and_dcpl_103;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1244" *)
  wire and_dcpl_105;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1245" *)
  wire and_dcpl_114;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2787" *)
  wire and_dcpl_1319;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3534" *)
  wire and_dcpl_1742;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1250" *)
  wire and_dcpl_204;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1251" *)
  wire and_dcpl_209;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1252" *)
  wire and_dcpl_217;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1253" *)
  wire and_dcpl_224;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1255" *)
  wire and_dcpl_228;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:998" *)
  wire and_dcpl_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1269" *)
  wire and_dcpl_301;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1281" *)
  wire and_dcpl_363;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:999" *)
  wire and_dcpl_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1288" *)
  wire and_dcpl_401;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1289" *)
  wire and_dcpl_407;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1290" *)
  wire and_dcpl_408;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1292" *)
  wire and_dcpl_409;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1293" *)
  wire and_dcpl_411;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1294" *)
  wire and_dcpl_417;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1295" *)
  wire and_dcpl_420;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1296" *)
  wire and_dcpl_424;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1297" *)
  wire and_dcpl_425;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1298" *)
  wire and_dcpl_433;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1300" *)
  wire and_dcpl_444;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1301" *)
  wire and_dcpl_446;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1303" *)
  wire and_dcpl_458;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1306" *)
  wire and_dcpl_473;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1307" *)
  wire and_dcpl_479;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1309" *)
  wire and_dcpl_481;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1311" *)
  wire and_dcpl_499;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1313" *)
  wire and_dcpl_535;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1320" *)
  wire and_dcpl_617;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1321" *)
  wire and_dcpl_626;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1323" *)
  wire and_dcpl_631;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1324" *)
  wire and_dcpl_648;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1000" *)
  wire and_dcpl_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1002" *)
  wire and_dcpl_73;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1239" *)
  wire and_dcpl_93;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1346" *)
  wire and_dcpl_942;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1348" *)
  wire and_dcpl_946;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1349" *)
  wire and_dcpl_950;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1351" *)
  wire and_dcpl_954;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1352" *)
  wire and_dcpl_958;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1354" *)
  wire and_dcpl_962;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1356" *)
  wire and_dcpl_966;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1357" *)
  wire and_dcpl_970;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1358" *)
  wire and_dcpl_974;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1360" *)
  wire and_dcpl_978;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1241" *)
  wire and_dcpl_98;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1362" *)
  wire and_dcpl_982;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1363" *)
  wire and_dcpl_987;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1365" *)
  wire and_dcpl_991;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1366" *)
  wire and_dcpl_995;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1367" *)
  wire and_dcpl_999;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5744" *)
  wire and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1012" *)
  wire and_tmp_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1014" *)
  wire and_tmp_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1016" *)
  wire and_tmp_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1147" *)
  wire and_tmp_165;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1150" *)
  wire and_tmp_166;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1153" *)
  wire and_tmp_168;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1156" *)
  wire and_tmp_169;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1165" *)
  wire and_tmp_171;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1176" *)
  wire and_tmp_175;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1021" *)
  wire and_tmp_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1024" *)
  wire and_tmp_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1264" *)
  wire and_tmp_225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1304" *)
  wire and_tmp_248;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1026" *)
  wire and_tmp_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1038" *)
  wire and_tmp_50;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1039" *)
  wire and_tmp_52;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1048" *)
  wire and_tmp_67;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1060" *)
  wire and_tmp_71;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1067" *)
  wire and_tmp_79;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1011" *)
  wire and_tmp_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1082" *)
  wire and_tmp_93;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1084" *)
  wire and_tmp_94;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1685" *)
  reg cfg_mode_eql_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1686" *)
  reg cfg_mode_eql_1_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1687" *)
  reg cfg_mode_eql_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:699" *)
  input cfg_mode_eql_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:720" *)
  wire cfg_mode_eql_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:694" *)
  input [31:0] cfg_offset_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:715" *)
  wire [31:0] cfg_offset_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1684" *)
  reg [1:0] cfg_out_precision_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2053" *)
  reg [1:0] cfg_out_precision_1_sva_st_113;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2088" *)
  reg [1:0] cfg_out_precision_1_sva_st_136;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2105" *)
  reg [1:0] cfg_out_precision_1_sva_st_144;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2109" *)
  reg [1:0] cfg_out_precision_1_sva_st_149;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2111" *)
  reg [1:0] cfg_out_precision_1_sva_st_154;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2112" *)
  reg [1:0] cfg_out_precision_1_sva_st_156;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3476" *)
  wire cfg_out_precision_and_32_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:698" *)
  input [1:0] cfg_out_precision_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:719" *)
  wire [1:0] cfg_out_precision_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2107" *)
  reg [1:0] cfg_proc_precision_1_sva_st_101;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2108" *)
  reg [1:0] cfg_proc_precision_1_sva_st_102;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2110" *)
  reg [1:0] cfg_proc_precision_1_sva_st_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2035" *)
  reg [1:0] cfg_proc_precision_1_sva_st_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2039" *)
  reg [1:0] cfg_proc_precision_1_sva_st_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2040" *)
  reg [1:0] cfg_proc_precision_1_sva_st_66;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2102" *)
  reg [1:0] cfg_proc_precision_1_sva_st_89;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2103" *)
  reg [1:0] cfg_proc_precision_1_sva_st_90;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3451" *)
  wire cfg_proc_precision_and_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3458" *)
  wire cfg_proc_precision_and_24_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3459" *)
  wire cfg_proc_precision_and_27_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3474" *)
  wire cfg_proc_precision_and_40_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3475" *)
  wire cfg_proc_precision_and_43_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:697" *)
  input [1:0] cfg_proc_precision_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:718" *)
  wire [1:0] cfg_proc_precision_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:695" *)
  input [15:0] cfg_scale_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:716" *)
  wire [15:0] cfg_scale_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1683" *)
  reg [5:0] cfg_truncate_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:696" *)
  input [5:0] cfg_truncate_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:717" *)
  wire [5:0] cfg_truncate_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3452" *)
  wire chn_idata_data_and_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3448" *)
  wire chn_idata_data_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2630" *)
  wire [15:0] chn_idata_data_mux1h_65_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2158" *)
  reg [28:0] chn_idata_data_sva_1_123_95_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2157" *)
  reg [28:0] chn_idata_data_sva_1_155_127_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2156" *)
  reg [28:0] chn_idata_data_sva_1_187_159_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2155" *)
  reg [28:0] chn_idata_data_sva_1_219_191_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2154" *)
  reg [28:0] chn_idata_data_sva_1_251_223_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2161" *)
  reg [27:0] chn_idata_data_sva_1_27_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2153" *)
  reg [28:0] chn_idata_data_sva_1_283_255_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2152" *)
  reg [28:0] chn_idata_data_sva_1_315_287_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2151" *)
  reg [28:0] chn_idata_data_sva_1_347_319_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2150" *)
  reg [28:0] chn_idata_data_sva_1_379_351_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2149" *)
  reg [28:0] chn_idata_data_sva_1_411_383_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2148" *)
  reg [28:0] chn_idata_data_sva_1_443_415_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2147" *)
  reg [28:0] chn_idata_data_sva_1_475_447_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2146" *)
  reg [28:0] chn_idata_data_sva_1_507_479_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2145" *)
  reg chn_idata_data_sva_1_511_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2160" *)
  reg [28:0] chn_idata_data_sva_1_59_31_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2159" *)
  reg [28:0] chn_idata_data_sva_1_91_63_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2175" *)
  reg [16:0] chn_idata_data_sva_2_111_95_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2174" *)
  reg [16:0] chn_idata_data_sva_2_143_127_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2178" *)
  reg [15:0] chn_idata_data_sva_2_15_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2173" *)
  reg [16:0] chn_idata_data_sva_2_175_159_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2172" *)
  reg [16:0] chn_idata_data_sva_2_207_191_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2171" *)
  reg [16:0] chn_idata_data_sva_2_239_223_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2170" *)
  reg [16:0] chn_idata_data_sva_2_271_255_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2169" *)
  reg [16:0] chn_idata_data_sva_2_303_287_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2168" *)
  reg [16:0] chn_idata_data_sva_2_335_319_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2167" *)
  reg [16:0] chn_idata_data_sva_2_367_351_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2166" *)
  reg [16:0] chn_idata_data_sva_2_399_383_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2165" *)
  reg [16:0] chn_idata_data_sva_2_431_415_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2164" *)
  reg [16:0] chn_idata_data_sva_2_463_447_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2177" *)
  reg [16:0] chn_idata_data_sva_2_47_31_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2163" *)
  reg [16:0] chn_idata_data_sva_2_495_479_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2162" *)
  reg chn_idata_data_sva_2_511_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2176" *)
  reg [16:0] chn_idata_data_sva_2_79_63_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2191" *)
  reg [16:0] chn_idata_data_sva_3_111_95_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2190" *)
  reg [16:0] chn_idata_data_sva_3_143_127_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2189" *)
  reg [16:0] chn_idata_data_sva_3_175_159_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2188" *)
  reg [16:0] chn_idata_data_sva_3_207_191_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2187" *)
  reg [16:0] chn_idata_data_sva_3_239_223_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2186" *)
  reg [16:0] chn_idata_data_sva_3_271_255_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2185" *)
  reg [16:0] chn_idata_data_sva_3_303_287_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2184" *)
  reg [16:0] chn_idata_data_sva_3_335_319_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2183" *)
  reg [16:0] chn_idata_data_sva_3_367_351_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2182" *)
  reg [16:0] chn_idata_data_sva_3_399_383_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2181" *)
  reg [16:0] chn_idata_data_sva_3_431_415_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2180" *)
  reg [16:0] chn_idata_data_sva_3_463_447_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2193" *)
  reg [16:0] chn_idata_data_sva_3_47_31_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2179" *)
  reg [16:0] chn_idata_data_sva_3_495_479_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2192" *)
  reg [16:0] chn_idata_data_sva_3_79_63_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:693" *)
  output chn_in_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:692" *)
  input chn_in_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:691" *)
  input [511:0] chn_in_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:710" *)
  wire chn_in_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:713" *)
  wire [511:0] chn_in_rsci_d_mxwt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:709" *)
  reg chn_in_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:712" *)
  reg chn_in_rsci_ld_core_psct;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2935" *)
  wire chn_in_rsci_ld_core_psct_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:703" *)
  input chn_in_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:704" *)
  output chn_in_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:711" *)
  wire chn_in_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1481" *)
  reg chn_odata_data_13_0_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3064" *)
  wire chn_odata_data_13_0_lpi_1_dfm_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4160" *)
  wire chn_odata_data_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2492" *)
  wire chn_out_and_32_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2493" *)
  wire chn_out_and_77_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2479" *)
  wire chn_out_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:702" *)
  output chn_out_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:701" *)
  input chn_out_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:700" *)
  output [271:0] chn_out_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:722" *)
  wire chn_out_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:787" *)
  reg chn_out_rsci_d_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:768" *)
  reg [8:0] chn_out_rsci_d_105_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:807" *)
  reg [3:0] chn_out_rsci_d_109_106;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:806" *)
  reg chn_out_rsci_d_110;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:767" *)
  reg chn_out_rsci_d_111;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:766" *)
  reg chn_out_rsci_d_112;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:765" *)
  reg [8:0] chn_out_rsci_d_121_113;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:805" *)
  reg [3:0] chn_out_rsci_d_125_122;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:804" *)
  reg chn_out_rsci_d_126;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:764" *)
  reg chn_out_rsci_d_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:763" *)
  reg chn_out_rsci_d_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:762" *)
  reg [8:0] chn_out_rsci_d_137_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:819" *)
  reg [3:0] chn_out_rsci_d_13_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:818" *)
  reg chn_out_rsci_d_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:803" *)
  reg [3:0] chn_out_rsci_d_141_138;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:802" *)
  reg chn_out_rsci_d_142;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:761" *)
  reg chn_out_rsci_d_143;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:760" *)
  reg chn_out_rsci_d_144;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:785" *)
  reg chn_out_rsci_d_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:759" *)
  reg [8:0] chn_out_rsci_d_153_145;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:801" *)
  reg [3:0] chn_out_rsci_d_157_154;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:800" *)
  reg chn_out_rsci_d_158;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:758" *)
  reg chn_out_rsci_d_159;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:784" *)
  reg chn_out_rsci_d_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:757" *)
  reg chn_out_rsci_d_160;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:756" *)
  reg [8:0] chn_out_rsci_d_169_161;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:799" *)
  reg [3:0] chn_out_rsci_d_173_170;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:798" *)
  reg chn_out_rsci_d_174;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:755" *)
  reg chn_out_rsci_d_175;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:754" *)
  reg chn_out_rsci_d_176;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:753" *)
  reg [8:0] chn_out_rsci_d_185_177;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:797" *)
  reg [3:0] chn_out_rsci_d_189_186;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:796" *)
  reg chn_out_rsci_d_190;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:752" *)
  reg chn_out_rsci_d_191;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:751" *)
  reg chn_out_rsci_d_192;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:750" *)
  reg [8:0] chn_out_rsci_d_201_193;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:795" *)
  reg [3:0] chn_out_rsci_d_205_202;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:794" *)
  reg chn_out_rsci_d_206;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:749" *)
  reg chn_out_rsci_d_207;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:748" *)
  reg chn_out_rsci_d_208;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:747" *)
  reg [8:0] chn_out_rsci_d_217_209;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:793" *)
  reg [3:0] chn_out_rsci_d_221_218;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:792" *)
  reg chn_out_rsci_d_222;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:746" *)
  reg chn_out_rsci_d_223;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:745" *)
  reg chn_out_rsci_d_224;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:744" *)
  reg [8:0] chn_out_rsci_d_233_225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:791" *)
  reg [3:0] chn_out_rsci_d_237_234;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:790" *)
  reg chn_out_rsci_d_238;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:743" *)
  reg chn_out_rsci_d_239;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:742" *)
  reg chn_out_rsci_d_240;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:741" *)
  reg [8:0] chn_out_rsci_d_249_241;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:789" *)
  reg [3:0] chn_out_rsci_d_253_250;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:788" *)
  reg chn_out_rsci_d_254;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:740" *)
  reg chn_out_rsci_d_255;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:739" *)
  reg chn_out_rsci_d_256;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:738" *)
  reg chn_out_rsci_d_257;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:737" *)
  reg chn_out_rsci_d_258;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:736" *)
  reg chn_out_rsci_d_259;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:783" *)
  reg [8:0] chn_out_rsci_d_25_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:735" *)
  reg chn_out_rsci_d_260;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:734" *)
  reg chn_out_rsci_d_261;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:733" *)
  reg chn_out_rsci_d_262;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:732" *)
  reg chn_out_rsci_d_263;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:731" *)
  reg chn_out_rsci_d_264;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:730" *)
  reg chn_out_rsci_d_265;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:729" *)
  reg chn_out_rsci_d_266;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:728" *)
  reg chn_out_rsci_d_267;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:727" *)
  reg chn_out_rsci_d_268;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:726" *)
  reg chn_out_rsci_d_269;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:725" *)
  reg chn_out_rsci_d_270;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:724" *)
  reg chn_out_rsci_d_271;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:817" *)
  reg [3:0] chn_out_rsci_d_29_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:816" *)
  reg chn_out_rsci_d_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:782" *)
  reg chn_out_rsci_d_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:781" *)
  reg chn_out_rsci_d_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:780" *)
  reg [8:0] chn_out_rsci_d_41_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:815" *)
  reg [3:0] chn_out_rsci_d_45_42;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:814" *)
  reg chn_out_rsci_d_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:779" *)
  reg chn_out_rsci_d_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:778" *)
  reg chn_out_rsci_d_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:777" *)
  reg [8:0] chn_out_rsci_d_57_49;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:813" *)
  reg [3:0] chn_out_rsci_d_61_58;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:812" *)
  reg chn_out_rsci_d_62;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:776" *)
  reg chn_out_rsci_d_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:775" *)
  reg chn_out_rsci_d_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:774" *)
  reg [8:0] chn_out_rsci_d_73_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:811" *)
  reg [3:0] chn_out_rsci_d_77_74;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:810" *)
  reg chn_out_rsci_d_78;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:773" *)
  reg chn_out_rsci_d_79;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:772" *)
  reg chn_out_rsci_d_80;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:771" *)
  reg [8:0] chn_out_rsci_d_89_81;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:809" *)
  reg [3:0] chn_out_rsci_d_93_90;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:808" *)
  reg chn_out_rsci_d_94;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:770" *)
  reg chn_out_rsci_d_95;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:769" *)
  reg chn_out_rsci_d_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:786" *)
  reg [8:0] chn_out_rsci_d_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:721" *)
  reg chn_out_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:705" *)
  input chn_out_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:706" *)
  output chn_out_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:723" *)
  wire chn_out_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:708" *)
  wire core_wen;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:714" *)
  wire core_wten;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6203" *)
  wire cvt_10_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2015" *)
  reg cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3059" *)
  wire cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3060" *)
  wire cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3654" *)
  wire cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6201" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1543" *)
  reg cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1945" *)
  reg [4:0] cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1444" *)
  reg cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1860" *)
  reg cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:867" *)
  wire cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6426" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3788" *)
  wire cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5368" *)
  wire [4:0] cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3425" *)
  wire cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1977" *)
  reg cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2793" *)
  wire [16:0] cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6531" *)
  wire cvt_10_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2926" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6532" *)
  wire [22:0] cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6238" *)
  wire [9:0] cvt_10_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1446" *)
  reg cvt_10_FpMantRNE_17U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:923" *)
  wire cvt_10_FpMantRNE_17U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6074" *)
  wire [9:0] cvt_10_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1380" *)
  reg cvt_10_FpMantRNE_24U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1748" *)
  reg cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:827" *)
  wire cvt_10_FpMantRNE_24U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3626" *)
  wire cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5971" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3606" *)
  wire cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5931" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:968" *)
  wire [4:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1653" *)
  reg cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2068" *)
  reg cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3607" *)
  wire cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5933" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2066" *)
  reg cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4406" *)
  wire [48:0] cvt_10_IntMulExt_33U_16U_49U_o_mul_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3702" *)
  wire cvt_10_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6570" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3665" *)
  wire cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6353" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_10_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3686" *)
  wire cvt_10_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6476" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4806" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_10_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1993" *)
  reg cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:939" *)
  wire cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5513" *)
  wire [17:0] cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6310" *)
  wire [17:0] cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:870" *)
  wire [49:0] cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6355" *)
  wire cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:868" *)
  wire cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:869" *)
  wire cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6144" *)
  wire [14:0] cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2586" *)
  wire cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6394" *)
  wire cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6395" *)
  wire [23:0] cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4407" *)
  wire [32:0] cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6206" *)
  wire cvt_11_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2013" *)
  reg cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3062" *)
  wire cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3063" *)
  wire cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3655" *)
  wire cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6204" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1520" *)
  reg cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1948" *)
  reg [4:0] cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1452" *)
  reg cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1868" *)
  reg cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:862" *)
  wire cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6428" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3789" *)
  wire cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5380" *)
  wire [4:0] cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3426" *)
  wire cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1978" *)
  reg cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2794" *)
  wire [16:0] cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6534" *)
  wire cvt_11_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2927" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6535" *)
  wire [22:0] cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6244" *)
  wire [9:0] cvt_11_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1454" *)
  reg cvt_11_FpMantRNE_17U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:922" *)
  wire cvt_11_FpMantRNE_17U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6083" *)
  wire [9:0] cvt_11_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1381" *)
  reg cvt_11_FpMantRNE_24U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1754" *)
  reg cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:826" *)
  wire cvt_11_FpMantRNE_24U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3625" *)
  wire cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5969" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3608" *)
  wire cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5935" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:965" *)
  wire [4:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1650" *)
  reg cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2071" *)
  reg cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3609" *)
  wire cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5937" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2069" *)
  reg cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4412" *)
  wire [48:0] cvt_11_IntMulExt_33U_16U_49U_o_mul_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3703" *)
  wire cvt_11_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6572" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3666" *)
  wire cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6356" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_11_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3687" *)
  wire cvt_11_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6480" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5183" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_11_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1992" *)
  reg cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:938" *)
  wire cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5510" *)
  wire [17:0] cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6314" *)
  wire [17:0] cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:865" *)
  wire [49:0] cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6361" *)
  wire cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:863" *)
  wire cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:864" *)
  wire cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6145" *)
  wire [14:0] cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2587" *)
  wire cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6396" *)
  wire cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6397" *)
  wire [23:0] cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4413" *)
  wire [32:0] cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6200" *)
  wire cvt_12_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2011" *)
  reg cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3056" *)
  wire cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3057" *)
  wire cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3653" *)
  wire cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6198" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1540" *)
  reg cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1951" *)
  reg [4:0] cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1460" *)
  reg cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1876" *)
  reg cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:857" *)
  wire cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6430" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3790" *)
  wire cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5399" *)
  wire [4:0] cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3427" *)
  wire cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1979" *)
  reg cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2795" *)
  wire [16:0] cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6537" *)
  wire cvt_12_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2928" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6538" *)
  wire [22:0] cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6250" *)
  wire [9:0] cvt_12_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1462" *)
  reg cvt_12_FpMantRNE_17U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:921" *)
  wire cvt_12_FpMantRNE_17U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6092" *)
  wire [9:0] cvt_12_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1382" *)
  reg cvt_12_FpMantRNE_24U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1760" *)
  reg cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:825" *)
  wire cvt_12_FpMantRNE_24U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3624" *)
  wire cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5967" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3610" *)
  wire cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5939" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:962" *)
  wire [4:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1647" *)
  reg cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2074" *)
  reg cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3611" *)
  wire cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5941" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2072" *)
  reg cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4409" *)
  wire [48:0] cvt_12_IntMulExt_33U_16U_49U_o_mul_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3704" *)
  wire cvt_12_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6574" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3667" *)
  wire cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6358" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_12_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3688" *)
  wire cvt_12_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6484" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5190" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_12_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1991" *)
  reg cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:937" *)
  wire cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5507" *)
  wire [17:0] cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6312" *)
  wire [17:0] cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:860" *)
  wire [49:0] cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6360" *)
  wire cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:858" *)
  wire cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:859" *)
  wire cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6146" *)
  wire [14:0] cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2588" *)
  wire cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6398" *)
  wire cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6399" *)
  wire [23:0] cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4410" *)
  wire [32:0] cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6192" *)
  wire cvt_13_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2009" *)
  reg cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3050" *)
  wire cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3051" *)
  wire cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3650" *)
  wire cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6190" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1525" *)
  reg cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1954" *)
  reg [4:0] cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1470" *)
  reg cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1884" *)
  reg cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:852" *)
  wire cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6432" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3791" *)
  wire cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5407" *)
  wire [4:0] cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3428" *)
  wire cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1980" *)
  reg cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2796" *)
  wire [16:0] cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6540" *)
  wire cvt_13_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2929" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6541" *)
  wire [22:0] cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6256" *)
  wire [9:0] cvt_13_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1472" *)
  reg cvt_13_FpMantRNE_17U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:920" *)
  wire cvt_13_FpMantRNE_17U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6101" *)
  wire [9:0] cvt_13_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1383" *)
  reg cvt_13_FpMantRNE_24U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1766" *)
  reg cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:824" *)
  wire cvt_13_FpMantRNE_24U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3623" *)
  wire cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5965" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3612" *)
  wire cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5943" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:959" *)
  wire [4:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1644" *)
  reg cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2077" *)
  reg cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3613" *)
  wire cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5945" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2075" *)
  reg cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4428" *)
  wire [48:0] cvt_13_IntMulExt_33U_16U_49U_o_mul_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3705" *)
  wire cvt_13_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6576" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3668" *)
  wire cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6362" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_13_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3689" *)
  wire cvt_13_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6488" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5169" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_13_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1990" *)
  reg cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:936" *)
  wire cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5504" *)
  wire [17:0] cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6322" *)
  wire [17:0] cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:855" *)
  wire [49:0] cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6373" *)
  wire cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:853" *)
  wire cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:854" *)
  wire cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6147" *)
  wire [14:0] cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2589" *)
  wire cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6400" *)
  wire cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6401" *)
  wire [23:0] cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4429" *)
  wire [32:0] cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6186" *)
  wire cvt_14_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2007" *)
  reg cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3046" *)
  wire cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3047" *)
  wire cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3648" *)
  wire cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6184" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1530" *)
  reg cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1957" *)
  reg [4:0] cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1477" *)
  reg cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1892" *)
  reg cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:847" *)
  wire cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6434" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3792" *)
  wire cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5427" *)
  wire [4:0] cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3429" *)
  wire cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1981" *)
  reg cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2797" *)
  wire [16:0] cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6543" *)
  wire cvt_14_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2930" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6544" *)
  wire [22:0] cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6262" *)
  wire [9:0] cvt_14_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1479" *)
  reg cvt_14_FpMantRNE_17U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:919" *)
  wire cvt_14_FpMantRNE_17U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6110" *)
  wire [9:0] cvt_14_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1384" *)
  reg cvt_14_FpMantRNE_24U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1772" *)
  reg cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:823" *)
  wire cvt_14_FpMantRNE_24U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3622" *)
  wire cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5963" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3614" *)
  wire cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5947" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:956" *)
  wire [4:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1641" *)
  reg cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2080" *)
  reg cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3615" *)
  wire cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5949" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2078" *)
  reg cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4415" *)
  wire [48:0] cvt_14_IntMulExt_33U_16U_49U_o_mul_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3708" *)
  wire cvt_14_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6582" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3669" *)
  wire cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6364" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_14_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3692" *)
  wire cvt_14_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6502" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5415" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_14_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1587" *)
  reg cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1989" *)
  reg cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:935" *)
  wire cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5501" *)
  wire [17:0] cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire [8:0] cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:850" *)
  wire [49:0] cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6366" *)
  wire cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:848" *)
  wire cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:849" *)
  wire cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6148" *)
  wire [14:0] cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2590" *)
  wire cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6402" *)
  wire cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6403" *)
  wire [23:0] cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4416" *)
  wire [32:0] cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6180" *)
  wire cvt_15_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2006" *)
  reg cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3646" *)
  wire cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6178" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1535" *)
  reg cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1960" *)
  reg [4:0] cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1485" *)
  reg cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1900" *)
  reg cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:842" *)
  wire cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6436" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3793" *)
  wire cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5436" *)
  wire [4:0] cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3430" *)
  wire cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1985" *)
  reg cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2798" *)
  wire [16:0] cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6546" *)
  wire cvt_15_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2931" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6547" *)
  wire [22:0] cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6268" *)
  wire [9:0] cvt_15_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1487" *)
  reg cvt_15_FpMantRNE_17U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:918" *)
  wire cvt_15_FpMantRNE_17U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6119" *)
  wire [9:0] cvt_15_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1385" *)
  reg cvt_15_FpMantRNE_24U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1778" *)
  reg cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:822" *)
  wire cvt_15_FpMantRNE_24U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3621" *)
  wire cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5961" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3616" *)
  wire cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5951" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:953" *)
  wire [4:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1638" *)
  reg cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2083" *)
  reg cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3617" *)
  wire cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5953" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2081" *)
  reg cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4425" *)
  wire [48:0] cvt_15_IntMulExt_33U_16U_49U_o_mul_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3706" *)
  wire cvt_15_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6578" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3670" *)
  wire cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6367" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_15_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3690" *)
  wire cvt_15_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6494" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5134" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_15_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1988" *)
  reg cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:934" *)
  wire cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5498" *)
  wire [17:0] cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6320" *)
  wire [17:0] cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:845" *)
  wire [49:0] cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6372" *)
  wire cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:843" *)
  wire cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:844" *)
  wire cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6149" *)
  wire [14:0] cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2591" *)
  wire cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6404" *)
  wire cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6405" *)
  wire [23:0] cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4426" *)
  wire [32:0] cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6172" *)
  wire cvt_16_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2004" *)
  reg cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3038" *)
  wire cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3039" *)
  wire cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3643" *)
  wire cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6170" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1533" *)
  reg cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1965" *)
  reg [4:0] cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1492" *)
  reg cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1908" *)
  reg cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:837" *)
  wire cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6438" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3794" *)
  wire cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5444" *)
  wire [4:0] cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3431" *)
  wire cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1986" *)
  reg cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2799" *)
  wire [16:0] cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6549" *)
  wire cvt_16_FpMantDecShiftRight_23U_8U_10U_carry_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2932" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6550" *)
  wire [22:0] cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6274" *)
  wire [9:0] cvt_16_FpMantRNE_17U_11U_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1494" *)
  reg cvt_16_FpMantRNE_17U_11U_else_and_4_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:917" *)
  wire cvt_16_FpMantRNE_17U_11U_else_and_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6128" *)
  wire [9:0] cvt_16_FpMantRNE_24U_11U_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1386" *)
  reg cvt_16_FpMantRNE_24U_11U_else_and_4_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1784" *)
  reg cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:821" *)
  wire cvt_16_FpMantRNE_24U_11U_else_and_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3620" *)
  wire cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5959" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3618" *)
  wire cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5955" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:950" *)
  wire [4:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1635" *)
  reg cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2086" *)
  reg cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3619" *)
  wire cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5957" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2084" *)
  reg cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4418" *)
  wire [48:0] cvt_16_IntMulExt_33U_16U_49U_o_mul_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3707" *)
  wire cvt_16_IntSaturation_17U_16U_else_if_acc_4_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6580" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3671" *)
  wire cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6369" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_16_IntSaturation_17U_16U_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3691" *)
  wire cvt_16_IntSaturation_17U_8U_else_if_acc_4_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6498" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5065" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_16_IntSaturation_17U_8U_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1987" *)
  reg cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:933" *)
  wire cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5463" *)
  wire [17:0] cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6318" *)
  wire [17:0] cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:840" *)
  wire [49:0] cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6371" *)
  wire cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:838" *)
  wire cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:839" *)
  wire cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6150" *)
  wire [14:0] cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2592" *)
  wire cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_24_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6406" *)
  wire cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6407" *)
  wire [23:0] cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4419" *)
  wire [32:0] cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6153" *)
  wire cvt_1_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2034" *)
  reg cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3636" *)
  wire cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6151" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1503" *)
  reg cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1912" *)
  reg [4:0] cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2087" *)
  reg cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:912" *)
  wire cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3672" *)
  wire cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6408" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5237" *)
  wire [4:0] cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3416" *)
  wire cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1967" *)
  reg cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6504" *)
  wire cvt_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2917" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6505" *)
  wire [22:0] cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5474" *)
  wire [9:0] cvt_1_FpMantRNE_17U_11U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1390" *)
  reg cvt_1_FpMantRNE_17U_11U_else_and_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:932" *)
  wire cvt_1_FpMantRNE_17U_11U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5993" *)
  wire [9:0] cvt_1_FpMantRNE_24U_11U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1371" *)
  reg cvt_1_FpMantRNE_24U_11U_else_and_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1695" *)
  reg cvt_1_FpMantRNE_24U_11U_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:836" *)
  wire cvt_1_FpMantRNE_24U_11U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3635" *)
  wire cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5989" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3588" *)
  wire cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5895" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:996" *)
  wire [4:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1681" *)
  reg cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2038" *)
  reg cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3589" *)
  wire cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5897" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2036" *)
  reg cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3693" *)
  wire cvt_1_IntSaturation_17U_16U_else_if_acc_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6552" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_1_IntSaturation_17U_16U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3656" *)
  wire cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6328" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_1_IntSaturation_17U_16U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3677" *)
  wire cvt_1_IntSaturation_17U_8U_else_if_acc_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6440" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_1_IntSaturation_17U_8U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3645" *)
  wire cvt_1_IntSaturation_17U_8U_if_acc_itm_10_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6176" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_1_IntSaturation_17U_8U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2089" *)
  reg cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2002" *)
  reg cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1789" *)
  reg cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:948" *)
  wire cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5540" *)
  wire [17:0] cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6326" *)
  wire [17:0] cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:915" *)
  wire [49:0] cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:913" *)
  wire cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6375" *)
  wire cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6135" *)
  wire [14:0] cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2577" *)
  wire cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:914" *)
  wire cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6376" *)
  wire cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6377" *)
  wire [23:0] cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4433" *)
  wire [32:0] cvt_1_IntSubExt_32U_32U_33U_o_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6156" *)
  wire cvt_2_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2032" *)
  reg cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3026" *)
  wire cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3027" *)
  wire cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3637" *)
  wire cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6154" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1506" *)
  reg cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1917" *)
  reg [4:0] cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1798" *)
  reg cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2091" *)
  reg cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:907" *)
  wire cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3673" *)
  wire cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6410" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5258" *)
  wire [4:0] cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3417" *)
  wire cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1968" *)
  reg cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6507" *)
  wire cvt_2_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2918" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6508" *)
  wire [22:0] cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4854" *)
  wire [9:0] cvt_2_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1395" *)
  reg cvt_2_FpMantRNE_17U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:931" *)
  wire cvt_2_FpMantRNE_17U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6002" *)
  wire [9:0] cvt_2_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1372" *)
  reg cvt_2_FpMantRNE_24U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1701" *)
  reg cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:835" *)
  wire cvt_2_FpMantRNE_24U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3634" *)
  wire cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5987" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3590" *)
  wire cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5899" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:993" *)
  wire [4:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1678" *)
  reg cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2043" *)
  reg cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3591" *)
  wire cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5901" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2041" *)
  reg cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3694" *)
  wire cvt_2_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6554" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3657" *)
  wire cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6330" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_2_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3678" *)
  wire cvt_2_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6444" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4832" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_2_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2001" *)
  reg cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2090" *)
  reg cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:947" *)
  wire cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5537" *)
  wire [17:0] cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6296" *)
  wire [17:0] cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:910" *)
  wire [49:0] cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6332" *)
  wire cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:908" *)
  wire cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:909" *)
  wire cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6136" *)
  wire [14:0] cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2578" *)
  wire cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6378" *)
  wire cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6379" *)
  wire [23:0] cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4388" *)
  wire [32:0] cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2937" *)
  wire cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6161" *)
  wire cvt_3_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2029" *)
  reg cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3029" *)
  wire cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3030" *)
  wire cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3639" *)
  wire cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6159" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1559" *)
  reg cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1922" *)
  reg [4:0] cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1805" *)
  reg cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2093" *)
  reg cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:902" *)
  wire cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3674" *)
  wire cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6412" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5275" *)
  wire [4:0] cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3418" *)
  wire cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1969" *)
  reg cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2784" *)
  wire [16:0] cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6510" *)
  wire cvt_3_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2919" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6511" *)
  wire [22:0] cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5267" *)
  wire [9:0] cvt_3_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1401" *)
  reg cvt_3_FpMantRNE_17U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:930" *)
  wire cvt_3_FpMantRNE_17U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6011" *)
  wire [9:0] cvt_3_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1373" *)
  reg cvt_3_FpMantRNE_24U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1707" *)
  reg cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:834" *)
  wire cvt_3_FpMantRNE_24U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3633" *)
  wire cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5985" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3592" *)
  wire cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5903" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:990" *)
  wire [4:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1675" *)
  reg cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2046" *)
  reg cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3593" *)
  wire cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5905" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2044" *)
  reg cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3695" *)
  wire cvt_3_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6556" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3658" *)
  wire cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6333" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_3_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3679" *)
  wire cvt_3_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6448" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3638" *)
  wire cvt_3_IntSaturation_17U_8U_if_acc_1_itm_10_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6157" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_3_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2094" *)
  reg cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2000" *)
  reg cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2092" *)
  reg cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:946" *)
  wire cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5534" *)
  wire [17:0] cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6300" *)
  wire [17:0] cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:905" *)
  wire [49:0] cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6338" *)
  wire cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:903" *)
  wire cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:904" *)
  wire cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6137" *)
  wire [14:0] cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2579" *)
  wire cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6380" *)
  wire cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6381" *)
  wire [23:0] cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4393" *)
  wire [32:0] cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6164" *)
  wire cvt_4_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2027" *)
  reg cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3032" *)
  wire cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3033" *)
  wire cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3640" *)
  wire cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6162" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1509" *)
  reg cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1925" *)
  reg [4:0] cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1405" *)
  reg cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1814" *)
  reg cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:897" *)
  wire cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6414" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3784" *)
  wire cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5291" *)
  wire [4:0] cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3419" *)
  wire cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1971" *)
  reg cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2786" *)
  wire [16:0] cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6513" *)
  wire cvt_4_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2920" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6514" *)
  wire [22:0] cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6211" *)
  wire [9:0] cvt_4_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1407" *)
  reg cvt_4_FpMantRNE_17U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:929" *)
  wire cvt_4_FpMantRNE_17U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6020" *)
  wire [9:0] cvt_4_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1374" *)
  reg cvt_4_FpMantRNE_24U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1713" *)
  reg cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:833" *)
  wire cvt_4_FpMantRNE_24U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3632" *)
  wire cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5983" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3594" *)
  wire cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5907" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:987" *)
  wire [4:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1672" *)
  reg cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2049" *)
  reg cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3595" *)
  wire cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5909" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2047" *)
  reg cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4390" *)
  wire [48:0] cvt_4_IntMulExt_33U_16U_49U_o_mul_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3696" *)
  wire cvt_4_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6558" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3659" *)
  wire cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6335" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_4_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3680" *)
  wire cvt_4_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6452" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4886" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_4_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1999" *)
  reg cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2095" *)
  reg cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:945" *)
  wire cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5531" *)
  wire [17:0] cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6298" *)
  wire [17:0] cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:900" *)
  wire [49:0] cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6337" *)
  wire cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:898" *)
  wire cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:899" *)
  wire cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6138" *)
  wire [14:0] cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2580" *)
  wire cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6382" *)
  wire cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6383" *)
  wire [23:0] cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4391" *)
  wire [32:0] cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6169" *)
  wire cvt_5_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2025" *)
  reg cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3642" *)
  wire cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6167" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1554" *)
  reg cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1930" *)
  reg [4:0] cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1412" *)
  reg cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1820" *)
  reg cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2097" *)
  reg cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:892" *)
  wire cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3675" *)
  wire cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6416" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5302" *)
  wire [4:0] cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3420" *)
  wire cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1972" *)
  reg cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2788" *)
  wire [16:0] cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6516" *)
  wire cvt_5_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2921" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6517" *)
  wire [22:0] cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6217" *)
  wire [9:0] cvt_5_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1414" *)
  reg cvt_5_FpMantRNE_17U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:928" *)
  wire cvt_5_FpMantRNE_17U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6029" *)
  wire [9:0] cvt_5_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1375" *)
  reg cvt_5_FpMantRNE_24U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1719" *)
  reg cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:832" *)
  wire cvt_5_FpMantRNE_24U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3631" *)
  wire cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5981" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3596" *)
  wire cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5911" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:984" *)
  wire [4:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1668" *)
  reg cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2052" *)
  reg cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3597" *)
  wire cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5913" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2050" *)
  reg cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3697" *)
  wire cvt_5_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6560" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3660" *)
  wire cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6339" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_5_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3681" *)
  wire cvt_5_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6456" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3641" *)
  wire cvt_5_IntSaturation_17U_8U_if_acc_1_itm_10_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6165" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_5_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2098" *)
  reg cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1998" *)
  reg cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2096" *)
  reg cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:944" *)
  wire cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5528" *)
  wire [17:0] cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6308" *)
  wire [17:0] cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:895" *)
  wire [49:0] cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6350" *)
  wire cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:893" *)
  wire cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:894" *)
  wire cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6139" *)
  wire [14:0] cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2581" *)
  wire cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6384" *)
  wire cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6385" *)
  wire [23:0] cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4404" *)
  wire [32:0] cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6175" *)
  wire cvt_6_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2023" *)
  reg cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3041" *)
  wire cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3042" *)
  wire cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3644" *)
  wire cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6173" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1551" *)
  reg cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1933" *)
  reg [4:0] cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1418" *)
  reg cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1828" *)
  reg cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:887" *)
  wire cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6418" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3785" *)
  wire cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5318" *)
  wire [4:0] cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3421" *)
  wire cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1973" *)
  reg cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2790" *)
  wire [16:0] cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6519" *)
  wire cvt_6_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2922" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6520" *)
  wire [22:0] cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6220" *)
  wire [9:0] cvt_6_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1420" *)
  reg cvt_6_FpMantRNE_17U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:927" *)
  wire cvt_6_FpMantRNE_17U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6038" *)
  wire [9:0] cvt_6_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1376" *)
  reg cvt_6_FpMantRNE_24U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1724" *)
  reg cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:831" *)
  wire cvt_6_FpMantRNE_24U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3630" *)
  wire cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5979" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3598" *)
  wire cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5915" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:980" *)
  wire [4:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1665" *)
  reg cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2056" *)
  reg cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3599" *)
  wire cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5917" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2054" *)
  reg cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4395" *)
  wire [48:0] cvt_6_IntMulExt_33U_16U_49U_o_mul_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3698" *)
  wire cvt_6_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6562" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3661" *)
  wire cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6341" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_6_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3682" *)
  wire cvt_6_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6460" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4973" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_6_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1997" *)
  reg cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2099" *)
  reg cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:943" *)
  wire cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5525" *)
  wire [17:0] cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6302" *)
  wire [17:0] cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:890" *)
  wire [49:0] cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6343" *)
  wire cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:888" *)
  wire cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:889" *)
  wire cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6140" *)
  wire [14:0] cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2582" *)
  wire cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6386" *)
  wire cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6387" *)
  wire [23:0] cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4396" *)
  wire [32:0] cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6183" *)
  wire cvt_7_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2021" *)
  reg cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3647" *)
  wire cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6181" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1512" *)
  reg cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1936" *)
  reg [4:0] cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1426" *)
  reg cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1836" *)
  reg cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:882" *)
  wire cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6420" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3786" *)
  wire cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5329" *)
  wire [4:0] cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3422" *)
  wire cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1974" *)
  reg cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2791" *)
  wire [16:0] cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6522" *)
  wire cvt_7_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2923" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6523" *)
  wire [22:0] cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6226" *)
  wire [9:0] cvt_7_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1428" *)
  reg cvt_7_FpMantRNE_17U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:926" *)
  wire cvt_7_FpMantRNE_17U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6047" *)
  wire [9:0] cvt_7_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1377" *)
  reg cvt_7_FpMantRNE_24U_11U_else_and_2_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1730" *)
  reg cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:830" *)
  wire cvt_7_FpMantRNE_24U_11U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3629" *)
  wire cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5977" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3600" *)
  wire cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5919" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:977" *)
  wire [4:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1662" *)
  reg cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2059" *)
  reg cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3601" *)
  wire cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5921" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2057" *)
  reg cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4401" *)
  wire [48:0] cvt_7_IntMulExt_33U_16U_49U_o_mul_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3699" *)
  wire cvt_7_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6564" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3662" *)
  wire cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6344" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_7_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3683" *)
  wire cvt_7_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6464" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5022" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_7_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1996" *)
  reg cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2100" *)
  reg cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:942" *)
  wire cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5522" *)
  wire [17:0] cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6306" *)
  wire [17:0] cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:885" *)
  wire [49:0] cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6349" *)
  wire cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:883" *)
  wire cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:884" *)
  wire cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6141" *)
  wire [14:0] cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2583" *)
  wire cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6388" *)
  wire cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6389" *)
  wire [23:0] cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4402" *)
  wire [32:0] cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6189" *)
  wire cvt_8_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2019" *)
  reg cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3649" *)
  wire cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6187" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1517" *)
  reg cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1939" *)
  reg [4:0] cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1433" *)
  reg cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1844" *)
  reg cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:877" *)
  wire cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6422" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3787" *)
  wire cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5344" *)
  wire [4:0] cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3423" *)
  wire cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1975" *)
  reg cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2792" *)
  wire [16:0] cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6525" *)
  wire cvt_8_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2924" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6526" *)
  wire [22:0] cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6232" *)
  wire [9:0] cvt_8_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1435" *)
  reg cvt_8_FpMantRNE_17U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:925" *)
  wire cvt_8_FpMantRNE_17U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6056" *)
  wire [9:0] cvt_8_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1378" *)
  reg cvt_8_FpMantRNE_24U_11U_else_and_3_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1736" *)
  reg cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:829" *)
  wire cvt_8_FpMantRNE_24U_11U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3628" *)
  wire cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5975" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3602" *)
  wire cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5923" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:974" *)
  wire [4:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1659" *)
  reg cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2062" *)
  reg cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3603" *)
  wire cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5925" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2060" *)
  reg cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4398" *)
  wire [48:0] cvt_8_IntMulExt_33U_16U_49U_o_mul_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3700" *)
  wire cvt_8_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6566" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3663" *)
  wire cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6346" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_8_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3684" *)
  wire cvt_8_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6468" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5102" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_8_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1995" *)
  reg cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2101" *)
  reg cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:941" *)
  wire cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5519" *)
  wire [17:0] cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6304" *)
  wire [17:0] cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:880" *)
  wire [49:0] cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6348" *)
  wire cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:878" *)
  wire cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:879" *)
  wire cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6142" *)
  wire [14:0] cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2584" *)
  wire cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6390" *)
  wire cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6391" *)
  wire [23:0] cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4399" *)
  wire [32:0] cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6197" *)
  wire cvt_9_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2017" *)
  reg cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3053" *)
  wire cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3054" *)
  wire cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3652" *)
  wire cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6195" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10" *)
  wire [11:0] cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1546" *)
  reg cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1942" *)
  reg [4:0] cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1851" *)
  reg cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2104" *)
  reg cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:872" *)
  wire cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3676" *)
  wire cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6424" *)
  (* unused_bits = "0 1 2 3" *)
  wire [4:0] cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5358" *)
  wire [4:0] cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3424" *)
  wire cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1976" *)
  reg cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6528" *)
  wire cvt_9_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2925" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12" *)
  wire [23:0] cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6529" *)
  wire [22:0] cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5162" *)
  wire [9:0] cvt_9_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1440" *)
  reg cvt_9_FpMantRNE_17U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:924" *)
  wire cvt_9_FpMantRNE_17U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6065" *)
  wire [9:0] cvt_9_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1379" *)
  reg cvt_9_FpMantRNE_24U_11U_else_and_1_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1742" *)
  reg cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:828" *)
  wire cvt_9_FpMantRNE_24U_11U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3627" *)
  wire cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5973" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3604" *)
  wire cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5927" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:971" *)
  wire [4:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1656" *)
  reg cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2065" *)
  reg cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3605" *)
  wire cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5929" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2063" *)
  reg cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3701" *)
  wire cvt_9_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6568" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3664" *)
  wire cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6351" *)
  (* unused_bits = "0 1" *)
  wire [2:0] cvt_9_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3685" *)
  wire cvt_9_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6472" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3651" *)
  wire cvt_9_IntSaturation_17U_8U_if_acc_1_itm_10_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6193" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] cvt_9_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2106" *)
  reg cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1994" *)
  reg cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1850" *)
  reg cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:940" *)
  wire cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5516" *)
  wire [17:0] cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6324" *)
  wire [17:0] cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:875" *)
  wire [49:0] cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6374" *)
  wire cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:873" *)
  wire cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:874" *)
  wire cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6143" *)
  wire [14:0] cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2585" *)
  wire cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6392" *)
  wire cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6393" *)
  wire [23:0] cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4431" *)
  wire [32:0] cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2219" *)
  wire cvt_and_147_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4006" *)
  wire cvt_and_231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4007" *)
  wire cvt_and_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3998" *)
  wire cvt_and_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3999" *)
  wire cvt_and_234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3994" *)
  wire cvt_and_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3995" *)
  wire cvt_and_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3985" *)
  wire cvt_and_237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3986" *)
  wire cvt_and_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3979" *)
  wire cvt_and_239_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3980" *)
  wire cvt_and_240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3972" *)
  wire cvt_and_241_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3973" *)
  wire cvt_and_242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3966" *)
  wire cvt_and_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3967" *)
  wire cvt_and_244_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3963" *)
  wire cvt_and_245_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3964" *)
  wire cvt_and_246_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3957" *)
  wire cvt_and_247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3958" *)
  wire cvt_and_248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3950" *)
  wire cvt_and_249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3951" *)
  wire cvt_and_250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3944" *)
  wire cvt_and_251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3945" *)
  wire cvt_and_252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3941" *)
  wire cvt_and_253_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3942" *)
  wire cvt_and_254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3936" *)
  wire cvt_and_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3937" *)
  wire cvt_and_256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3932" *)
  wire cvt_and_257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3933" *)
  wire cvt_and_258_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3926" *)
  wire cvt_and_259_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3927" *)
  wire cvt_and_260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3923" *)
  wire cvt_and_261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3924" *)
  wire cvt_and_262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2934" *)
  wire cvt_and_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3389" *)
  wire cvt_asn_319;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3390" *)
  wire cvt_asn_321;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3391" *)
  wire cvt_asn_323;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3392" *)
  wire cvt_asn_327;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3393" *)
  wire cvt_asn_329;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3394" *)
  wire cvt_asn_333;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3395" *)
  wire cvt_asn_335;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3396" *)
  wire cvt_asn_339;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3397" *)
  wire cvt_asn_341;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3398" *)
  wire cvt_asn_345;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3399" *)
  wire cvt_asn_347;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3400" *)
  wire cvt_asn_351;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3401" *)
  wire cvt_asn_353;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3402" *)
  wire cvt_asn_357;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3403" *)
  wire cvt_asn_359;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3404" *)
  wire cvt_asn_363;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3405" *)
  wire cvt_asn_365;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3406" *)
  wire cvt_asn_369;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3407" *)
  wire cvt_asn_371;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3408" *)
  wire cvt_asn_375;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3409" *)
  wire cvt_asn_377;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3410" *)
  wire cvt_asn_381;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3411" *)
  wire cvt_asn_383;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3412" *)
  wire cvt_asn_387;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3413" *)
  wire cvt_asn_389;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3414" *)
  wire cvt_asn_393;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3415" *)
  wire cvt_asn_399;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2576" *)
  wire cvt_cvt_nand_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2522" *)
  wire cvt_else_and_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2523" *)
  wire cvt_else_and_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3463" *)
  wire cvt_else_and_24_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3464" *)
  wire cvt_else_and_34_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2521" *)
  wire cvt_else_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2226" *)
  wire cvt_else_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2225" *)
  wire cvt_else_equal_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2198" *)
  wire cvt_else_equal_tmp_10_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2208" *)
  wire cvt_else_equal_tmp_15_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1422" *)
  reg cvt_else_equal_tmp_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2207" *)
  wire cvt_else_equal_tmp_16_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2214" *)
  wire cvt_else_equal_tmp_18_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2213" *)
  wire cvt_else_equal_tmp_19_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2220" *)
  wire cvt_else_equal_tmp_21_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2218" *)
  wire cvt_else_equal_tmp_22_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2232" *)
  wire cvt_else_equal_tmp_27_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1448" *)
  reg cvt_else_equal_tmp_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2231" *)
  wire cvt_else_equal_tmp_28_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2229" *)
  wire cvt_else_equal_tmp_30_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2228" *)
  wire cvt_else_equal_tmp_31_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1464" *)
  reg cvt_else_equal_tmp_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2223" *)
  wire cvt_else_equal_tmp_33_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1465" *)
  reg cvt_else_equal_tmp_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2222" *)
  wire cvt_else_equal_tmp_34_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2217" *)
  wire cvt_else_equal_tmp_36_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2216" *)
  wire cvt_else_equal_tmp_37_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2211" *)
  wire cvt_else_equal_tmp_39_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2196" *)
  wire cvt_else_equal_tmp_3_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2210" *)
  wire cvt_else_equal_tmp_40_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2205" *)
  wire cvt_else_equal_tmp_42_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2204" *)
  wire cvt_else_equal_tmp_43_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1496" *)
  reg cvt_else_equal_tmp_45;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2202" *)
  wire cvt_else_equal_tmp_45_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1497" *)
  reg cvt_else_equal_tmp_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2201" *)
  wire cvt_else_equal_tmp_46_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2195" *)
  wire cvt_else_equal_tmp_4_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1396" *)
  reg cvt_else_equal_tmp_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1409" *)
  reg cvt_else_equal_tmp_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2199" *)
  wire cvt_else_equal_tmp_9_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4075" *)
  wire cvt_else_mux1h_103_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4072" *)
  wire cvt_else_mux1h_105_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4016" *)
  wire cvt_else_mux1h_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4086" *)
  wire cvt_else_mux1h_122_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4083" *)
  wire cvt_else_mux1h_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4097" *)
  wire cvt_else_mux1h_141_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4094" *)
  wire cvt_else_mux1h_143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4108" *)
  wire cvt_else_mux1h_160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4105" *)
  wire cvt_else_mux1h_162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4119" *)
  wire cvt_else_mux1h_179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4116" *)
  wire cvt_else_mux1h_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4130" *)
  wire cvt_else_mux1h_198_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4127" *)
  wire cvt_else_mux1h_200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4141" *)
  wire cvt_else_mux1h_217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4138" *)
  wire cvt_else_mux1h_219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4152" *)
  wire cvt_else_mux1h_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4149" *)
  wire cvt_else_mux1h_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4162" *)
  wire cvt_else_mux1h_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4173" *)
  wire cvt_else_mux1h_274_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4170" *)
  wire cvt_else_mux1h_276_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4031" *)
  wire cvt_else_mux1h_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4183" *)
  wire cvt_else_mux1h_292_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4176" *)
  wire cvt_else_mux1h_295_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4028" *)
  wire cvt_else_mux1h_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4042" *)
  wire cvt_else_mux1h_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4039" *)
  wire cvt_else_mux1h_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4053" *)
  wire cvt_else_mux1h_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4050" *)
  wire cvt_else_mux1h_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4064" *)
  wire cvt_else_mux1h_84_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4061" *)
  wire cvt_else_mux1h_86_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4020" *)
  wire cvt_else_mux1h_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6208" *)
  wire cvt_else_mux_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6210" *)
  wire cvt_else_mux_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6209" *)
  wire cvt_else_mux_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2227" *)
  wire cvt_else_nor_dfs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1456" *)
  reg cvt_else_nor_dfs_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2230" *)
  wire cvt_else_nor_dfs_10_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1466" *)
  reg cvt_else_nor_dfs_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2224" *)
  wire cvt_else_nor_dfs_11_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2212" *)
  wire cvt_else_nor_dfs_13_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2206" *)
  wire cvt_else_nor_dfs_14_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1498" *)
  reg cvt_else_nor_dfs_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2203" *)
  wire cvt_else_nor_dfs_15_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2197" *)
  wire cvt_else_nor_dfs_1_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1397" *)
  reg cvt_else_nor_dfs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2200" *)
  wire cvt_else_nor_dfs_3_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2209" *)
  wire cvt_else_nor_dfs_5_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2215" *)
  wire cvt_else_nor_dfs_6_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2221" *)
  wire cvt_else_nor_dfs_7_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2233" *)
  wire cvt_else_nor_dfs_9_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4078" *)
  wire cvt_if_mux_100_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4011" *)
  wire cvt_if_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4098" *)
  wire cvt_if_mux_113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4089" *)
  wire cvt_if_mux_115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4109" *)
  wire cvt_if_mux_128_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4100" *)
  wire cvt_if_mux_130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4120" *)
  wire cvt_if_mux_143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4111" *)
  wire cvt_if_mux_145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4131" *)
  wire cvt_if_mux_158_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4122" *)
  wire cvt_if_mux_160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4142" *)
  wire cvt_if_mux_173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4133" *)
  wire cvt_if_mux_175_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4153" *)
  wire cvt_if_mux_188_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4144" *)
  wire cvt_if_mux_190_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4163" *)
  wire cvt_if_mux_203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4155" *)
  wire cvt_if_mux_205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4174" *)
  wire cvt_if_mux_218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4165" *)
  wire cvt_if_mux_220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4184" *)
  wire cvt_if_mux_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4178" *)
  wire cvt_if_mux_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4032" *)
  wire cvt_if_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4023" *)
  wire cvt_if_mux_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4043" *)
  wire cvt_if_mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4034" *)
  wire cvt_if_mux_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4054" *)
  wire cvt_if_mux_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4045" *)
  wire cvt_if_mux_55_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4065" *)
  wire cvt_if_mux_68_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4056" *)
  wire cvt_if_mux_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4076" *)
  wire cvt_if_mux_83_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4067" *)
  wire cvt_if_mux_85_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4021" *)
  wire cvt_if_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4087" *)
  wire cvt_if_mux_98_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2234" *)
  wire cvt_if_unequal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4015" *)
  wire cvt_mux_2280_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4010" *)
  wire cvt_mux_2281_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4027" *)
  wire cvt_mux_2284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4022" *)
  wire cvt_mux_2285_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4038" *)
  wire cvt_mux_2288_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4033" *)
  wire cvt_mux_2289_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4049" *)
  wire cvt_mux_2292_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4044" *)
  wire cvt_mux_2293_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4060" *)
  wire cvt_mux_2296_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4055" *)
  wire cvt_mux_2297_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4071" *)
  wire cvt_mux_2300_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4066" *)
  wire cvt_mux_2301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4082" *)
  wire cvt_mux_2304_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4077" *)
  wire cvt_mux_2305_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4093" *)
  wire cvt_mux_2308_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4088" *)
  wire cvt_mux_2309_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4104" *)
  wire cvt_mux_2312_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4099" *)
  wire cvt_mux_2313_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4115" *)
  wire cvt_mux_2316_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4110" *)
  wire cvt_mux_2317_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4126" *)
  wire cvt_mux_2320_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4121" *)
  wire cvt_mux_2321_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4137" *)
  wire cvt_mux_2324_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4132" *)
  wire cvt_mux_2325_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4148" *)
  wire cvt_mux_2328_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4143" *)
  wire cvt_mux_2329_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4159" *)
  wire cvt_mux_2332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4154" *)
  wire cvt_mux_2333_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4169" *)
  wire cvt_mux_2336_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4164" *)
  wire cvt_mux_2337_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4175" *)
  wire cvt_mux_2340_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4182" *)
  wire cvt_mux_2341_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4030" *)
  wire cvt_mux_2346_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4041" *)
  wire cvt_mux_2348_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4052" *)
  wire cvt_mux_2350_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4063" *)
  wire cvt_mux_2352_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4074" *)
  wire cvt_mux_2354_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4172" *)
  wire cvt_mux_2356_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4085" *)
  wire cvt_mux_2358_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4096" *)
  wire cvt_mux_2360_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4107" *)
  wire cvt_mux_2362_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4118" *)
  wire cvt_mux_2364_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4129" *)
  wire cvt_mux_2366_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4161" *)
  wire cvt_mux_2368_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4140" *)
  wire cvt_mux_2370_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4151" *)
  wire cvt_mux_2372_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4019" *)
  wire cvt_mux_2373_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2482" *)
  wire cvt_or_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2483" *)
  wire cvt_or_12_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2484" *)
  wire cvt_or_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2485" *)
  wire cvt_or_18_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2486" *)
  wire cvt_or_20_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2487" *)
  wire cvt_or_22_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2488" *)
  wire cvt_or_24_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2489" *)
  wire cvt_or_26_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2490" *)
  wire cvt_or_28_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2480" *)
  wire cvt_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2491" *)
  wire cvt_or_30_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4018" *)
  wire cvt_or_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2481" *)
  wire cvt_or_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2478" *)
  wire cvt_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1688" *)
  reg cvt_unequal_tmp_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1689" *)
  reg cvt_unequal_tmp_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1690" *)
  reg cvt_unequal_tmp_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:820" *)
  wire [1:0] fsm_output;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3432" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3433" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3434" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3435" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3436" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3437" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3438" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3439" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3440" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3441" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3442" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3443" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3444" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3445" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3446" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3447" *)
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2194" *)
  wire main_stage_en_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1499" *)
  reg main_stage_v_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2940" *)
  wire main_stage_v_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1500" *)
  reg main_stage_v_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2985" *)
  wire main_stage_v_2_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1501" *)
  reg main_stage_v_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3023" *)
  wire main_stage_v_3_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5222" *)
  wire mux_1000_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5226" *)
  wire mux_1001_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5228" *)
  wire mux_1002_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5225" *)
  wire mux_1003_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5234" *)
  wire mux_1004_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5247" *)
  wire mux_1010_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5245" *)
  wire mux_1011_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5255" *)
  wire mux_1012_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6737" *)
  wire mux_1013_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6736" *)
  wire mux_1014_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5254" *)
  wire mux_1016_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5257" *)
  wire mux_1017_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5253" *)
  wire mux_1018_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5270" *)
  wire mux_1027_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5284" *)
  wire mux_1034_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5283" *)
  wire mux_1035_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6743" *)
  wire mux_1040_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6744" *)
  wire mux_1042_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5290" *)
  wire mux_1044_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5289" *)
  wire mux_1045_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6745" *)
  wire mux_1046_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6746" *)
  wire mux_1048_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5286" *)
  wire mux_1050_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5285" *)
  wire mux_1051_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5287" *)
  wire mux_1052_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3782" *)
  wire mux_1053_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5288" *)
  wire mux_1054_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5312" *)
  wire mux_1069_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5310" *)
  wire mux_1070_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3521" *)
  wire mux_1071_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6748" *)
  wire mux_1072_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6747" *)
  wire mux_1073_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5316" *)
  wire mux_1075_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5317" *)
  wire mux_1076_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5315" *)
  wire mux_1077_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6752" *)
  wire mux_1086_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6751" *)
  wire mux_1087_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5327" *)
  wire mux_1089_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5328" *)
  wire mux_1090_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5326" *)
  wire mux_1091_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6586" *)
  wire mux_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4207" *)
  wire mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6759" *)
  wire mux_1102_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6760" *)
  wire mux_1104_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5339" *)
  wire mux_1106_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5338" *)
  wire mux_1107_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6761" *)
  wire mux_1108_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3526" *)
  wire mux_110_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6762" *)
  wire mux_1110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5342" *)
  wire mux_1112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5341" *)
  wire mux_1113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5343" *)
  wire mux_1114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5340" *)
  wire mux_1115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5337" *)
  wire mux_1116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2693" *)
  wire mux_1126_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5356" *)
  wire mux_1127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5367" *)
  wire mux_1133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5366" *)
  wire mux_1134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2733" *)
  wire mux_1142_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6763" *)
  wire mux_1151_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5379" *)
  wire mux_1153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5378" *)
  wire mux_1154_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5377" *)
  wire mux_1163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5391" *)
  wire mux_1172_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5390" *)
  wire mux_1173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5389" *)
  wire mux_1174_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5396" *)
  wire mux_1175_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5395" *)
  wire mux_1176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5394" *)
  wire mux_1177_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5393" *)
  wire mux_1178_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5388" *)
  wire mux_1179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5587" *)
  wire mux_118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5878" *)
  wire mux_119_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4210" *)
  wire mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5420" *)
  wire mux_1202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5419" *)
  wire mux_1203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5417" *)
  wire mux_1204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5425" *)
  wire mux_1211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5424" *)
  wire mux_1212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5422" *)
  wire mux_1213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5880" *)
  wire mux_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5585" *)
  wire mux_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5454" *)
  wire mux_1252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5881" *)
  wire mux_125_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5452" *)
  wire mux_1262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5457" *)
  wire mux_1265_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5456" *)
  wire mux_1266_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5459" *)
  wire mux_1267_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5461" *)
  wire mux_1268_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6769" *)
  wire mux_1269_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6774" *)
  wire mux_1271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6773" *)
  wire mux_1272_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6772" *)
  wire mux_1273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6771" *)
  wire mux_1274_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6770" *)
  wire mux_1275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6775" *)
  wire mux_1281_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5873" *)
  wire mux_1283_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5872" *)
  wire mux_1284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5871" *)
  wire mux_1285_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5870" *)
  wire mux_1286_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4213" *)
  wire mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5586" *)
  wire mux_130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5883" *)
  wire mux_131_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6776" *)
  wire mux_1325_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6781" *)
  wire mux_1327_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6780" *)
  wire mux_1328_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6779" *)
  wire mux_1329_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6778" *)
  wire mux_1330_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6777" *)
  wire mux_1331_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6782" *)
  wire mux_1338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3730" *)
  wire mux_133_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6783" *)
  wire mux_1340_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5546" *)
  wire mux_1342_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5545" *)
  wire mux_1343_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5544" *)
  wire mux_1344_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5543" *)
  wire mux_1345_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3777" *)
  wire mux_134_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4215" *)
  wire mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6787" *)
  wire mux_1405_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6786" *)
  wire mux_1406_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6785" *)
  wire mux_1407_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6784" *)
  wire mux_1408_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5877" *)
  wire mux_1412_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5876" *)
  wire mux_1413_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5875" *)
  wire mux_1414_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5874" *)
  wire mux_1415_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6791" *)
  wire mux_1416_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6790" *)
  wire mux_1417_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6789" *)
  wire mux_1418_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5555" *)
  wire mux_1420_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5554" *)
  wire mux_1421_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5553" *)
  wire mux_1423_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5552" *)
  wire mux_1424_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5551" *)
  wire mux_1425_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5550" *)
  wire mux_1426_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5549" *)
  wire mux_1427_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5548" *)
  wire mux_1428_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5547" *)
  wire mux_1429_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6798" *)
  wire mux_1430_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6797" *)
  wire mux_1431_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6796" *)
  wire mux_1432_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6795" *)
  wire mux_1433_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6794" *)
  wire mux_1434_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2692" *)
  wire mux_1436_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3761" *)
  wire mux_1437_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5562" *)
  wire mux_1438_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5561" *)
  wire mux_1439_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5886" *)
  wire mux_143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5560" *)
  wire mux_1441_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5559" *)
  wire mux_1442_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5563" *)
  wire mux_1458_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3527" *)
  wire mux_1460_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5568" *)
  wire mux_1461_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3748" *)
  wire mux_1463_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2694" *)
  wire mux_1464_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5567" *)
  wire mux_1465_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3732" *)
  wire mux_1466_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5572" *)
  wire mux_1467_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5576" *)
  wire mux_1470_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5574" *)
  wire mux_1471_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5571" *)
  wire mux_1472_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3763" *)
  wire mux_1489_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6591" *)
  wire mux_148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5581" *)
  wire mux_1490_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2730" *)
  wire mux_1494_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5580" *)
  wire mux_1495_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5588" *)
  wire mux_149_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4214" *)
  wire mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5888" *)
  wire mux_150_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5583" *)
  wire mux_1519_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3764" *)
  wire mux_1521_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5589" *)
  wire mux_152_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5592" *)
  wire mux_1531_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5591" *)
  wire mux_1532_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5590" *)
  wire mux_1533_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5594" *)
  wire mux_1534_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5597" *)
  wire mux_1535_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5600" *)
  wire mux_1536_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5603" *)
  wire mux_1537_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5606" *)
  wire mux_1538_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5609" *)
  wire mux_1539_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5890" *)
  wire mux_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5612" *)
  wire mux_1540_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5615" *)
  wire mux_1541_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5618" *)
  wire mux_1542_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5621" *)
  wire mux_1543_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5624" *)
  wire mux_1544_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5627" *)
  wire mux_1545_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5630" *)
  wire mux_1546_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5633" *)
  wire mux_1547_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5636" *)
  wire mux_1548_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5639" *)
  wire mux_1549_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4424" *)
  wire mux_154_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5642" *)
  wire mux_1550_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5645" *)
  wire mux_1551_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5648" *)
  wire mux_1552_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5651" *)
  wire mux_1553_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5654" *)
  wire mux_1554_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5657" *)
  wire mux_1555_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5660" *)
  wire mux_1556_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5663" *)
  wire mux_1557_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5666" *)
  wire mux_1558_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5669" *)
  wire mux_1559_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4423" *)
  wire mux_155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5672" *)
  wire mux_1560_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5675" *)
  wire mux_1561_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5678" *)
  wire mux_1562_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5681" *)
  wire mux_1563_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5684" *)
  wire mux_1564_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5687" *)
  wire mux_1565_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5691" *)
  wire mux_1567_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5692" *)
  wire mux_1568_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5690" *)
  wire mux_1569_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5696" *)
  wire mux_1571_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5697" *)
  wire mux_1572_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5695" *)
  wire mux_1573_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5701" *)
  wire mux_1575_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5702" *)
  wire mux_1576_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5700" *)
  wire mux_1577_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5706" *)
  wire mux_1579_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5707" *)
  wire mux_1580_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5705" *)
  wire mux_1581_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5711" *)
  wire mux_1583_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5712" *)
  wire mux_1584_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5710" *)
  wire mux_1585_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5716" *)
  wire mux_1587_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5717" *)
  wire mux_1588_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5715" *)
  wire mux_1589_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5721" *)
  wire mux_1590_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5720" *)
  wire mux_1591_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5728" *)
  wire mux_1593_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5729" *)
  wire mux_1594_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5727" *)
  wire mux_1595_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5733" *)
  wire mux_1597_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5734" *)
  wire mux_1598_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5732" *)
  wire mux_1599_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4421" *)
  wire mux_159_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4220" *)
  wire mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5738" *)
  wire mux_1601_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5739" *)
  wire mux_1602_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5737" *)
  wire mux_1603_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5743" *)
  wire mux_1604_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5742" *)
  wire mux_1605_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5750" *)
  wire mux_1607_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5751" *)
  wire mux_1608_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5749" *)
  wire mux_1609_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5755" *)
  wire mux_1611_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5756" *)
  wire mux_1612_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5754" *)
  wire mux_1613_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5760" *)
  wire mux_1615_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5761" *)
  wire mux_1616_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5759" *)
  wire mux_1617_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5765" *)
  wire mux_1619_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5766" *)
  wire mux_1620_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5764" *)
  wire mux_1621_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5770" *)
  wire mux_1623_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5771" *)
  wire mux_1624_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5769" *)
  wire mux_1625_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5774" *)
  wire mux_1626_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5776" *)
  wire mux_1627_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4435" *)
  wire mux_162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5781" *)
  wire mux_1632_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5780" *)
  wire mux_1633_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5783" *)
  wire mux_1638_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5782" *)
  wire mux_1639_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4437" *)
  wire mux_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5779" *)
  wire mux_1640_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5787" *)
  wire mux_1643_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5786" *)
  wire mux_1644_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5789" *)
  wire mux_1647_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5788" *)
  wire mux_1648_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5785" *)
  wire mux_1649_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5790" *)
  wire mux_1653_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3750" *)
  wire mux_1654_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5794" *)
  wire mux_1658_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5793" *)
  wire mux_1659_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5792" *)
  wire mux_1660_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5797" *)
  wire mux_1661_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5798" *)
  wire mux_1662_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5796" *)
  wire mux_1663_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3713" *)
  wire mux_166_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5802" *)
  wire mux_1672_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5801" *)
  wire mux_1673_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5800" *)
  wire mux_1674_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4439" *)
  wire mux_167_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5806" *)
  wire mux_1683_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5805" *)
  wire mux_1684_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5804" *)
  wire mux_1685_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5828" *)
  wire mux_1687_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5831" *)
  wire mux_1689_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5834" *)
  wire mux_1692_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5837" *)
  wire mux_1694_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5840" *)
  wire mux_1697_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4440" *)
  wire mux_169_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4219" *)
  wire mux_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5843" *)
  wire mux_1700_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5846" *)
  wire mux_1704_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5849" *)
  wire mux_1707_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5852" *)
  wire mux_1711_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5855" *)
  wire mux_1715_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5858" *)
  wire mux_1720_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5861" *)
  wire mux_1727_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5864" *)
  wire mux_1734_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5867" *)
  wire mux_1743_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4512" *)
  wire mux_1750_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4511" *)
  wire mux_1751_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4510" *)
  wire mux_1752_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4532" *)
  wire mux_1757_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4530" *)
  wire mux_1758_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4441" *)
  wire mux_175_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4558" *)
  wire mux_1760_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3740" *)
  wire mux_1761_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3517" *)
  wire mux_1762_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4602" *)
  wire mux_1772_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3741" *)
  wire mux_1779_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4639" *)
  wire mux_1780_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4658" *)
  wire mux_1785_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4679" *)
  wire mux_1788_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4706" *)
  wire mux_1790_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4705" *)
  wire mux_1791_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4724" *)
  wire mux_1794_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4729" *)
  wire mux_1796_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4727" *)
  wire mux_1797_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4726" *)
  wire mux_1798_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4723" *)
  wire mux_1799_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4222" *)
  wire mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4760" *)
  wire mux_1807_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4759" *)
  wire mux_1808_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4792" *)
  wire mux_1814_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4790" *)
  wire mux_1815_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4789" *)
  wire mux_1816_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4788" *)
  wire mux_1817_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4864" *)
  wire mux_1828_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4866" *)
  wire mux_1830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4863" *)
  wire mux_1831_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5014" *)
  wire mux_1832_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6807" *)
  wire mux_1836_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6803" *)
  wire mux_1839_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6804" *)
  wire mux_1841_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6809" *)
  wire mux_1846_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3759" *)
  wire mux_1849_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3718" *)
  wire mux_1851_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3771" *)
  wire mux_1852_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4916" *)
  wire mux_1859_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3746" *)
  wire mux_1864_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4961" *)
  wire mux_1867_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6811" *)
  wire mux_1876_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3745" *)
  wire mux_1881_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3507" *)
  wire mux_1882_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4990" *)
  wire mux_1886_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5012" *)
  wire mux_1888_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5010" *)
  wire mux_1889_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6595" *)
  wire mux_188_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5024" *)
  wire mux_1892_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4226" *)
  wire mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6813" *)
  wire mux_1903_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5089" *)
  wire mux_1909_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4443" *)
  wire mux_190_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5104" *)
  wire mux_1916_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4442" *)
  wire mux_191_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6815" *)
  wire mux_1927_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4444" *)
  wire mux_192_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5144" *)
  wire mux_1930_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5143" *)
  wire mux_1933_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6817" *)
  wire mux_1940_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6819" *)
  wire mux_1943_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6821" *)
  wire mux_1953_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6823" *)
  wire mux_1964_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2933" *)
  wire mux_1966_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4225" *)
  wire mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4192" *)
  wire mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5435" *)
  wire mux_2000_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5481" *)
  wire mux_2010_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5480" *)
  wire mux_2011_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5483" *)
  wire mux_2012_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5484" *)
  wire mux_2013_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5482" *)
  wire mux_2014_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5478" *)
  wire mux_2015_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5488" *)
  wire mux_2017_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5491" *)
  wire mux_2018_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5489" *)
  wire mux_2019_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2732" *)
  wire mux_201_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5486" *)
  wire mux_2020_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5827" *)
  wire mux_207_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5826" *)
  wire mux_208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4231" *)
  wire mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4533" *)
  wire mux_2170_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4636" *)
  wire mux_2171_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4515" *)
  wire mux_2172_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4514" *)
  wire mux_2173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4513" *)
  wire mux_2174_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4535" *)
  wire mux_2175_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4534" *)
  wire mux_2176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4563" *)
  wire mux_2177_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4562" *)
  wire mux_2178_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4561" *)
  wire mux_2179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4605" *)
  wire mux_2183_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4604" *)
  wire mux_2185_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4603" *)
  wire mux_2186_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4682" *)
  wire mux_2193_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4681" *)
  wire mux_2195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4680" *)
  wire mux_2196_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4230" *)
  wire mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6829" *)
  wire mux_2200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6828" *)
  wire mux_2201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6830" *)
  wire mux_2202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6827" *)
  wire mux_2203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6826" *)
  wire mux_2204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6825" *)
  wire mux_2205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6833" *)
  wire mux_2207_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6832" *)
  wire mux_2208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4736" *)
  wire mux_2210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4735" *)
  wire mux_2211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4734" *)
  wire mux_2212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4733" *)
  wire mux_2213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4732" *)
  wire mux_2214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4765" *)
  wire mux_2215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4764" *)
  wire mux_2216_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4763" *)
  wire mux_2217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4762" *)
  wire mux_2218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4796" *)
  wire mux_2219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4795" *)
  wire mux_2221_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4794" *)
  wire mux_2222_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4793" *)
  wire mux_2223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4868" *)
  wire mux_2224_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4883" *)
  wire mux_2225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4882" *)
  wire mux_2226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4907" *)
  wire mux_2227_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2723" *)
  wire mux_2230_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4963" *)
  wire mux_2231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4964" *)
  wire mux_2232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4988" *)
  wire mux_2233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5090" *)
  wire mux_2236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5092" *)
  wire mux_2237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5093" *)
  wire mux_2239_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5494" *)
  wire mux_2248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5493" *)
  wire mux_2249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5241" *)
  wire mux_2250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5243" *)
  wire mux_2251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5262" *)
  wire mux_2252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5264" *)
  wire mux_2253_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5279" *)
  wire mux_2254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5281" *)
  wire mux_2255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5295" *)
  wire mux_2256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5297" *)
  wire mux_2257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5306" *)
  wire mux_2258_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5308" *)
  wire mux_2259_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5322" *)
  wire mux_2260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5324" *)
  wire mux_2261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5333" *)
  wire mux_2262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5335" *)
  wire mux_2263_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5348" *)
  wire mux_2264_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5350" *)
  wire mux_2265_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5362" *)
  wire mux_2266_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5364" *)
  wire mux_2267_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5372" *)
  wire mux_2268_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5374" *)
  wire mux_2269_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5384" *)
  wire mux_2270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5386" *)
  wire mux_2271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5403" *)
  wire mux_2272_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5405" *)
  wire mux_2273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5411" *)
  wire mux_2274_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5413" *)
  wire mux_2275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5431" *)
  wire mux_2276_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5433" *)
  wire mux_2277_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5440" *)
  wire mux_2278_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5442" *)
  wire mux_2279_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5448" *)
  wire mux_2280_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5450" *)
  wire mux_2281_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6835" *)
  wire mux_2299_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4233" *)
  wire mux_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3930" *)
  wire mux_2301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3929" *)
  wire mux_2302_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6836" *)
  wire mux_2303_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6837" *)
  wire mux_2305_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3939" *)
  wire mux_2307_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3938" *)
  wire mux_2308_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6838" *)
  wire mux_2309_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6839" *)
  wire mux_2311_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3948" *)
  wire mux_2313_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3947" *)
  wire mux_2314_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6840" *)
  wire mux_2315_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6841" *)
  wire mux_2317_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3954" *)
  wire mux_2319_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3953" *)
  wire mux_2320_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6842" *)
  wire mux_2322_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6843" *)
  wire mux_2324_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3961" *)
  wire mux_2326_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3960" *)
  wire mux_2327_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6844" *)
  wire mux_2329_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4447" *)
  wire mux_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3970" *)
  wire mux_2331_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3969" *)
  wire mux_2332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6845" *)
  wire mux_2333_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6846" *)
  wire mux_2335_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3976" *)
  wire mux_2337_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3975" *)
  wire mux_2338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6847" *)
  wire mux_2341_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3983" *)
  wire mux_2343_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3982" *)
  wire mux_2344_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6848" *)
  wire mux_2346_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3989" *)
  wire mux_2348_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3988" *)
  wire mux_2349_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6849" *)
  wire mux_2350_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6850" *)
  wire mux_2352_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3992" *)
  wire mux_2354_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3991" *)
  wire mux_2355_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6851" *)
  wire mux_2356_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6852" *)
  wire mux_2358_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4446" *)
  wire mux_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4003" *)
  wire mux_2360_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4002" *)
  wire mux_2361_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4001" *)
  wire mux_2362_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4452" *)
  wire mux_237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4451" *)
  wire mux_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4237" *)
  wire mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4455" *)
  wire mux_241_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4454" *)
  wire mux_242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4450" *)
  wire mux_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6603" *)
  wire mux_244_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4458" *)
  wire mux_246_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4457" *)
  wire mux_247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4461" *)
  wire mux_248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4236" *)
  wire mux_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6609" *)
  wire mux_250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6612" *)
  wire mux_252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4466" *)
  wire mux_254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4465" *)
  wire mux_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4464" *)
  wire mux_256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4463" *)
  wire mux_257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4242" *)
  wire mux_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4470" *)
  wire mux_260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4469" *)
  wire mux_261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4473" *)
  wire mux_264_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4472" *)
  wire mux_265_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4471" *)
  wire mux_266_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4468" *)
  wire mux_267_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4241" *)
  wire mux_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4476" *)
  wire mux_270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4475" *)
  wire mux_271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3726" *)
  wire mux_272_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4477" *)
  wire mux_273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4478" *)
  wire mux_275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4483" *)
  wire mux_279_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4245" *)
  wire mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4482" *)
  wire mux_280_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4485" *)
  wire mux_283_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4484" *)
  wire mux_284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4481" *)
  wire mux_285_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4488" *)
  wire mux_288_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4487" *)
  wire mux_289_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4244" *)
  wire mux_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4494" *)
  wire mux_290_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4491" *)
  wire mux_291_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4498" *)
  wire mux_295_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4497" *)
  wire mux_296_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4250" *)
  wire mux_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4190" *)
  wire mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4501" *)
  wire mux_300_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4500" *)
  wire mux_301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4496" *)
  wire mux_302_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4505" *)
  wire mux_306_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4504" *)
  wire mux_307_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6624" *)
  wire mux_308_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4249" *)
  wire mux_30_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6625" *)
  wire mux_310_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6626" *)
  wire mux_312_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4507" *)
  wire mux_314_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4506" *)
  wire mux_315_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4503" *)
  wire mux_316_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4255" *)
  wire mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3528" *)
  wire mux_320_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4516" *)
  wire mux_322_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4519" *)
  wire mux_327_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4520" *)
  wire mux_328_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4518" *)
  wire mux_329_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4254" *)
  wire mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4524" *)
  wire mux_332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4523" *)
  wire mux_333_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4526" *)
  wire mux_336_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4525" *)
  wire mux_337_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4522" *)
  wire mux_338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4259" *)
  wire mux_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4540" *)
  wire mux_341_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4538" *)
  wire mux_342_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2726" *)
  wire mux_344_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4544" *)
  wire mux_347_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4542" *)
  wire mux_348_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4258" *)
  wire mux_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4548" *)
  wire mux_352_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4547" *)
  wire mux_353_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4551" *)
  wire mux_357_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4550" *)
  wire mux_358_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4546" *)
  wire mux_359_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4264" *)
  wire mux_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4555" *)
  wire mux_363_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4554" *)
  wire mux_364_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6636" *)
  wire mux_369_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4263" *)
  wire mux_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4557" *)
  wire mux_371_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4556" *)
  wire mux_372_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4553" *)
  wire mux_373_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5809" *)
  wire mux_377_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4564" *)
  wire mux_378_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4269" *)
  wire mux_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3512" *)
  wire mux_382_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4566" *)
  wire mux_383_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4571" *)
  wire mux_387_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4570" *)
  wire mux_388_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4268" *)
  wire mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4574" *)
  wire mux_392_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4573" *)
  wire mux_393_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4569" *)
  wire mux_394_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4578" *)
  wire mux_398_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4577" *)
  wire mux_399_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4197" *)
  wire mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6642" *)
  wire mux_404_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4580" *)
  wire mux_406_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4579" *)
  wire mux_407_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4576" *)
  wire mux_408_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4273" *)
  wire mux_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3770" *)
  wire mux_417_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4584" *)
  wire mux_418_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4272" *)
  wire mux_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4589" *)
  wire mux_423_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4588" *)
  wire mux_424_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4592" *)
  wire mux_429_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4276" *)
  wire mux_42_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4591" *)
  wire mux_430_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4587" *)
  wire mux_431_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4596" *)
  wire mux_436_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4595" *)
  wire mux_437_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4280" *)
  wire mux_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4598" *)
  wire mux_442_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4597" *)
  wire mux_443_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4594" *)
  wire mux_444_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5811" *)
  wire mux_449_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4279" *)
  wire mux_44_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4606" *)
  wire mux_450_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4607" *)
  wire mux_453_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5813" *)
  wire mux_454_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4609" *)
  wire mux_456_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4608" *)
  wire mux_458_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4283" *)
  wire mux_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4613" *)
  wire mux_461_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4612" *)
  wire mux_462_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4615" *)
  wire mux_465_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4614" *)
  wire mux_466_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4611" *)
  wire mux_467_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4287" *)
  wire mux_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4618" *)
  wire mux_471_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4617" *)
  wire mux_472_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2727" *)
  wire mux_474_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4622" *)
  wire mux_477_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4620" *)
  wire mux_478_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4286" *)
  wire mux_47_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4626" *)
  wire mux_482_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4625" *)
  wire mux_483_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6660" *)
  wire mux_486_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4629" *)
  wire mux_488_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4628" *)
  wire mux_489_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4292" *)
  wire mux_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4624" *)
  wire mux_490_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4633" *)
  wire mux_494_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4632" *)
  wire mux_495_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4291" *)
  wire mux_49_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4196" *)
  wire mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6663" *)
  wire mux_500_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4635" *)
  wire mux_503_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4634" *)
  wire mux_504_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4631" *)
  wire mux_505_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4294" *)
  wire mux_50_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4642" *)
  wire mux_515_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4640" *)
  wire mux_516_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4298" *)
  wire mux_51_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4646" *)
  wire mux_520_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4645" *)
  wire mux_521_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6668" *)
  wire mux_524_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4649" *)
  wire mux_526_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4648" *)
  wire mux_527_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4644" *)
  wire mux_528_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4297" *)
  wire mux_52_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4653" *)
  wire mux_532_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4652" *)
  wire mux_533_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6672" *)
  wire mux_538_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4303" *)
  wire mux_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6671" *)
  wire mux_540_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4655" *)
  wire mux_542_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4654" *)
  wire mux_543_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4651" *)
  wire mux_544_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4302" *)
  wire mux_54_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4662" *)
  wire mux_555_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4659" *)
  wire mux_556_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4306" *)
  wire mux_55_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4666" *)
  wire mux_561_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4665" *)
  wire mux_562_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4669" *)
  wire mux_567_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4668" *)
  wire mux_568_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4664" *)
  wire mux_569_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4305" *)
  wire mux_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4673" *)
  wire mux_574_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4672" *)
  wire mux_575_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6679" *)
  wire mux_576_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4311" *)
  wire mux_57_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4675" *)
  wire mux_581_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4674" *)
  wire mux_582_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4671" *)
  wire mux_583_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4310" *)
  wire mux_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4687" *)
  wire mux_593_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4684" *)
  wire mux_594_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4691" *)
  wire mux_598_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4690" *)
  wire mux_599_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4316" *)
  wire mux_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4188" *)
  wire mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4694" *)
  wire mux_603_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4693" *)
  wire mux_604_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4689" *)
  wire mux_605_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4698" *)
  wire mux_609_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4315" *)
  wire mux_60_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4697" *)
  wire mux_610_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6692" *)
  wire mux_611_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4701" *)
  wire mux_615_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4700" *)
  wire mux_616_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4696" *)
  wire mux_617_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4319" *)
  wire mux_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4711" *)
  wire mux_629_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4323" *)
  wire mux_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4708" *)
  wire mux_630_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4715" *)
  wire mux_635_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4714" *)
  wire mux_636_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6698" *)
  wire mux_637_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4322" *)
  wire mux_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4718" *)
  wire mux_642_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4717" *)
  wire mux_643_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4713" *)
  wire mux_644_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4328" *)
  wire mux_64_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4327" *)
  wire mux_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2731" *)
  wire mux_660_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4330" *)
  wire mux_66_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4742" *)
  wire mux_670_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4739" *)
  wire mux_671_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4746" *)
  wire mux_676_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4745" *)
  wire mux_677_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4334" *)
  wire mux_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4749" *)
  wire mux_682_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4748" *)
  wire mux_683_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4744" *)
  wire mux_684_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4753" *)
  wire mux_689_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4333" *)
  wire mux_68_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4752" *)
  wire mux_690_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6710" *)
  wire mux_691_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4755" *)
  wire mux_696_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4754" *)
  wire mux_697_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4751" *)
  wire mux_698_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4339" *)
  wire mux_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4338" *)
  wire mux_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4770" *)
  wire mux_714_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4767" *)
  wire mux_715_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4342" *)
  wire mux_71_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4774" *)
  wire mux_721_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4773" *)
  wire mux_722_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4777" *)
  wire mux_728_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4776" *)
  wire mux_729_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4341" *)
  wire mux_72_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4772" *)
  wire mux_730_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4781" *)
  wire mux_736_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4780" *)
  wire mux_737_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6723" *)
  wire mux_738_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4347" *)
  wire mux_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4784" *)
  wire mux_744_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4783" *)
  wire mux_745_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4779" *)
  wire mux_746_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4346" *)
  wire mux_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4352" *)
  wire mux_75_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2738" *)
  wire mux_767_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4351" *)
  wire mux_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5815" *)
  wire mux_770_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4355" *)
  wire mux_77_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3762" *)
  wire mux_786_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5817" *)
  wire mux_789_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4359" *)
  wire mux_78_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4801" *)
  wire mux_792_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4802" *)
  wire mux_793_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4800" *)
  wire mux_794_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4804" *)
  wire mux_796_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5820" *)
  wire mux_798_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5819" *)
  wire mux_799_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4358" *)
  wire mux_79_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4204" *)
  wire mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4805" *)
  wire mux_800_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5823" *)
  wire mux_801_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5825" *)
  wire mux_802_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5822" *)
  wire mux_803_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4810" *)
  wire mux_805_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4812" *)
  wire mux_806_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4809" *)
  wire mux_807_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4816" *)
  wire mux_808_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4818" *)
  wire mux_809_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4364" *)
  wire mux_80_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4815" *)
  wire mux_810_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4808" *)
  wire mux_811_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4822" *)
  wire mux_812_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2688" *)
  wire mux_813_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4825" *)
  wire mux_814_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4820" *)
  wire mux_815_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4828" *)
  wire mux_816_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4830" *)
  wire mux_817_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4827" *)
  wire mux_818_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4836" *)
  wire mux_819_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4363" *)
  wire mux_81_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4839" *)
  wire mux_821_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4834" *)
  wire mux_822_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4845" *)
  wire mux_823_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4844" *)
  wire mux_825_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4843" *)
  wire mux_826_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2690" *)
  wire mux_827_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4850" *)
  wire mux_828_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4841" *)
  wire mux_829_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4366" *)
  wire mux_82_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4872" *)
  wire mux_830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4875" *)
  wire mux_832_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4870" *)
  wire mux_833_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4890" *)
  wire mux_834_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4893" *)
  wire mux_836_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4888" *)
  wire mux_837_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4911" *)
  wire mux_838_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4370" *)
  wire mux_83_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4914" *)
  wire mux_840_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4909" *)
  wire mux_841_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4921" *)
  wire mux_842_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4920" *)
  wire mux_843_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4924" *)
  wire mux_844_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4919" *)
  wire mux_845_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4928" *)
  wire mux_846_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4930" *)
  wire mux_847_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4927" *)
  wire mux_848_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4918" *)
  wire mux_849_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4369" *)
  wire mux_84_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4934" *)
  wire mux_850_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4937" *)
  wire mux_852_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4932" *)
  wire mux_853_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4947" *)
  wire mux_854_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4946" *)
  wire mux_855_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4945" *)
  wire mux_856_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4950" *)
  wire mux_857_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4949" *)
  wire mux_858_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4944" *)
  wire mux_859_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4375" *)
  wire mux_85_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4968" *)
  wire mux_860_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4971" *)
  wire mux_862_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4966" *)
  wire mux_863_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4977" *)
  wire mux_864_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4980" *)
  wire mux_866_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4975" *)
  wire mux_867_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4995" *)
  wire mux_868_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4994" *)
  wire mux_869_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4374" *)
  wire mux_86_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4998" *)
  wire mux_870_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4993" *)
  wire mux_871_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5002" *)
  wire mux_872_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5004" *)
  wire mux_873_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5001" *)
  wire mux_874_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4992" *)
  wire mux_875_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5017" *)
  wire mux_876_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5020" *)
  wire mux_878_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5015" *)
  wire mux_879_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4377" *)
  wire mux_87_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5029" *)
  wire mux_880_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5028" *)
  wire mux_881_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5032" *)
  wire mux_882_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5027" *)
  wire mux_883_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5036" *)
  wire mux_884_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5038" *)
  wire mux_885_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5035" *)
  wire mux_886_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5026" *)
  wire mux_887_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5042" *)
  wire mux_888_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4381" *)
  wire mux_88_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5045" *)
  wire mux_890_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5040" *)
  wire mux_891_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5052" *)
  wire mux_892_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5050" *)
  wire mux_894_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5049" *)
  wire mux_895_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5058" *)
  wire mux_897_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5056" *)
  wire mux_898_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5047" *)
  wire mux_899_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4380" *)
  wire mux_89_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4202" *)
  wire mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5073" *)
  wire mux_902_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5075" *)
  wire mux_903_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5072" *)
  wire mux_904_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5069" *)
  wire mux_906_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5079" *)
  wire mux_908_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5067" *)
  wire mux_909_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4386" *)
  wire mux_90_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5097" *)
  wire mux_910_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5100" *)
  wire mux_912_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5095" *)
  wire mux_913_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5109" *)
  wire mux_914_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5108" *)
  wire mux_915_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5112" *)
  wire mux_916_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5107" *)
  wire mux_917_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5117" *)
  wire mux_918_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5120" *)
  wire mux_919_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4385" *)
  wire mux_91_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5116" *)
  wire mux_920_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5106" *)
  wire mux_921_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5123" *)
  wire mux_922_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5126" *)
  wire mux_924_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5121" *)
  wire mux_925_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5148" *)
  wire mux_926_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5151" *)
  wire mux_928_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5146" *)
  wire mux_929_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5824" *)
  wire mux_92_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5155" *)
  wire mux_930_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5158" *)
  wire mux_932_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5153" *)
  wire mux_933_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5178" *)
  wire mux_934_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5181" *)
  wire mux_936_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5176" *)
  wire mux_937_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5192" *)
  wire mux_938_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5196" *)
  wire mux_939_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5194" *)
  wire mux_940_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5193" *)
  wire mux_943_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5200" *)
  wire mux_948_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5203" *)
  wire mux_949_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5202" *)
  wire mux_950_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5205" *)
  wire mux_951_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5207" *)
  wire mux_952_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5204" *)
  wire mux_953_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5201" *)
  wire mux_954_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5208" *)
  wire mux_959_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5211" *)
  wire mux_964_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6732" *)
  wire mux_969_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6755" *)
  wire mux_976_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5212" *)
  wire mux_982_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5217" *)
  wire mux_984_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5216" *)
  wire mux_985_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5219" *)
  wire mux_988_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3733" *)
  wire mux_989_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5218" *)
  wire mux_990_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5215" *)
  wire mux_991_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5221" *)
  wire mux_995_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4208" *)
  wire mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4185" *)
  wire mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1161" *)
  wire mux_tmp_1015;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1162" *)
  wire mux_tmp_1038;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1164" *)
  wire mux_tmp_1039;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1167" *)
  wire mux_tmp_1041;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1168" *)
  wire mux_tmp_1043;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1169" *)
  wire mux_tmp_1047;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1170" *)
  wire mux_tmp_1049;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1171" *)
  wire mux_tmp_1074;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1172" *)
  wire mux_tmp_1088;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1173" *)
  wire mux_tmp_1100;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1175" *)
  wire mux_tmp_1101;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1178" *)
  wire mux_tmp_1103;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1179" *)
  wire mux_tmp_1105;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1180" *)
  wire mux_tmp_1109;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1181" *)
  wire mux_tmp_1111;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1013" *)
  wire mux_tmp_114;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1182" *)
  wire mux_tmp_1152;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1015" *)
  wire mux_tmp_117;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1183" *)
  wire mux_tmp_1196;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1184" *)
  wire mux_tmp_1197;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1018" *)
  wire mux_tmp_120;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1022" *)
  wire mux_tmp_122;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1187" *)
  wire mux_tmp_1225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1188" *)
  wire mux_tmp_1226;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1189" *)
  wire mux_tmp_1227;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1023" *)
  wire mux_tmp_123;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1190" *)
  wire mux_tmp_1264;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1193" *)
  wire mux_tmp_1270;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1194" *)
  wire mux_tmp_1276;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1195" *)
  wire mux_tmp_1280;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1196" *)
  wire mux_tmp_1282;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1025" *)
  wire mux_tmp_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1197" *)
  wire mux_tmp_1326;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1198" *)
  wire mux_tmp_1332;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1199" *)
  wire mux_tmp_1337;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1200" *)
  wire mux_tmp_1339;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1201" *)
  wire mux_tmp_1341;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1202" *)
  wire mux_tmp_1409;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1203" *)
  wire mux_tmp_1419;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1206" *)
  wire mux_tmp_1435;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1207" *)
  wire mux_tmp_1469;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1027" *)
  wire mux_tmp_151;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1211" *)
  wire mux_tmp_1566;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1213" *)
  wire mux_tmp_1570;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1215" *)
  wire mux_tmp_1574;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1217" *)
  wire mux_tmp_1578;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1219" *)
  wire mux_tmp_1582;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1221" *)
  wire mux_tmp_1586;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1223" *)
  wire mux_tmp_1592;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1225" *)
  wire mux_tmp_1596;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1227" *)
  wire mux_tmp_1600;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1229" *)
  wire mux_tmp_1606;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1028" *)
  wire mux_tmp_161;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1231" *)
  wire mux_tmp_1610;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1233" *)
  wire mux_tmp_1614;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1235" *)
  wire mux_tmp_1618;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1237" *)
  wire mux_tmp_1622;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1287" *)
  wire mux_tmp_1813;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1030" *)
  wire mux_tmp_189;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1310" *)
  wire mux_tmp_1899;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1032" *)
  wire mux_tmp_199;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1033" *)
  wire mux_tmp_200;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2607" *)
  wire mux_tmp_2203;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2609" *)
  wire mux_tmp_2206;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3536" *)
  wire mux_tmp_2294;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3538" *)
  wire mux_tmp_2298;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3539" *)
  wire mux_tmp_2300;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3541" *)
  wire mux_tmp_2304;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3542" *)
  wire mux_tmp_2306;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3544" *)
  wire mux_tmp_2310;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3545" *)
  wire mux_tmp_2312;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3547" *)
  wire mux_tmp_2315;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3548" *)
  wire mux_tmp_2317;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3549" *)
  wire mux_tmp_2319;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3551" *)
  wire mux_tmp_2322;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3552" *)
  wire mux_tmp_2324;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3554" *)
  wire mux_tmp_2328;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3555" *)
  wire mux_tmp_2330;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3556" *)
  wire mux_tmp_2334;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3557" *)
  wire mux_tmp_2336;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3559" *)
  wire mux_tmp_2339;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3560" *)
  wire mux_tmp_2341;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3562" *)
  wire mux_tmp_2345;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3563" *)
  wire mux_tmp_2347;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3565" *)
  wire mux_tmp_2351;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3566" *)
  wire mux_tmp_2353;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1035" *)
  wire mux_tmp_236;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1036" *)
  wire mux_tmp_239;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1037" *)
  wire mux_tmp_245;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1040" *)
  wire mux_tmp_249;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1041" *)
  wire mux_tmp_251;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1042" *)
  wire mux_tmp_253;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1043" *)
  wire mux_tmp_259;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1044" *)
  wire mux_tmp_263;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1049" *)
  wire mux_tmp_294;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1050" *)
  wire mux_tmp_298;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1051" *)
  wire mux_tmp_299;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1052" *)
  wire mux_tmp_305;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1054" *)
  wire mux_tmp_309;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1055" *)
  wire mux_tmp_311;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1056" *)
  wire mux_tmp_313;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1057" *)
  wire mux_tmp_317;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1059" *)
  wire mux_tmp_321;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1062" *)
  wire mux_tmp_345;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1063" *)
  wire mux_tmp_351;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1064" *)
  wire mux_tmp_356;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1065" *)
  wire mux_tmp_370;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1068" *)
  wire mux_tmp_386;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1010" *)
  wire mux_tmp_39;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1069" *)
  wire mux_tmp_391;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1070" *)
  wire mux_tmp_405;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1072" *)
  wire mux_tmp_415;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1073" *)
  wire mux_tmp_416;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1074" *)
  wire mux_tmp_421;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1075" *)
  wire mux_tmp_422;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1076" *)
  wire mux_tmp_427;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1077" *)
  wire mux_tmp_428;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1078" *)
  wire mux_tmp_435;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1079" *)
  wire mux_tmp_440;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1080" *)
  wire mux_tmp_441;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1083" *)
  wire mux_tmp_455;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1086" *)
  wire mux_tmp_481;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1087" *)
  wire mux_tmp_487;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1088" *)
  wire mux_tmp_502;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1090" *)
  wire mux_tmp_519;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1091" *)
  wire mux_tmp_525;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1092" *)
  wire mux_tmp_541;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1094" *)
  wire mux_tmp_560;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1095" *)
  wire mux_tmp_565;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1096" *)
  wire mux_tmp_566;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1097" *)
  wire mux_tmp_577;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1098" *)
  wire mux_tmp_578;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1099" *)
  wire mux_tmp_579;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1100" *)
  wire mux_tmp_580;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1101" *)
  wire mux_tmp_585;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1102" *)
  wire mux_tmp_591;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1103" *)
  wire mux_tmp_592;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1104" *)
  wire mux_tmp_597;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1008" *)
  wire mux_tmp_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1105" *)
  wire mux_tmp_600;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1106" *)
  wire mux_tmp_601;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1107" *)
  wire mux_tmp_602;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1108" *)
  wire mux_tmp_612;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1109" *)
  wire mux_tmp_613;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1110" *)
  wire mux_tmp_614;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1112" *)
  wire mux_tmp_634;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1113" *)
  wire mux_tmp_638;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1114" *)
  wire mux_tmp_639;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1115" *)
  wire mux_tmp_640;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1116" *)
  wire mux_tmp_641;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1118" *)
  wire mux_tmp_658;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1119" *)
  wire mux_tmp_678;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1120" *)
  wire mux_tmp_679;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1121" *)
  wire mux_tmp_680;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1122" *)
  wire mux_tmp_681;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1123" *)
  wire mux_tmp_692;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1124" *)
  wire mux_tmp_693;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1125" *)
  wire mux_tmp_694;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1126" *)
  wire mux_tmp_695;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1128" *)
  wire mux_tmp_719;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1129" *)
  wire mux_tmp_720;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1130" *)
  wire mux_tmp_723;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1131" *)
  wire mux_tmp_724;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1132" *)
  wire mux_tmp_725;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1133" *)
  wire mux_tmp_726;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1134" *)
  wire mux_tmp_727;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1135" *)
  wire mux_tmp_739;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1136" *)
  wire mux_tmp_740;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1137" *)
  wire mux_tmp_741;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1138" *)
  wire mux_tmp_742;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1139" *)
  wire mux_tmp_743;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1141" *)
  wire mux_tmp_765;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1142" *)
  wire mux_tmp_766;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1145" *)
  wire mux_tmp_944;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1146" *)
  wire mux_tmp_945;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1148" *)
  wire mux_tmp_946;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1149" *)
  wire mux_tmp_947;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1151" *)
  wire mux_tmp_960;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1152" *)
  wire mux_tmp_961;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1154" *)
  wire mux_tmp_962;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1155" *)
  wire mux_tmp_963;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1157" *)
  wire mux_tmp_986;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1158" *)
  wire mux_tmp_987;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1159" *)
  wire mux_tmp_992;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1160" *)
  wire mux_tmp_994;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4972" *)
  wire nand_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4981" *)
  wire nand_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2553" *)
  wire nand_133_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2552" *)
  wire nand_135_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2551" *)
  wire nand_137_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2550" *)
  wire nand_139_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5021" *)
  wire nand_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2549" *)
  wire nand_141_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2548" *)
  wire nand_143_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2547" *)
  wire nand_145_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2546" *)
  wire nand_147_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2545" *)
  wire nand_149_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2544" *)
  wire nand_151_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2543" *)
  wire nand_153_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2542" *)
  wire nand_156_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2541" *)
  wire nand_158_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5046" *)
  wire nand_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2540" *)
  wire nand_160_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2539" *)
  wire nand_162_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2538" *)
  wire nand_164_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5051" *)
  wire nand_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3725" *)
  wire nand_171_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5053" *)
  wire nand_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2537" *)
  wire nand_190_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5426" *)
  wire nand_199_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5421" *)
  wire nand_201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2737" *)
  wire nand_202_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5037" *)
  wire nand_204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5003" *)
  wire nand_205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4929" *)
  wire nand_206_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2689" *)
  wire nand_207_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4817" *)
  wire nand_208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2501" *)
  wire nand_219_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5101" *)
  wire nand_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4728" *)
  wire nand_225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5119" *)
  wire nand_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6801" *)
  wire nand_230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4353" *)
  wire nand_231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4317" *)
  wire nand_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4281" *)
  wire nand_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4270" *)
  wire nand_234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4256" *)
  wire nand_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5127" *)
  wire nand_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5152" *)
  wire nand_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5159" *)
  wire nand_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5182" *)
  wire nand_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4826" *)
  wire nand_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4840" *)
  wire nand_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5418" *)
  wire nand_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5423" *)
  wire nand_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4847" *)
  wire nand_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4707" *)
  wire nand_51_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4876" *)
  wire nand_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4894" *)
  wire nand_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4915" *)
  wire nand_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4938" *)
  wire nand_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6594" *)
  wire nand_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1163" *)
  wire nand_tmp_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1174" *)
  wire nand_tmp_36;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1205" *)
  wire nand_tmp_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3243" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3246" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3249" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3252" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3255" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3258" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2714" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3219" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3222" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3225" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3228" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3231" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3234" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3237" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3240" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3261" *)
  (* unused_bits = "16" *)
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3361" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3363" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3365" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3367" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3369" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3371" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3343" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3345" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3347" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3349" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3351" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3353" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3355" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3357" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3359" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3373" *)
  (* unused_bits = "17" *)
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1734" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1740" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2;
  wire [4:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2377" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2373" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2369" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2365" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2361" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2357" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2413" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2409" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2405" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2401" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2397" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2393" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2389" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2385" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2381" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2353" *)
  (* unused_bits = "11" *)
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2958" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2960" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2962" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2964" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2966" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2968" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2970" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2972" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2942" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2944" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2946" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2948" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2950" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2952" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2954" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2956" *)
  (* unused_bits = "3" *)
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2443" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2441" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2439" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2437" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2435" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2433" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2461" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2459" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2457" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2455" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2453" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2451" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2449" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2447" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2445" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2431" *)
  (* unused_bits = "45" *)
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7261" *)
  wire [271:0] nl_NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_inst_chn_out_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6202" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire [4:0] nl_cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6427" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5369" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7062" *)
  wire [16:0] nl_cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7204" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  wire [22:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7201" *)
  wire [3:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6533" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6239" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_10_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6075" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_10_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5972" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5932" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:969" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5934" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6571" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6354" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_10_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6477" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4807" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_10_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5514" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6311" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6875" *)
  wire [111:0] nl_cvt_10_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:871" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [40:0] nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6959" *)
  wire [5:0] nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4408" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7066" *)
  wire [16:0] nl_cvt_10_leading_sign_17_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6205" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire [4:0] nl_cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6429" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5381" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7070" *)
  wire [16:0] nl_cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7213" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  wire [22:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7210" *)
  wire [3:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6536" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6245" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_11_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6084" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_11_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5970" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5936" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:966" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5938" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6573" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6357" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_11_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6481" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5184" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_11_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5511" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6315" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6881" *)
  wire [111:0] nl_cvt_11_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:866" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [40:0] nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6965" *)
  wire [5:0] nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4414" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7074" *)
  wire [16:0] nl_cvt_11_leading_sign_17_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6199" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire [4:0] nl_cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6431" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5400" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7078" *)
  wire [16:0] nl_cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7222" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  wire [22:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7219" *)
  wire [3:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6539" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6251" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_12_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6093" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_12_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5968" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5940" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:963" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5942" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6575" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6359" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_12_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6485" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5191" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_12_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5508" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6313" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6878" *)
  wire [111:0] nl_cvt_12_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:861" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [40:0] nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6971" *)
  wire [5:0] nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4411" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7082" *)
  wire [16:0] nl_cvt_12_leading_sign_17_0_3_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6191" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire [4:0] nl_cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6433" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5408" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7086" *)
  wire [16:0] nl_cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7231" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  wire [22:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7228" *)
  wire [3:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6542" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6257" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_13_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6102" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_13_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5966" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5944" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:960" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5946" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6577" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6363" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_13_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6489" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5170" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_13_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5505" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6323" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6893" *)
  wire [111:0] nl_cvt_13_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:856" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [40:0] nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6977" *)
  wire [5:0] nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4430" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7090" *)
  wire [16:0] nl_cvt_13_leading_sign_17_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6185" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire [4:0] nl_cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6435" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5428" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7094" *)
  wire [16:0] nl_cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7240" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  wire [22:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7237" *)
  wire [3:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6545" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6263" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_14_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6111" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_14_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5964" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5948" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:957" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5950" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6583" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6365" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_14_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6503" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5416" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_14_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5502" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6884" *)
  wire [111:0] nl_cvt_14_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:851" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [40:0] nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6983" *)
  wire [5:0] nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4417" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7098" *)
  wire [16:0] nl_cvt_14_leading_sign_17_0_3_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6179" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire [4:0] nl_cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6437" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5437" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7102" *)
  wire [16:0] nl_cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7249" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  wire [22:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7246" *)
  wire [3:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6548" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6269" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_15_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6120" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_15_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5962" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5952" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:954" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5954" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6579" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6368" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_15_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6495" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5135" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_15_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5499" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6321" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6890" *)
  wire [111:0] nl_cvt_15_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:846" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [40:0] nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6989" *)
  wire [5:0] nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4427" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7106" *)
  wire [16:0] nl_cvt_15_leading_sign_17_0_3_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6171" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl;
  wire [4:0] nl_cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6439" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5445" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7110" *)
  wire [16:0] nl_cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7258" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg_s;
  wire [22:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7255" *)
  wire [3:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6551" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6275" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_16_FpMantRNE_17U_11U_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6129" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_16_FpMantRNE_24U_11U_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5960" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5956" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:951" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5958" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6581" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6370" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_16_IntSaturation_17U_16U_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6499" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5066" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_16_IntSaturation_17U_8U_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5464" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6319" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6887" *)
  wire [111:0] nl_cvt_16_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_4_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:841" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp;
  wire [40:0] nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_a;
  wire [2:0] nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4420" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7114" *)
  wire [16:0] nl_cvt_16_leading_sign_17_0_4_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6152" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl;
  wire [4:0] nl_cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6409" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5238" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6998" *)
  wire [16:0] nl_cvt_1_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7123" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s;
  wire [22:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7120" *)
  wire [3:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6506" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5475" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_1_FpMantRNE_17U_11U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5994" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_1_FpMantRNE_24U_11U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5990" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5896" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:997" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5898" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6553" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_1_IntSaturation_17U_16U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6329" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_1_IntSaturation_17U_16U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6441" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_1_IntSaturation_17U_8U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6177" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_1_IntSaturation_17U_8U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5541" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6327" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6899" *)
  wire [111:0] nl_cvt_1_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:916" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp;
  wire [40:0] nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6905" *)
  wire [5:0] nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4434" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_1_IntSubExt_32U_32U_33U_o_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7001" *)
  wire [16:0] nl_cvt_1_leading_sign_17_0_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6155" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire [4:0] nl_cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6411" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5259" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7004" *)
  wire [16:0] nl_cvt_2_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7132" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  wire [22:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7129" *)
  wire [3:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6509" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4855" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_2_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6003" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_2_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5988" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5900" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:994" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5902" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6555" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6331" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_2_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6445" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4833" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_2_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5538" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6297" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6854" *)
  wire [111:0] nl_cvt_2_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:911" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [40:0] nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6911" *)
  wire [5:0] nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4389" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7007" *)
  wire [16:0] nl_cvt_2_leading_sign_17_0_1_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6160" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire [4:0] nl_cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6413" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5276" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7010" *)
  wire [16:0] nl_cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7141" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  wire [22:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7138" *)
  wire [3:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6512" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5268" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_3_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6012" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_3_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5986" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5904" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:991" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5906" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6557" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6334" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_3_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6449" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6158" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_3_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5535" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6301" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6860" *)
  wire [111:0] nl_cvt_3_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:906" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [40:0] nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6917" *)
  wire [5:0] nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4394" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7013" *)
  wire [16:0] nl_cvt_3_leading_sign_17_0_1_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6163" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire [4:0] nl_cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6415" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5292" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7016" *)
  wire [16:0] nl_cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7150" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  wire [22:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7147" *)
  wire [3:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6515" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6212" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_4_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6021" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_4_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5984" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5908" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:988" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5910" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6559" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6336" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_4_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6453" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4887" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_4_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5532" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6299" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6857" *)
  wire [111:0] nl_cvt_4_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:901" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [40:0] nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  wire [4:0] nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4392" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7020" *)
  wire [16:0] nl_cvt_4_leading_sign_17_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6168" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1931" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6417" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5303" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7024" *)
  wire [16:0] nl_cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7159" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  wire [22:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7156" *)
  wire [3:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6518" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6218" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_5_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6030" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_5_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5982" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5912" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:985" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5914" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6561" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6340" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_5_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6457" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6166" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_5_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5529" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6309" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6872" *)
  wire [111:0] nl_cvt_5_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:896" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [40:0] nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6929" *)
  wire [5:0] nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4405" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7028" *)
  wire [16:0] nl_cvt_5_leading_sign_17_0_1_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6174" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1934" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6419" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5319" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7032" *)
  wire [16:0] nl_cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7168" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  wire [22:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7165" *)
  wire [3:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6521" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6221" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_6_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6039" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_6_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5980" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5916" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:981" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5918" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6563" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6342" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_6_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6461" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4974" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_6_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5526" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6303" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6863" *)
  wire [111:0] nl_cvt_6_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:891" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [40:0] nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6935" *)
  wire [5:0] nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4397" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7036" *)
  wire [16:0] nl_cvt_6_leading_sign_17_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6182" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1937" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6421" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5330" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7040" *)
  wire [16:0] nl_cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7177" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  wire [22:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7174" *)
  wire [3:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6524" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6227" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_7_FpMantRNE_17U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6048" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_7_FpMantRNE_24U_11U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5978" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5920" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:978" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5922" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6565" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6345" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_7_IntSaturation_17U_16U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6465" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5023" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_7_IntSaturation_17U_8U_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5523" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6307" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6869" *)
  wire [111:0] nl_cvt_7_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:886" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [40:0] nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6941" *)
  wire [5:0] nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4403" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7044" *)
  wire [16:0] nl_cvt_7_leading_sign_17_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6188" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1940" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6423" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5345" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7048" *)
  wire [16:0] nl_cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7186" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  wire [22:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7183" *)
  wire [3:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6527" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6233" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_8_FpMantRNE_17U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6057" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_8_FpMantRNE_24U_11U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5976" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5924" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:975" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5926" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6567" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6347" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_8_IntSaturation_17U_16U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6469" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5103" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_8_IntSaturation_17U_8U_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5520" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6305" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6866" *)
  wire [111:0] nl_cvt_8_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:881" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [40:0] nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6947" *)
  wire [5:0] nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4400" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7052" *)
  wire [16:0] nl_cvt_8_leading_sign_17_0_3_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6196" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 12" *)
  wire [12:0] nl_cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1943" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6425" *)
  (* unused_bits = "0 1 2 3 5" *)
  wire [5:0] nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5359" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7056" *)
  wire [16:0] nl_cvt_9_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7195" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  wire [22:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7192" *)
  wire [3:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6530" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5163" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_9_FpMantRNE_17U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6066" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_cvt_9_FpMantRNE_24U_11U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5974" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5928" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:972" *)
  (* unused_bits = "5" *)
  wire [5:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5930" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6569" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6352" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_cvt_9_IntSaturation_17U_16U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6473" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6194" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_cvt_9_IntSaturation_17U_8U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5517" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6325" *)
  (* unused_bits = "18" *)
  wire [18:0] nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6896" *)
  wire [111:0] nl_cvt_9_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:876" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [40:0] nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6953" *)
  wire [5:0] nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4432" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7059" *)
  wire [16:0] nl_cvt_9_leading_sign_17_0_1_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6806" *)
  wire nor_1025_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4982" *)
  wire nor_1033_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4953" *)
  wire nor_1040_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3744" *)
  wire nor_1048_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4899" *)
  wire nor_1049_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6805" *)
  wire nor_1053_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2502" *)
  wire nor_1056_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6802" *)
  wire nor_1063_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2561" *)
  wire nor_1099_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2555" *)
  wire nor_1185_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2556" *)
  wire nor_1186_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5775" *)
  wire nor_1195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5747" *)
  wire nor_1198_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5725" *)
  wire nor_1200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5688" *)
  wire nor_1201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5689" *)
  wire nor_1202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5685" *)
  wire nor_1203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5686" *)
  wire nor_1204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5682" *)
  wire nor_1205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5683" *)
  wire nor_1206_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5679" *)
  wire nor_1207_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5680" *)
  wire nor_1208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5676" *)
  wire nor_1209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5677" *)
  wire nor_1210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5673" *)
  wire nor_1211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5674" *)
  wire nor_1212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5670" *)
  wire nor_1213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5671" *)
  wire nor_1214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5667" *)
  wire nor_1215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5668" *)
  wire nor_1216_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5664" *)
  wire nor_1217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5665" *)
  wire nor_1218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5661" *)
  wire nor_1219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5662" *)
  wire nor_1220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5658" *)
  wire nor_1221_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5659" *)
  wire nor_1222_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5655" *)
  wire nor_1223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5656" *)
  wire nor_1224_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5652" *)
  wire nor_1225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5653" *)
  wire nor_1226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5649" *)
  wire nor_1227_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5650" *)
  wire nor_1228_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5646" *)
  wire nor_1229_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5647" *)
  wire nor_1230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5643" *)
  wire nor_1231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5644" *)
  wire nor_1232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5640" *)
  wire nor_1233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5641" *)
  wire nor_1234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5637" *)
  wire nor_1235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5638" *)
  wire nor_1236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5634" *)
  wire nor_1237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5635" *)
  wire nor_1238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5631" *)
  wire nor_1239_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5632" *)
  wire nor_1240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5628" *)
  wire nor_1241_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5629" *)
  wire nor_1242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5625" *)
  wire nor_1243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5626" *)
  wire nor_1244_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5622" *)
  wire nor_1245_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5623" *)
  wire nor_1246_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5619" *)
  wire nor_1247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5620" *)
  wire nor_1248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5616" *)
  wire nor_1249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5617" *)
  wire nor_1250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5613" *)
  wire nor_1251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5614" *)
  wire nor_1252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5610" *)
  wire nor_1253_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5611" *)
  wire nor_1254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5607" *)
  wire nor_1255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5608" *)
  wire nor_1256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5604" *)
  wire nor_1257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5605" *)
  wire nor_1258_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5601" *)
  wire nor_1259_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5602" *)
  wire nor_1260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5598" *)
  wire nor_1261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5599" *)
  wire nor_1262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5595" *)
  wire nor_1263_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5596" *)
  wire nor_1264_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5584" *)
  wire nor_1271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5579" *)
  wire nor_1287_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5570" *)
  wire nor_1301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5575" *)
  wire nor_1302_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5577" *)
  wire nor_1303_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5566" *)
  wire nor_1305_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5564" *)
  wire nor_1306_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3491" *)
  wire nor_1309_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3500" *)
  wire nor_1310_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5558" *)
  wire nor_1314_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2695" *)
  wire nor_1320_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5458" *)
  wire nor_1338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5455" *)
  wire nor_1351_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6766" *)
  wire nor_1371_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6767" *)
  wire nor_1372_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6768" *)
  wire nor_1373_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6764" *)
  wire nor_1387_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6765" *)
  wire nor_1388_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5397" *)
  wire nor_1403_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5376" *)
  wire nor_1415_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5357" *)
  wire nor_1433_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5352" *)
  wire nor_1434_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6757" *)
  wire nor_1446_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6753" *)
  wire nor_1455_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5314" *)
  wire nor_1463_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6749" *)
  wire nor_1464_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5311" *)
  wire nor_1465_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5313" *)
  wire nor_1466_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3754" *)
  wire nor_1486_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6741" *)
  wire nor_1487_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3722" *)
  wire nor_1488_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3723" *)
  wire nor_1489_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5271" *)
  wire nor_1498_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3721" *)
  wire nor_1500_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5256" *)
  wire nor_1508_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5246" *)
  wire nor_1510_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5248" *)
  wire nor_1511_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5235" *)
  wire nor_1519_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2518" *)
  wire nor_151_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5236" *)
  wire nor_1521_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5227" *)
  wire nor_1523_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5229" *)
  wire nor_1524_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5230" *)
  wire nor_1525_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5223" *)
  wire nor_1526_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5224" *)
  wire nor_1527_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6734" *)
  wire nor_1534_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6735" *)
  wire nor_1535_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5220" *)
  wire nor_1536_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5213" *)
  wire nor_1537_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5214" *)
  wire nor_1538_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6733" *)
  wire nor_1545_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5209" *)
  wire nor_1547_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5210" *)
  wire nor_1548_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5206" *)
  wire nor_1555_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2574" *)
  wire nor_1556_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5195" *)
  wire nor_1557_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5199" *)
  wire nor_1558_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5179" *)
  wire nor_1563_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5156" *)
  wire nor_1566_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5149" *)
  wire nor_1569_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5124" *)
  wire nor_1572_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5110" *)
  wire nor_1574_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5111" *)
  wire nor_1575_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5113" *)
  wire nor_1577_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5114" *)
  wire nor_1578_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5115" *)
  wire nor_1579_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5098" *)
  wire nor_1583_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5070" *)
  wire nor_1584_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5071" *)
  wire nor_1585_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5078" *)
  wire nor_1588_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2531" *)
  wire nor_1589_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5043" *)
  wire nor_1596_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5030" *)
  wire nor_1598_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5031" *)
  wire nor_1599_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5033" *)
  wire nor_1602_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5034" *)
  wire nor_1603_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5018" *)
  wire nor_1608_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4996" *)
  wire nor_1610_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4997" *)
  wire nor_1611_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4999" *)
  wire nor_1614_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5000" *)
  wire nor_1615_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4978" *)
  wire nor_1620_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4969" *)
  wire nor_1623_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2513" *)
  wire nor_1624_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4948" *)
  wire nor_1625_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2571" *)
  wire nor_1626_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4951" *)
  wire nor_1628_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2519" *)
  wire nor_1629_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2514" *)
  wire nor_1630_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4935" *)
  wire nor_1634_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4922" *)
  wire nor_1636_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4923" *)
  wire nor_1637_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4925" *)
  wire nor_1640_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4926" *)
  wire nor_1641_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4912" *)
  wire nor_1646_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4891" *)
  wire nor_1649_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4873" *)
  wire nor_1652_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4842" *)
  wire nor_1653_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4849" *)
  wire nor_1655_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4837" *)
  wire nor_1658_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4829" *)
  wire nor_1659_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4831" *)
  wire nor_1661_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2505" *)
  wire nor_1664_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4823" *)
  wire nor_1665_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2509" *)
  wire nor_1666_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4811" *)
  wire nor_1667_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2511" *)
  wire nor_1669_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4813" *)
  wire nor_1670_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4814" *)
  wire nor_1671_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2503" *)
  wire nor_1672_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4799" *)
  wire nor_1674_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4798" *)
  wire nor_1683_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6730" *)
  wire nor_1685_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6731" *)
  wire nor_1686_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6728" *)
  wire nor_1687_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6729" *)
  wire nor_1689_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4782" *)
  wire nor_1697_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4785" *)
  wire nor_1698_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6724" *)
  wire nor_1699_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6725" *)
  wire nor_1700_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6726" *)
  wire nor_1701_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6727" *)
  wire nor_1702_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4775" *)
  wire nor_1708_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4778" *)
  wire nor_1709_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6719" *)
  wire nor_1711_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6720" *)
  wire nor_1712_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6721" *)
  wire nor_1713_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6722" *)
  wire nor_1714_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6716" *)
  wire nor_1718_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6717" *)
  wire nor_1719_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6714" *)
  wire nor_1728_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6715" *)
  wire nor_1730_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4756" *)
  wire nor_1737_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6711" *)
  wire nor_1738_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6712" *)
  wire nor_1739_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6713" *)
  wire nor_1740_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4747" *)
  wire nor_1745_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4750" *)
  wire nor_1746_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6707" *)
  wire nor_1748_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6708" *)
  wire nor_1749_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6709" *)
  wire nor_1750_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4738" *)
  wire nor_1761_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6705" *)
  wire nor_1762_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6703" *)
  wire nor_1764_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6704" *)
  wire nor_1766_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3716" *)
  wire nor_1772_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4719" *)
  wire nor_1773_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6700" *)
  wire nor_1774_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6701" *)
  wire nor_1775_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6702" *)
  wire nor_1776_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6697" *)
  wire nor_1780_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6695" *)
  wire nor_1787_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6696" *)
  wire nor_1789_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4699" *)
  wire nor_1793_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4702" *)
  wire nor_1794_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6693" *)
  wire nor_1795_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6694" *)
  wire nor_1796_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4692" *)
  wire nor_1800_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4695" *)
  wire nor_1801_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6690" *)
  wire nor_1803_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6691" *)
  wire nor_1804_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6688" *)
  wire nor_1807_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4688" *)
  wire nor_1809_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6687" *)
  wire nor_1810_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4676" *)
  wire nor_1814_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6681" *)
  wire nor_1815_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6682" *)
  wire nor_1816_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6683" *)
  wire nor_1817_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4667" *)
  wire nor_1822_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4670" *)
  wire nor_1823_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6678" *)
  wire nor_1827_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6675" *)
  wire nor_1828_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6673" *)
  wire nor_1838_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2528" *)
  wire nor_183_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6674" *)
  wire nor_1840_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4647" *)
  wire nor_1847_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4650" *)
  wire nor_1848_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6667" *)
  wire nor_1851_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6665" *)
  wire nor_1858_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6666" *)
  wire nor_1860_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4627" *)
  wire nor_1868_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4630" *)
  wire nor_1869_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6659" *)
  wire nor_1872_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4619" *)
  wire nor_1875_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6657" *)
  wire nor_1882_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6658" *)
  wire nor_1884_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6656" *)
  wire nor_1891_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6654" *)
  wire nor_1892_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6655" *)
  wire nor_1894_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3769" *)
  wire nor_1898_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6652" *)
  wire nor_1901_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6653" *)
  wire nor_1902_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6651" *)
  wire nor_1906_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4590" *)
  wire nor_1907_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4593" *)
  wire nor_1908_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6650" *)
  wire nor_1911_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6646" *)
  wire nor_1912_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6647" *)
  wire nor_1915_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4583" *)
  wire nor_1917_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6645" *)
  wire nor_1919_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6643" *)
  wire nor_1922_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6644" *)
  wire nor_1924_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4572" *)
  wire nor_1931_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4575" *)
  wire nor_1932_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6639" *)
  wire nor_1935_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4565" *)
  wire nor_1939_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6637" *)
  wire nor_1942_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6638" *)
  wire nor_1944_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4549" *)
  wire nor_1951_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4552" *)
  wire nor_1952_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6633" *)
  wire nor_1955_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4541" *)
  wire nor_1958_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6632" *)
  wire nor_1959_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4539" *)
  wire nor_1962_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6630" *)
  wire nor_1964_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6631" *)
  wire nor_1966_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6629" *)
  wire nor_1974_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6627" *)
  wire nor_1975_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6628" *)
  wire nor_1977_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3715" *)
  wire nor_1980_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6623" *)
  wire nor_1983_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4499" *)
  wire nor_1984_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4502" *)
  wire nor_1985_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6620" *)
  wire nor_1987_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6619" *)
  wire nor_1988_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4495" *)
  wire nor_1991_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4489" *)
  wire nor_1992_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4490" *)
  wire nor_1993_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6617" *)
  wire nor_1995_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6618" *)
  wire nor_1997_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3504" *)
  wire nor_2004_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3505" *)
  wire nor_2005_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6615" *)
  wire nor_2007_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6616" *)
  wire nor_2009_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3503" *)
  wire nor_2011_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6614" *)
  wire nor_2013_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6613" *)
  wire nor_2015_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4459" *)
  wire nor_2016_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4460" *)
  wire nor_2017_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4453" *)
  wire nor_2020_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6602" *)
  wire nor_2021_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6601" *)
  wire nor_2022_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4445" *)
  wire nor_2026_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6599" *)
  wire nor_2027_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6600" *)
  wire nor_2028_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6596" *)
  wire nor_2029_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2494" *)
  wire nor_2040_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4438" *)
  wire nor_2046_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3711" *)
  wire nor_2047_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4436" *)
  wire nor_2048_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6593" *)
  wire nor_2049_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6592" *)
  wire nor_2050_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6590" *)
  wire nor_2052_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6589" *)
  wire nor_2054_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6588" *)
  wire nor_2055_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6587" *)
  wire nor_2056_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4378" *)
  wire nor_2057_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4379" *)
  wire nor_2058_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4367" *)
  wire nor_2059_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4368" *)
  wire nor_2060_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4356" *)
  wire nor_2061_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4357" *)
  wire nor_2062_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4331" *)
  wire nor_2063_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4332" *)
  wire nor_2064_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4320" *)
  wire nor_2065_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4321" *)
  wire nor_2066_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4295" *)
  wire nor_2067_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4296" *)
  wire nor_2068_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4284" *)
  wire nor_2069_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4285" *)
  wire nor_2070_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4234" *)
  wire nor_2071_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4235" *)
  wire nor_2072_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4223" *)
  wire nor_2073_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4224" *)
  wire nor_2074_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4211" *)
  wire nor_2075_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4212" *)
  wire nor_2076_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4186" *)
  wire nor_2081_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4187" *)
  wire nor_2082_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2691" *)
  wire nor_2099_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4865" *)
  wire nor_2100_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4867" *)
  wire nor_2101_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5582" *)
  wire nor_2110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5573" *)
  wire nor_2113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5569" *)
  wire nor_2114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5578" *)
  wire nor_2127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5565" *)
  wire nor_2130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3492" *)
  wire nor_213_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5011" *)
  wire nor_2142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5013" *)
  wire nor_2143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3525" *)
  wire nor_2150_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2725" *)
  wire nor_2219_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5495" *)
  wire nor_2251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5497" *)
  wire nor_2252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5091" *)
  wire nor_2269_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4884" *)
  wire nor_2284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2722" *)
  wire nor_2285_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4797" *)
  wire nor_2287_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4766" *)
  wire nor_2290_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4683" *)
  wire nor_2300_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3758" *)
  wire nor_2326_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5451" *)
  wire nor_2396_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5443" *)
  wire nor_2401_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5434" *)
  wire nor_2406_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5414" *)
  wire nor_2411_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5375" *)
  wire nor_2425_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5365" *)
  wire nor_2429_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5351" *)
  wire nor_2433_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5336" *)
  wire nor_2437_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5325" *)
  wire nor_2441_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5309" *)
  wire nor_2445_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5298" *)
  wire nor_2449_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5282" *)
  wire nor_2453_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5265" *)
  wire nor_2457_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5244" *)
  wire nor_2461_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2594" *)
  wire nor_45_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2495" *)
  wire nor_50_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2563" *)
  wire nor_57_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2526" *)
  wire nor_63_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2534" *)
  wire nor_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1257" *)
  wire nor_tmp_636;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1019" *)
  wire not_tmp_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1204" *)
  wire not_tmp_1709;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1260" *)
  wire not_tmp_2254;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1302" *)
  wire not_tmp_2422;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1045" *)
  wire not_tmp_249;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1046" *)
  wire not_tmp_269;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1047" *)
  wire not_tmp_270;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1058" *)
  wire not_tmp_312;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1061" *)
  wire not_tmp_336;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1066" *)
  wire not_tmp_388;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1071" *)
  wire not_tmp_436;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1081" *)
  wire not_tmp_497;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1085" *)
  wire not_tmp_520;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1089" *)
  wire not_tmp_580;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1093" *)
  wire not_tmp_638;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1111" *)
  wire not_tmp_757;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1117" *)
  wire not_tmp_811;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1127" *)
  wire not_tmp_899;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1140" *)
  wire not_tmp_989;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:689" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:690" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3860" *)
  wire oWidth_aWidth_bWidth_prb;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3864" *)
  wire oWidth_aWidth_bWidth_prb_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3900" *)
  wire oWidth_aWidth_bWidth_prb_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3904" *)
  wire oWidth_aWidth_bWidth_prb_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3908" *)
  wire oWidth_aWidth_bWidth_prb_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3912" *)
  wire oWidth_aWidth_bWidth_prb_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3916" *)
  wire oWidth_aWidth_bWidth_prb_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3920" *)
  wire oWidth_aWidth_bWidth_prb_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3868" *)
  wire oWidth_aWidth_bWidth_prb_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3872" *)
  wire oWidth_aWidth_bWidth_prb_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3876" *)
  wire oWidth_aWidth_bWidth_prb_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3880" *)
  wire oWidth_aWidth_bWidth_prb_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3884" *)
  wire oWidth_aWidth_bWidth_prb_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3888" *)
  wire oWidth_aWidth_bWidth_prb_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3892" *)
  wire oWidth_aWidth_bWidth_prb_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3896" *)
  wire oWidth_aWidth_bWidth_prb_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3859" *)
  wire oWidth_mWidth_prb;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3863" *)
  wire oWidth_mWidth_prb_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3899" *)
  wire oWidth_mWidth_prb_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3903" *)
  wire oWidth_mWidth_prb_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3907" *)
  wire oWidth_mWidth_prb_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3911" *)
  wire oWidth_mWidth_prb_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3915" *)
  wire oWidth_mWidth_prb_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3919" *)
  wire oWidth_mWidth_prb_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3867" *)
  wire oWidth_mWidth_prb_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3871" *)
  wire oWidth_mWidth_prb_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3875" *)
  wire oWidth_mWidth_prb_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3879" *)
  wire oWidth_mWidth_prb_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3883" *)
  wire oWidth_mWidth_prb_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3887" *)
  wire oWidth_mWidth_prb_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3891" *)
  wire oWidth_mWidth_prb_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3895" *)
  wire oWidth_mWidth_prb_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6706" *)
  wire or_1015_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4289" *)
  wire or_101_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4293" *)
  wire or_103_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6718" *)
  wire or_1072_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4300" *)
  wire or_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5816" *)
  wire or_1118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4304" *)
  wire or_111_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5818" *)
  wire or_1134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5821" *)
  wire or_1145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4307" *)
  wire or_114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2507" *)
  wire or_1157_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2512" *)
  wire or_1159_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4308" *)
  wire or_116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2506" *)
  wire or_1176_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2517" *)
  wire or_1196_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3498" *)
  wire or_1198_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4312" *)
  wire or_119_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4193" *)
  wire or_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4846" *)
  wire or_1201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2524" *)
  wire or_1202_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4851" *)
  wire or_1209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4313" *)
  wire or_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4318" *)
  wire or_126_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4952" *)
  wire or_1280_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4325" *)
  wire or_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4329" *)
  wire or_134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5054" *)
  wire or_1374_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5048" *)
  wire or_1375_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5057" *)
  wire or_1379_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5059" *)
  wire or_1383_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5074" *)
  wire or_1393_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5077" *)
  wire or_1396_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5076" *)
  wire or_1399_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4194" *)
  wire or_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5080" *)
  wire or_1402_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5081" *)
  wire or_1409_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4336" *)
  wire or_140_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4340" *)
  wire or_142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5118" *)
  wire or_1431_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4343" *)
  wire or_145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4344" *)
  wire or_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5197" *)
  wire or_1483_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5198" *)
  wire or_1484_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4199" *)
  wire or_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4348" *)
  wire or_150_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4349" *)
  wire or_152_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4354" *)
  wire or_157_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2527" *)
  wire or_1587_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2557" *)
  wire or_1596_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2558" *)
  wire or_1625_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4361" *)
  wire or_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6742" *)
  wire or_1643_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6740" *)
  wire or_1644_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3467" *)
  wire or_1659_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4365" *)
  wire or_165_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2559" *)
  wire or_1693_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4372" *)
  wire or_171_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3468" *)
  wire or_1720_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4376" *)
  wire or_173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6754" *)
  wire or_1745_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3469" *)
  wire or_1752_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6758" *)
  wire or_1773_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6756" *)
  wire or_1774_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3470" *)
  wire or_1789_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4383" *)
  wire or_179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4206" *)
  wire or_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4387" *)
  wire or_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2560" *)
  wire or_1829_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3710" *)
  wire or_183_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3471" *)
  wire or_1851_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3729" *)
  wire or_186_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3472" *)
  wire or_1892_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5398" *)
  wire or_1918_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2575" *)
  wire or_1919_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3473" *)
  wire or_1925_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4203" *)
  wire or_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3734" *)
  wire or_2140_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5879" *)
  wire or_217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6788" *)
  wire or_2232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5557" *)
  wire or_2242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6792" *)
  wire or_2245_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6793" *)
  wire or_2246_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5556" *)
  wire or_2251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5882" *)
  wire or_226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2536" *)
  wire or_2289_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6800" *)
  wire or_2306_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5884" *)
  wire or_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6584" *)
  wire or_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5593" *)
  wire or_2433_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5885" *)
  wire or_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5887" *)
  wire or_263_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5829" *)
  wire or_2688_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5830" *)
  wire or_2691_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5832" *)
  wire or_2696_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5833" *)
  wire or_2699_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5835" *)
  wire or_2705_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5836" *)
  wire or_2709_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5889" *)
  wire or_270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5838" *)
  wire or_2714_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5839" *)
  wire or_2717_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5841" *)
  wire or_2723_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5842" *)
  wire or_2727_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5844" *)
  wire or_2733_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5845" *)
  wire or_2737_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5847" *)
  wire or_2744_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5848" *)
  wire or_2749_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5850" *)
  wire or_2754_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5851" *)
  wire or_2758_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5891" *)
  wire or_275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5853" *)
  wire or_2764_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5854" *)
  wire or_2768_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5856" *)
  wire or_2774_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5857" *)
  wire or_2778_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5859" *)
  wire or_2784_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5860" *)
  wire or_2789_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5862" *)
  wire or_2796_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5863" *)
  wire or_2802_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5865" *)
  wire or_2809_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5866" *)
  wire or_2815_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5868" *)
  wire or_2823_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5869" *)
  wire or_2830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4209" *)
  wire or_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2510" *)
  wire or_300_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3712" *)
  wire or_303_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3529" *)
  wire or_3063_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3714" *)
  wire or_306_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4531" *)
  wire or_3070_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2515" *)
  wire or_309_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3743" *)
  wire or_3151_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4725" *)
  wire or_3170_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4761" *)
  wire or_3196_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4791" *)
  wire or_3220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2572" *)
  wire or_3538_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2573" *)
  wire or_3542_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5479" *)
  wire or_3597_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4217" *)
  wire or_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5485" *)
  wire or_3600_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5487" *)
  wire or_3606_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5490" *)
  wire or_3607_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5492" *)
  wire or_3609_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3724" *)
  wire or_3623_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3735" *)
  wire or_3696_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3756" *)
  wire or_3774_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6597" *)
  wire or_378_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4221" *)
  wire or_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3499" *)
  wire or_3817_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5232" *)
  wire or_3841_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5251" *)
  wire or_3850_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5273" *)
  wire or_3860_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6215" *)
  wire or_3872_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5300" *)
  wire or_3879_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6224" *)
  wire or_3891_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6230" *)
  wire or_3900_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6236" *)
  wire or_3911_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5354" *)
  wire or_3920_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6242" *)
  wire or_3932_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6248" *)
  wire or_3942_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6254" *)
  wire or_3953_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6260" *)
  wire or_3965_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6266" *)
  wire or_3977_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6272" *)
  wire or_3989_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6278" *)
  wire or_3999_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3717" *)
  wire or_400_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2496" *)
  wire or_419_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2497" *)
  wire or_423_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2525" *)
  wire or_425_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6604" *)
  wire or_429_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6605" *)
  wire or_431_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4722" *)
  wire or_4348_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6606" *)
  wire or_434_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4228" *)
  wire or_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6611" *)
  wire or_445_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6607" *)
  wire or_448_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2498" *)
  wire or_451_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2535" *)
  wire or_4524_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5039" *)
  wire or_4526_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5005" *)
  wire or_4528_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4931" *)
  wire or_4530_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4819" *)
  wire or_4532_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2500" *)
  wire or_4535_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2567" *)
  wire or_4536_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2719" *)
  wire or_4550_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3531" *)
  wire or_4559_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4537" *)
  wire or_4569_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4232" *)
  wire or_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3515" *)
  wire or_461_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6831" *)
  wire or_4667_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6834" *)
  wire or_4675_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2721" *)
  wire or_4709_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2724" *)
  wire or_4714_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4885" *)
  wire or_4718_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4962" *)
  wire or_4745_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2739" *)
  wire or_4749_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4965" *)
  wire or_4755_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2740" *)
  wire or_4788_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5094" *)
  wire or_4793_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5807" *)
  wire or_479_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5496" *)
  wire or_4857_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3466" *)
  wire or_4862_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3487" *)
  wire or_5038_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3488" *)
  wire or_5053_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3489" *)
  wire or_5069_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3490" *)
  wire or_5086_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2564" *)
  wire or_510_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2499" *)
  wire or_513_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3581" *)
  wire or_5174_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3580" *)
  wire or_5175_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3579" *)
  wire or_5176_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3578" *)
  wire or_5177_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3577" *)
  wire or_5178_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3576" *)
  wire or_5179_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3575" *)
  wire or_5180_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3574" *)
  wire or_5181_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3573" *)
  wire or_5182_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3572" *)
  wire or_5183_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3571" *)
  wire or_5184_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3570" *)
  wire or_5185_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3569" *)
  wire or_5186_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3568" *)
  wire or_5187_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3567" *)
  wire or_5188_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3583" *)
  wire or_5189_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4239" *)
  wire or_51_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6622" *)
  wire or_520_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3584" *)
  wire or_5254_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3731" *)
  wire or_5379_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4243" *)
  wire or_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5808" *)
  wire or_547_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4246" *)
  wire or_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2593" *)
  wire or_578_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4247" *)
  wire or_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6635" *)
  wire or_599_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2566" *)
  wire or_600_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4251" *)
  wire or_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5810" *)
  wire or_626_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4252" *)
  wire or_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6641" *)
  wire or_645_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4257" *)
  wire or_68_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6649" *)
  wire or_690_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4260" *)
  wire or_71_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5812" *)
  wire or_724_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:5814" *)
  wire or_733_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4261" *)
  wire or_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4265" *)
  wire or_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6662" *)
  wire or_784_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4266" *)
  wire or_78_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6664" *)
  wire or_795_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6670" *)
  wire or_828_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4271" *)
  wire or_83_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6585" *)
  wire or_86_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6677" *)
  wire or_871_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4274" *)
  wire or_88_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6684" *)
  wire or_894_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6685" *)
  wire or_898_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4277" *)
  wire or_90_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6689" *)
  wire or_921_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4282" *)
  wire or_95_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4716" *)
  wire or_961_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:4191" *)
  wire or_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1254" *)
  wire or_dcpl_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1256" *)
  wire or_dcpl_109;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1258" *)
  wire or_dcpl_110;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1259" *)
  wire or_dcpl_111;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1262" *)
  wire or_dcpl_113;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1263" *)
  wire or_dcpl_114;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1265" *)
  wire or_dcpl_115;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1266" *)
  wire or_dcpl_116;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1267" *)
  wire or_dcpl_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1268" *)
  wire or_dcpl_120;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1270" *)
  wire or_dcpl_124;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1271" *)
  wire or_dcpl_125;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1272" *)
  wire or_dcpl_126;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1273" *)
  wire or_dcpl_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1274" *)
  wire or_dcpl_130;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1275" *)
  wire or_dcpl_131;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1276" *)
  wire or_dcpl_132;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1277" *)
  wire or_dcpl_133;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1280" *)
  wire or_dcpl_136;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1282" *)
  wire or_dcpl_137;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1283" *)
  wire or_dcpl_139;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1284" *)
  wire or_dcpl_140;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1285" *)
  wire or_dcpl_143;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1286" *)
  wire or_dcpl_144;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1291" *)
  wire or_dcpl_147;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1246" *)
  wire or_dcpl_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1299" *)
  wire or_dcpl_151;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1247" *)
  wire or_dcpl_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1305" *)
  wire or_dcpl_160;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1308" *)
  wire or_dcpl_163;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1312" *)
  wire or_dcpl_178;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1314" *)
  wire or_dcpl_181;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1315" *)
  wire or_dcpl_184;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1316" *)
  wire or_dcpl_188;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1317" *)
  wire or_dcpl_195;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1318" *)
  wire or_dcpl_197;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1319" *)
  wire or_dcpl_210;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1322" *)
  wire or_dcpl_243;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1326" *)
  wire or_dcpl_277;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1248" *)
  wire or_dcpl_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1249" *)
  wire or_dcpl_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1327" *)
  wire or_dcpl_320;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1328" *)
  wire or_dcpl_322;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1329" *)
  wire or_dcpl_324;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1330" *)
  wire or_dcpl_326;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1331" *)
  wire or_dcpl_328;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1332" *)
  wire or_dcpl_330;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1333" *)
  wire or_dcpl_332;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1334" *)
  wire or_dcpl_334;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1335" *)
  wire or_dcpl_336;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1336" *)
  wire or_dcpl_338;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1337" *)
  wire or_dcpl_340;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1338" *)
  wire or_dcpl_342;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1339" *)
  wire or_dcpl_344;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1340" *)
  wire or_dcpl_346;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1341" *)
  wire or_dcpl_348;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1342" *)
  wire or_dcpl_350;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1343" *)
  wire or_dcpl_353;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1344" *)
  wire or_dcpl_386;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1345" *)
  wire or_dcpl_389;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1347" *)
  wire or_dcpl_399;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1240" *)
  wire or_dcpl_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1350" *)
  wire or_dcpl_420;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1353" *)
  wire or_dcpl_439;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1355" *)
  wire or_dcpl_448;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1359" *)
  wire or_dcpl_480;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1361" *)
  wire or_dcpl_490;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1364" *)
  wire or_dcpl_511;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1369" *)
  wire or_dcpl_612;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3535" *)
  wire or_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1143" *)
  wire or_tmp_1375;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1144" *)
  wire or_tmp_1393;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1166" *)
  wire or_tmp_1650;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1177" *)
  wire or_tmp_1780;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1007" *)
  wire or_tmp_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1185" *)
  wire or_tmp_1981;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1186" *)
  wire or_tmp_1992;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1017" *)
  wire or_tmp_213;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1191" *)
  wire or_tmp_2136;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1192" *)
  wire or_tmp_2139;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1020" *)
  wire or_tmp_218;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1009" *)
  wire or_tmp_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1208" *)
  wire or_tmp_2432;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1209" *)
  wire or_tmp_2466;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1210" *)
  wire or_tmp_2469;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1212" *)
  wire or_tmp_2569;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1214" *)
  wire or_tmp_2571;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1216" *)
  wire or_tmp_2573;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1218" *)
  wire or_tmp_2575;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1220" *)
  wire or_tmp_2577;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1222" *)
  wire or_tmp_2579;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1224" *)
  wire or_tmp_2588;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1226" *)
  wire or_tmp_2590;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1228" *)
  wire or_tmp_2595;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1230" *)
  wire or_tmp_2604;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1232" *)
  wire or_tmp_2606;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1234" *)
  wire or_tmp_2608;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1236" *)
  wire or_tmp_2610;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1238" *)
  wire or_tmp_2612;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1261" *)
  wire or_tmp_2960;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1278" *)
  wire or_tmp_3025;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1279" *)
  wire or_tmp_3032;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1029" *)
  wire or_tmp_306;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1325" *)
  wire or_tmp_3379;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1370" *)
  wire or_tmp_3487;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2595" *)
  wire or_tmp_3763;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2597" *)
  wire or_tmp_3768;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1031" *)
  wire or_tmp_378;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2606" *)
  wire or_tmp_3826;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2608" *)
  wire or_tmp_3832;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2611" *)
  wire or_tmp_3840;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2613" *)
  wire or_tmp_3849;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1034" *)
  wire or_tmp_389;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3537" *)
  wire or_tmp_4080;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3540" *)
  wire or_tmp_4081;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3543" *)
  wire or_tmp_4082;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3546" *)
  wire or_tmp_4084;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3550" *)
  wire or_tmp_4086;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3553" *)
  wire or_tmp_4087;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3558" *)
  wire or_tmp_4092;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3561" *)
  wire or_tmp_4095;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3564" *)
  wire or_tmp_4097;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3582" *)
  wire or_tmp_4102;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:1053" *)
  wire or_tmp_533;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2682" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2681" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2680" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2679" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2676" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2675" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2672" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2671" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2668" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2667" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2664" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2663" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2656" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2655" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2658" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2657" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2662" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2661" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2666" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2665" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2670" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2669" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2674" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2673" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2678" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2677" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2660" *)
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2659" *)
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2642" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2641" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2644" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2643" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2646" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2645" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2648" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2647" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2650" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2649" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2652" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2651" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2632" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2631" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2634" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2633" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2636" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2635" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2638" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2637" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2640" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2639" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2654" *)
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2653" *)
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2898" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2897" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2901" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2900" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2904" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2903" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2907" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2906" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2910" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2909" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2913" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2912" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2871" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2870" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2874" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2873" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2877" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2876" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2880" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2879" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2883" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2882" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2886" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2885" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2889" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2888" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2892" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2891" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2895" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2894" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2916" *)
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2915" *)
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2683" *)
  reg [4:0] reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2684" *)
  reg [9:0] reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3450" *)
  reg [1:0] reg_cfg_proc_precision_1_sva_st_40_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2686" *)
  reg [4:0] reg_chn_idata_data_sva_3_15_0_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2687" *)
  reg [9:0] reg_chn_idata_data_sva_3_15_0_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2685" *)
  reg reg_chn_idata_data_sva_3_15_0_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:2533" *)
  reg reg_chn_out_rsci_ld_core_psct_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3508" *)
  wire reg_cvt_else_cvt_else_nor_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:3524" *)
  reg reg_cvt_else_nor_dfs_9_cse;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0 = _03847_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10137" *) 1'b1;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl = { 1'b1, _04190_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10141" *) 7'b1110001;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl = chn_in_rsci_d_mxwt[30:24] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10145" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0 = _03848_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10149" *) 1'b1;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = { 1'b1, _04191_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10153" *) 7'b1110001;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = chn_in_rsci_d_mxwt[62:56] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10157" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0 = _03849_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10161" *) 1'b1;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = { 1'b1, _04192_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10165" *) 7'b1110001;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = chn_in_rsci_d_mxwt[94:88] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10169" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0 = _03850_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10173" *) 1'b1;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = { 1'b1, _04193_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10177" *) 7'b1110001;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = chn_in_rsci_d_mxwt[126:120] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10181" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0 = _03851_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10185" *) 1'b1;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = { 1'b1, _04194_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10189" *) 7'b1110001;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = chn_in_rsci_d_mxwt[158:152] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10193" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0 = _03852_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10197" *) 1'b1;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = { 1'b1, _04195_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10201" *) 7'b1110001;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = chn_in_rsci_d_mxwt[190:184] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10205" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0 = _03853_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10209" *) 1'b1;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = { 1'b1, _04196_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10213" *) 7'b1110001;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = chn_in_rsci_d_mxwt[222:216] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10217" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0 = _03854_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10221" *) 1'b1;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = { 1'b1, _04197_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10225" *) 7'b1110001;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = chn_in_rsci_d_mxwt[254:248] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10229" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0 = _03855_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10233" *) 1'b1;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = { 1'b1, _04198_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10237" *) 7'b1110001;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = chn_in_rsci_d_mxwt[286:280] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10241" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0 = _03856_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10245" *) 1'b1;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = { 1'b1, _04199_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10249" *) 7'b1110001;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = chn_in_rsci_d_mxwt[318:312] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10253" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0 = _03857_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10257" *) 1'b1;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = { 1'b1, _04200_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10261" *) 7'b1110001;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = chn_in_rsci_d_mxwt[350:344] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10265" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0 = _03858_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10269" *) 1'b1;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = { 1'b1, _04201_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10273" *) 7'b1110001;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = chn_in_rsci_d_mxwt[382:376] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10277" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0 = _03859_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10281" *) 1'b1;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = { 1'b1, _04202_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10285" *) 7'b1110001;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = chn_in_rsci_d_mxwt[414:408] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10289" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0 = _03860_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10293" *) 1'b1;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = { 1'b1, _04203_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10297" *) 7'b1110001;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = chn_in_rsci_d_mxwt[446:440] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10301" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0 = _03861_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10305" *) 1'b1;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = { 1'b1, _04204_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10309" *) 7'b1110001;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = chn_in_rsci_d_mxwt[478:472] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10313" *) 8'b11001101;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0 = _03862_[2:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10317" *) 1'b1;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl = { 1'b1, _04205_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10321" *) 7'b1110001;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl = chn_in_rsci_d_mxwt[510:504] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10325" *) 8'b11001101;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl = chn_in_rsci_d_mxwt[510:503] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10329" *) 9'b101110001;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = chn_in_rsci_d_mxwt[478:471] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10333" *) 9'b101110001;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = chn_in_rsci_d_mxwt[446:439] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10337" *) 9'b101110001;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = chn_in_rsci_d_mxwt[414:407] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10341" *) 9'b101110001;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = chn_in_rsci_d_mxwt[382:375] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10345" *) 9'b101110001;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = chn_in_rsci_d_mxwt[350:343] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10349" *) 9'b101110001;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = chn_in_rsci_d_mxwt[318:311] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10353" *) 9'b101110001;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = chn_in_rsci_d_mxwt[286:279] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10357" *) 9'b101110001;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = chn_in_rsci_d_mxwt[254:247] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10361" *) 9'b101110001;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = chn_in_rsci_d_mxwt[222:215] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10365" *) 9'b101110001;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = chn_in_rsci_d_mxwt[190:183] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10369" *) 9'b101110001;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = chn_in_rsci_d_mxwt[158:151] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10373" *) 9'b101110001;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = chn_in_rsci_d_mxwt[126:119] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10377" *) 9'b101110001;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = chn_in_rsci_d_mxwt[94:87] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10381" *) 9'b101110001;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = chn_in_rsci_d_mxwt[62:55] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10385" *) 9'b101110001;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl = chn_in_rsci_d_mxwt[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10389" *) 9'b101110001;
  assign cvt_1_FpMantRNE_24U_11U_else_acc_nl = chn_idata_data_sva_1_27_0_1[22:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10393" *) FpMantRNE_24U_11U_else_carry_1_sva_2;
  assign cvt_2_FpMantRNE_24U_11U_else_acc_1_nl = chn_idata_data_sva_1_59_31_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10419" *) FpMantRNE_24U_11U_else_carry_2_sva_2;
  assign cvt_3_FpMantRNE_24U_11U_else_acc_1_nl = chn_idata_data_sva_1_91_63_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10445" *) FpMantRNE_24U_11U_else_carry_3_sva_2;
  assign cvt_4_FpMantRNE_24U_11U_else_acc_2_nl = chn_idata_data_sva_1_123_95_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10471" *) FpMantRNE_24U_11U_else_carry_4_sva_2;
  assign cvt_5_FpMantRNE_24U_11U_else_acc_1_nl = chn_idata_data_sva_1_155_127_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10497" *) FpMantRNE_24U_11U_else_carry_5_sva_2;
  assign cvt_6_FpMantRNE_24U_11U_else_acc_2_nl = chn_idata_data_sva_1_187_159_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10523" *) FpMantRNE_24U_11U_else_carry_6_sva_2;
  assign cvt_7_FpMantRNE_24U_11U_else_acc_2_nl = chn_idata_data_sva_1_219_191_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10549" *) FpMantRNE_24U_11U_else_carry_7_sva_2;
  assign cvt_8_FpMantRNE_24U_11U_else_acc_3_nl = chn_idata_data_sva_1_251_223_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10575" *) FpMantRNE_24U_11U_else_carry_8_sva_2;
  assign cvt_9_FpMantRNE_24U_11U_else_acc_1_nl = chn_idata_data_sva_1_283_255_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10601" *) FpMantRNE_24U_11U_else_carry_9_sva_2;
  assign cvt_10_FpMantRNE_24U_11U_else_acc_2_nl = chn_idata_data_sva_1_315_287_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10627" *) FpMantRNE_24U_11U_else_carry_10_sva_2;
  assign cvt_11_FpMantRNE_24U_11U_else_acc_2_nl = chn_idata_data_sva_1_347_319_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10653" *) FpMantRNE_24U_11U_else_carry_11_sva_2;
  assign cvt_12_FpMantRNE_24U_11U_else_acc_3_nl = chn_idata_data_sva_1_379_351_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10679" *) FpMantRNE_24U_11U_else_carry_12_sva_2;
  assign cvt_13_FpMantRNE_24U_11U_else_acc_2_nl = chn_idata_data_sva_1_411_383_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10705" *) FpMantRNE_24U_11U_else_carry_13_sva_2;
  assign cvt_14_FpMantRNE_24U_11U_else_acc_3_nl = chn_idata_data_sva_1_443_415_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10731" *) FpMantRNE_24U_11U_else_carry_14_sva_2;
  assign cvt_15_FpMantRNE_24U_11U_else_acc_3_nl = chn_idata_data_sva_1_475_447_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10757" *) FpMantRNE_24U_11U_else_carry_15_sva_2;
  assign cvt_16_FpMantRNE_24U_11U_else_acc_4_nl = chn_idata_data_sva_1_507_479_1[23:14] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10783" *) FpMantRNE_24U_11U_else_carry_sva_2;
  assign cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl = { 1'b1, cvt_1_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_nl, _04240_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11011" *) 1'b1;
  assign cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl = { 1'b1, cvt_2_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl, _04243_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11021" *) 1'b1;
  assign cvt_3_IntSaturation_17U_8U_if_acc_1_nl = { _00171_[10], _00171_[10], _00171_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11028" *) 1'b1;
  assign cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl = { 1'b1, cvt_3_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl, _04246_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11035" *) 1'b1;
  assign cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl = { 1'b1, cvt_4_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl, _04249_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11044" *) 1'b1;
  assign cvt_5_IntSaturation_17U_8U_if_acc_1_nl = { _00172_[10], _00172_[10], _00172_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11050" *) 1'b1;
  assign cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl = { 1'b1, cvt_5_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl, _04252_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11057" *) 1'b1;
  assign cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl = { 1'b1, cvt_16_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_4_nl, _04255_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11066" *) 1'b1;
  assign cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl = { 1'b1, cvt_6_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl, _04258_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11075" *) 1'b1;
  assign cvt_1_IntSaturation_17U_8U_if_acc_nl = { _00173_[10], _00173_[10], _00173_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11081" *) 1'b1;
  assign cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl = { 1'b1, cvt_15_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl, _04261_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11088" *) 1'b1;
  assign cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl = { 1'b1, cvt_7_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl, _04264_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11098" *) 1'b1;
  assign cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl = { 1'b1, cvt_14_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl, _04267_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11107" *) 1'b1;
  assign cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl = { 1'b1, cvt_8_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl, _04270_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11116" *) 1'b1;
  assign cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl = { 1'b1, cvt_13_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl, _04273_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11125" *) 1'b1;
  assign cvt_9_IntSaturation_17U_8U_if_acc_1_nl = { _00174_[10], _00174_[10], _00174_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11131" *) 1'b1;
  assign cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl = { 1'b1, cvt_9_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl, _04276_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11138" *) 1'b1;
  assign cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl = { 1'b1, cvt_12_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl, _04279_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11147" *) 1'b1;
  assign cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl = { 1'b1, cvt_10_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl, _04282_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11156" *) 1'b1;
  assign cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl = { 1'b1, cvt_11_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl, _04285_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11165" *) 1'b1;
  assign cvt_4_FpMantRNE_17U_11U_else_acc_2_nl = cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11250" *) FpMantRNE_17U_11U_else_carry_4_sva;
  assign cvt_5_FpMantRNE_17U_11U_else_acc_1_nl = cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11264" *) FpMantRNE_17U_11U_else_carry_5_sva;
  assign cvt_6_FpMantRNE_17U_11U_else_acc_2_nl = cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11270" *) FpMantRNE_17U_11U_else_carry_6_sva;
  assign cvt_7_FpMantRNE_17U_11U_else_acc_2_nl = cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11284" *) FpMantRNE_17U_11U_else_carry_7_sva;
  assign cvt_8_FpMantRNE_17U_11U_else_acc_3_nl = cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11298" *) FpMantRNE_17U_11U_else_carry_8_sva;
  assign cvt_10_FpMantRNE_17U_11U_else_acc_2_nl = cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11312" *) FpMantRNE_17U_11U_else_carry_10_sva;
  assign cvt_11_FpMantRNE_17U_11U_else_acc_2_nl = cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11326" *) FpMantRNE_17U_11U_else_carry_11_sva;
  assign cvt_12_FpMantRNE_17U_11U_else_acc_3_nl = cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11340" *) FpMantRNE_17U_11U_else_carry_12_sva;
  assign cvt_13_FpMantRNE_17U_11U_else_acc_2_nl = cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11354" *) FpMantRNE_17U_11U_else_carry_13_sva;
  assign cvt_14_FpMantRNE_17U_11U_else_acc_3_nl = cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11368" *) FpMantRNE_17U_11U_else_carry_14_sva;
  assign cvt_15_FpMantRNE_17U_11U_else_acc_3_nl = cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11382" *) FpMantRNE_17U_11U_else_carry_15_sva;
  assign cvt_16_FpMantRNE_17U_11U_else_acc_4_nl = cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11396" *) FpMantRNE_17U_11U_else_carry_sva;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp = { _04310_, chn_in_rsci_d_mxwt[506:503] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11526" *) 1'b1;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = { _04312_, chn_in_rsci_d_mxwt[474:471] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11533" *) 1'b1;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = { _04314_, chn_in_rsci_d_mxwt[442:439] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11540" *) 1'b1;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = { _04316_, chn_in_rsci_d_mxwt[410:407] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11547" *) 1'b1;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = { _04318_, chn_in_rsci_d_mxwt[378:375] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11554" *) 1'b1;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = { _04320_, chn_in_rsci_d_mxwt[346:343] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11561" *) 1'b1;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = { _04322_, chn_in_rsci_d_mxwt[314:311] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11568" *) 1'b1;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = { _04324_, chn_in_rsci_d_mxwt[282:279] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11575" *) 1'b1;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = { _04326_, chn_in_rsci_d_mxwt[250:247] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11582" *) 1'b1;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = { _04328_, chn_in_rsci_d_mxwt[218:215] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11589" *) 1'b1;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = { _04330_, chn_in_rsci_d_mxwt[186:183] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11596" *) 1'b1;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = { _04331_, chn_in_rsci_d_mxwt[154:151] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11601" *) 1'b1;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = { _04333_, chn_in_rsci_d_mxwt[122:119] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11610" *) 1'b1;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = { _04335_, chn_in_rsci_d_mxwt[90:87] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11617" *) 1'b1;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = { _04337_, chn_in_rsci_d_mxwt[58:55] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11624" *) 1'b1;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp = { _04339_, chn_in_rsci_d_mxwt[26:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11631" *) 1'b1;
  assign cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_2_sva_2, IntShiftRightSat_49U_6U_17U_o_16_2_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2, IntShiftRightSat_49U_6U_17U_o_0_2_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11756" *) 1'b1;
  assign cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_4_sva_2, IntShiftRightSat_49U_6U_17U_o_16_4_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2, IntShiftRightSat_49U_6U_17U_o_0_4_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11762" *) 1'b1;
  assign cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_3_sva_3, IntShiftRightSat_49U_6U_17U_o_16_3_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2, IntShiftRightSat_49U_6U_17U_o_0_3_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11768" *) 1'b1;
  assign cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_6_sva_2, IntShiftRightSat_49U_6U_17U_o_16_6_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2, IntShiftRightSat_49U_6U_17U_o_0_6_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11774" *) 1'b1;
  assign cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_8_sva_2, IntShiftRightSat_49U_6U_17U_o_16_8_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2, IntShiftRightSat_49U_6U_17U_o_0_8_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11780" *) 1'b1;
  assign cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_7_sva_2, IntShiftRightSat_49U_6U_17U_o_16_7_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2, IntShiftRightSat_49U_6U_17U_o_0_7_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11786" *) 1'b1;
  assign cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_5_sva_3, IntShiftRightSat_49U_6U_17U_o_16_5_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2, IntShiftRightSat_49U_6U_17U_o_0_5_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11792" *) 1'b1;
  assign cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_10_sva_2, IntShiftRightSat_49U_6U_17U_o_16_10_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2, IntShiftRightSat_49U_6U_17U_o_0_10_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11798" *) 1'b1;
  assign cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_12_sva_2, IntShiftRightSat_49U_6U_17U_o_16_12_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2, IntShiftRightSat_49U_6U_17U_o_0_12_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11807" *) 1'b1;
  assign cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_11_sva_2, IntShiftRightSat_49U_6U_17U_o_16_11_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2, IntShiftRightSat_49U_6U_17U_o_0_11_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11813" *) 1'b1;
  assign { _03864_[17:9], cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl } = { IntShiftRightSat_49U_6U_17U_o_16_14_sva_2, IntShiftRightSat_49U_6U_17U_o_16_14_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2, IntShiftRightSat_49U_6U_17U_o_0_14_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11822" *) 1'b1;
  assign cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl = { IntShiftRightSat_49U_6U_17U_o_16_sva_2, IntShiftRightSat_49U_6U_17U_o_16_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_sva_2, IntShiftRightSat_49U_6U_17U_o_0_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11828" *) 1'b1;
  assign cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_15_sva_2, IntShiftRightSat_49U_6U_17U_o_16_15_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2, IntShiftRightSat_49U_6U_17U_o_0_15_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11834" *) 1'b1;
  assign cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_13_sva_2, IntShiftRightSat_49U_6U_17U_o_16_13_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2, IntShiftRightSat_49U_6U_17U_o_0_13_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11840" *) 1'b1;
  assign cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_9_sva_3, IntShiftRightSat_49U_6U_17U_o_16_9_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2, IntShiftRightSat_49U_6U_17U_o_0_9_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11846" *) 1'b1;
  assign cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl = { IntShiftRightSat_49U_6U_17U_o_16_1_sva_3, IntShiftRightSat_49U_6U_17U_o_16_1_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2, IntShiftRightSat_49U_6U_17U_o_0_1_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11852" *) 1'b1;
  assign cvt_1_IntSaturation_17U_16U_if_acc_nl = { _00187_[2], _00187_[2], _00187_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11889" *) 1'b1;
  assign cvt_2_IntSaturation_17U_16U_if_acc_1_nl = { _00188_[2], _00188_[2], _00188_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11893" *) 1'b1;
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11930" *) cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  assign cvt_3_IntSaturation_17U_16U_if_acc_1_nl = { _00189_[2], _00189_[2], _00189_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11937" *) 1'b1;
  assign cvt_4_IntSaturation_17U_16U_if_acc_2_nl = { or_dcpl_109, or_dcpl_109, _00190_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11941" *) 1'b1;
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11978" *) cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12018" *) cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  assign cvt_5_IntSaturation_17U_16U_if_acc_1_nl = { or_dcpl_111, or_dcpl_111, _00191_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12025" *) 1'b1;
  assign cvt_6_IntSaturation_17U_16U_if_acc_2_nl = { or_dcpl_114, or_dcpl_114, _00192_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12029" *) 1'b1;
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12066" *) cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  assign cvt_7_IntSaturation_17U_16U_if_acc_2_nl = { or_dcpl_116, or_dcpl_116, _00193_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12073" *) 1'b1;
  assign cvt_8_IntSaturation_17U_16U_if_acc_3_nl = { or_dcpl_120, or_dcpl_120, _00194_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12077" *) 1'b1;
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12114" *) cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12154" *) cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12194" *) cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  assign cvt_9_IntSaturation_17U_16U_if_acc_1_nl = { _00195_[2], _00195_[2], _00195_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12201" *) 1'b1;
  assign cvt_10_IntSaturation_17U_16U_if_acc_2_nl = { or_dcpl_125, or_dcpl_125, _00196_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12205" *) 1'b1;
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12242" *) cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  assign cvt_11_IntSaturation_17U_16U_if_acc_2_nl = { or_dcpl_127, or_dcpl_127, _00197_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12249" *) 1'b1;
  assign cvt_12_IntSaturation_17U_16U_if_acc_3_nl = { or_dcpl_131, or_dcpl_131, _00198_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12253" *) 1'b1;
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12290" *) cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12330" *) cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  assign cvt_13_IntSaturation_17U_16U_if_acc_2_nl = { or_dcpl_133, or_dcpl_133, _00199_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12337" *) 1'b1;
  assign cvt_14_IntSaturation_17U_16U_if_acc_3_nl = { or_dcpl_137, or_dcpl_137, _00200_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12341" *) 1'b1;
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12378" *) cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  assign cvt_15_IntSaturation_17U_16U_if_acc_3_nl = { or_dcpl_140, or_dcpl_140, _00201_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12385" *) 1'b1;
  assign cvt_16_IntSaturation_17U_16U_if_acc_4_nl = { or_dcpl_144, or_dcpl_144, _00202_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12389" *) 1'b1;
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12426" *) cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_8_nl;
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12466" *) cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12506" *) cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12546" *) cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp = { IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[111], IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[111:63] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12586" *) cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12610" *) cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12638" *) cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12666" *) cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12694" *) cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12722" *) cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12750" *) cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12778" *) cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12806" *) cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12834" *) cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12862" *) cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12890" *) cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12918" *) cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12946" *) cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12974" *) cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13002" *) cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva = { IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[74], IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[74:31] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13030" *) cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_8_nl;
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl = { 1'b1, _04485_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13042" *) 1'b1;
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = { 1'b1, _04486_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13051" *) 1'b1;
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = { 1'b1, _04487_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13060" *) 1'b1;
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = { 1'b1, _04488_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13069" *) 1'b1;
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = { 1'b1, _04489_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13078" *) 1'b1;
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = { 1'b1, _04490_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13087" *) 1'b1;
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = { 1'b1, _04491_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13096" *) 1'b1;
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = { 1'b1, _04492_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13105" *) 1'b1;
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = { 1'b1, _04493_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13114" *) 1'b1;
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = { 1'b1, _04494_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13123" *) 1'b1;
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = { 1'b1, _04495_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13132" *) 1'b1;
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = { 1'b1, _04496_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13141" *) 1'b1;
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = { 1'b1, _04497_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13150" *) 1'b1;
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = { 1'b1, _04498_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13159" *) 1'b1;
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = { 1'b1, _04499_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13168" *) 1'b1;
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl = { 1'b1, _04500_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13177" *) 1'b1;
  assign cvt_1_IntSaturation_17U_8U_else_if_acc_nl = { IntShiftRightSat_49U_6U_17U_o_16_1_sva_4, IntShiftRightSat_49U_6U_17U_o_16_1_sva_4, reg_chn_idata_data_sva_3_15_0_1_reg, reg_chn_idata_data_sva_3_15_0_2_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13189" *) 1'b1;
  assign cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_2_sva_3, IntShiftRightSat_49U_6U_17U_o_16_2_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13203" *) 1'b1;
  assign cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_3_sva_4, IntShiftRightSat_49U_6U_17U_o_16_3_sva_4, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13221" *) 1'b1;
  assign cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_4_sva_3, IntShiftRightSat_49U_6U_17U_o_16_4_sva_3, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[14:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13234" *) 1'b1;
  assign cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_5_sva_4, IntShiftRightSat_49U_6U_17U_o_16_5_sva_4, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13248" *) 1'b1;
  assign cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_6_sva_3, IntShiftRightSat_49U_6U_17U_o_16_6_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13262" *) 1'b1;
  assign cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_7_sva_3, IntShiftRightSat_49U_6U_17U_o_16_7_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13276" *) 1'b1;
  assign cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_8_sva_3, IntShiftRightSat_49U_6U_17U_o_16_8_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13290" *) 1'b1;
  assign cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_9_sva_4, IntShiftRightSat_49U_6U_17U_o_16_9_sva_4, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13304" *) 1'b1;
  assign cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_10_sva_3, IntShiftRightSat_49U_6U_17U_o_16_10_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13318" *) 1'b1;
  assign cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_11_sva_3, IntShiftRightSat_49U_6U_17U_o_16_11_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13332" *) 1'b1;
  assign cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_12_sva_3, IntShiftRightSat_49U_6U_17U_o_16_12_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13346" *) 1'b1;
  assign cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_13_sva_3, IntShiftRightSat_49U_6U_17U_o_16_13_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13360" *) 1'b1;
  assign cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_15_sva_3, IntShiftRightSat_49U_6U_17U_o_16_15_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13383" *) 1'b1;
  assign cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl = { IntShiftRightSat_49U_6U_17U_o_16_sva_3, IntShiftRightSat_49U_6U_17U_o_16_sva_3, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg, reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13397" *) 1'b1;
  assign cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_14_sva_3, IntShiftRightSat_49U_6U_17U_o_16_14_sva_3, reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg, reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg[9:6] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13409" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva = { _04518_, _04519_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13417" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva = { _04520_, _04521_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13422" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva = { _04522_, _04523_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13427" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva = { _04524_, _04525_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13432" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva = { _04526_, _04527_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13437" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva = { _04528_, _04529_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13442" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva = { _04530_, _04531_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13447" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva = { _04532_, _04533_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13452" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva = { _04534_, _04535_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13457" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva = { _04536_, _04537_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13462" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva = { _04538_, _04539_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13467" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva = { _04540_, _04541_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13472" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva = { _04542_, _04543_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13477" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva = { _04544_, _04545_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13482" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva = { _04546_, _04547_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13487" *) 1'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva = { _04548_, _04549_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13492" *) 1'b1;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva = cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13532" *) cvt_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl;
  assign cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13537" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva = cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13548" *) cvt_2_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  assign cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13553" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva = cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13564" *) cvt_3_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  assign cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13569" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva = cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13580" *) cvt_4_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  assign cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13585" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva = cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13596" *) cvt_5_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  assign cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13601" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva = cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13612" *) cvt_6_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  assign cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13617" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva = cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13628" *) cvt_7_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  assign cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13633" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva = cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13644" *) cvt_8_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  assign cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13649" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva = cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13660" *) cvt_9_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  assign cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13665" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva = cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13676" *) cvt_10_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  assign cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13681" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva = cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13692" *) cvt_11_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  assign cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13697" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva = cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13708" *) cvt_12_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  assign cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13713" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva = cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13724" *) cvt_13_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  assign cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13729" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva = cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13740" *) cvt_14_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  assign cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13745" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva = cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13756" *) cvt_15_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  assign cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13761" *) 23'b11111111111111111111111;
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva = cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_itm[23:13] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13772" *) cvt_16_FpMantDecShiftRight_23U_8U_10U_carry_and_4_nl;
  assign cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl = FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13777" *) 23'b11111111111111111111111;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva = _00203_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13913" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva = _00204_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13917" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva = _00205_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13921" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva = _00206_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13925" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva = _00207_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13929" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva = _00208_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13933" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva = _00209_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13937" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva = _00210_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13941" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva = _00211_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13945" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva = _00212_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13949" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva = _00213_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13953" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva = _00214_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13957" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva = _00215_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13961" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva = _00216_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13965" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva = _00217_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13969" *) 1'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva = _00218_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13973" *) 1'b1;
  assign cvt_1_IntSaturation_17U_16U_else_if_acc_nl = { IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14008" *) 1'b1;
  assign cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14012" *) 1'b1;
  assign cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14016" *) 1'b1;
  assign cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14020" *) 1'b1;
  assign cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14024" *) 1'b1;
  assign cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14028" *) 1'b1;
  assign cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14032" *) 1'b1;
  assign cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14036" *) 1'b1;
  assign cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14040" *) 1'b1;
  assign cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14044" *) 1'b1;
  assign cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14048" *) 1'b1;
  assign cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14052" *) 1'b1;
  assign cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14056" *) 1'b1;
  assign cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14060" *) 1'b1;
  assign cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl = { IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14064" *) 1'b1;
  assign cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0[14] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14068" *) 1'b1;
  assign nl_cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2 = _00219_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22484" *) 5'b11101;
  assign nl_cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 = _00220_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22490" *) 5'b11101;
  assign nl_cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 = _00221_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22493" *) 5'b11101;
  assign nl_cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = _00222_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22496" *) 5'b11101;
  assign nl_cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0] = _00223_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22499" *) 5'b11101;
  assign nl_cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0] = _00224_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22503" *) 5'b11101;
  assign nl_cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0] = _00225_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22506" *) 5'b11101;
  assign nl_cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2[4:0] = _00226_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22509" *) 5'b11101;
  assign nl_cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = _00227_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22512" *) 5'b11101;
  assign nl_cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = _00228_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22515" *) 5'b11101;
  assign nl_cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = _00229_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22518" *) 5'b11101;
  assign nl_cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 = _00230_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22521" *) 5'b11101;
  assign nl_cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0] = _00231_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22524" *) 5'b11101;
  assign nl_cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 = _00232_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22527" *) 5'b11101;
  assign nl_cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 = _00233_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22530" *) 5'b11101;
  assign nl_cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2 = _00234_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22535" *) 5'b11101;
  assign cvt_10_IntSaturation_17U_8U_if_acc_2_nl = { _00175_[10], _00175_[10], _00175_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22847" *) 1'b1;
  assign cvt_2_IntSaturation_17U_8U_if_acc_1_nl = { _00176_[10], _00176_[10], _00176_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22850" *) 1'b1;
  assign cvt_4_IntSaturation_17U_8U_if_acc_2_nl = { _00177_[10], _00177_[10], _00177_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22853" *) 1'b1;
  assign cvt_6_IntSaturation_17U_8U_if_acc_2_nl = { _00178_[10], _00178_[10], _00178_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22856" *) 1'b1;
  assign cvt_7_IntSaturation_17U_8U_if_acc_2_nl = { _00179_[10], _00179_[10], _00179_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22859" *) 1'b1;
  assign cvt_16_IntSaturation_17U_8U_if_acc_4_nl = { _00180_[10], _00180_[10], _00180_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22862" *) 1'b1;
  assign cvt_8_IntSaturation_17U_8U_if_acc_3_nl = { _00181_[10], _00181_[10], _00181_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22865" *) 1'b1;
  assign cvt_15_IntSaturation_17U_8U_if_acc_3_nl = { _00182_[10], _00182_[10], _00182_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22868" *) 1'b1;
  assign cvt_13_IntSaturation_17U_8U_if_acc_2_nl = { _00183_[10], _00183_[10], _00183_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22871" *) 1'b1;
  assign cvt_11_IntSaturation_17U_8U_if_acc_2_nl = { _00184_[10], _00184_[10], _00184_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22874" *) 1'b1;
  assign cvt_12_IntSaturation_17U_8U_if_acc_3_nl = { _00185_[10], _00185_[10], _00185_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22877" *) 1'b1;
  assign cvt_3_FpMantRNE_17U_11U_else_acc_1_nl = cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22942" *) FpMantRNE_17U_11U_else_carry_3_sva;
  assign cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl = { IntShiftRightSat_49U_6U_17U_o_16_sva_2, IntShiftRightSat_49U_6U_17U_o_16_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_sva_2, IntShiftRightSat_49U_6U_17U_o_0_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23206" *) 18'b111111111111111111;
  assign cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_15_sva_2, IntShiftRightSat_49U_6U_17U_o_16_15_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2, IntShiftRightSat_49U_6U_17U_o_0_15_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23212" *) 18'b111111111111111111;
  assign cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_14_sva_2, IntShiftRightSat_49U_6U_17U_o_16_14_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2, IntShiftRightSat_49U_6U_17U_o_0_14_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23218" *) 18'b111111111111111111;
  assign cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_13_sva_2, IntShiftRightSat_49U_6U_17U_o_16_13_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2, IntShiftRightSat_49U_6U_17U_o_0_13_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23224" *) 18'b111111111111111111;
  assign cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_12_sva_2, IntShiftRightSat_49U_6U_17U_o_16_12_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2, IntShiftRightSat_49U_6U_17U_o_0_12_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23230" *) 18'b111111111111111111;
  assign cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_11_sva_2, IntShiftRightSat_49U_6U_17U_o_16_11_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2, IntShiftRightSat_49U_6U_17U_o_0_11_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23236" *) 18'b111111111111111111;
  assign cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_10_sva_2, IntShiftRightSat_49U_6U_17U_o_16_10_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2, IntShiftRightSat_49U_6U_17U_o_0_10_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23242" *) 18'b111111111111111111;
  assign cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_9_sva_3, IntShiftRightSat_49U_6U_17U_o_16_9_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2, IntShiftRightSat_49U_6U_17U_o_0_9_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23248" *) 18'b111111111111111111;
  assign cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = { IntShiftRightSat_49U_6U_17U_o_16_8_sva_2, IntShiftRightSat_49U_6U_17U_o_16_8_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2, IntShiftRightSat_49U_6U_17U_o_0_8_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23254" *) 18'b111111111111111111;
  assign cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_7_sva_2, IntShiftRightSat_49U_6U_17U_o_16_7_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2, IntShiftRightSat_49U_6U_17U_o_0_7_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23260" *) 18'b111111111111111111;
  assign cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_6_sva_2, IntShiftRightSat_49U_6U_17U_o_16_6_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2, IntShiftRightSat_49U_6U_17U_o_0_6_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23266" *) 18'b111111111111111111;
  assign cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_5_sva_3, IntShiftRightSat_49U_6U_17U_o_16_5_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2, IntShiftRightSat_49U_6U_17U_o_0_5_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23272" *) 18'b111111111111111111;
  assign cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = { IntShiftRightSat_49U_6U_17U_o_16_4_sva_2, IntShiftRightSat_49U_6U_17U_o_16_4_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2, IntShiftRightSat_49U_6U_17U_o_0_4_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23278" *) 18'b111111111111111111;
  assign cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_3_sva_3, IntShiftRightSat_49U_6U_17U_o_16_3_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2, IntShiftRightSat_49U_6U_17U_o_0_3_sva_3 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23284" *) 18'b111111111111111111;
  assign cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = { IntShiftRightSat_49U_6U_17U_o_16_2_sva_2, IntShiftRightSat_49U_6U_17U_o_16_2_sva_2, IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2, IntShiftRightSat_49U_6U_17U_o_0_2_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23290" *) 18'b111111111111111111;
  assign cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl = { IntShiftRightSat_49U_6U_17U_o_16_1_sva_3, IntShiftRightSat_49U_6U_17U_o_16_1_sva_3, IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2, IntShiftRightSat_49U_6U_17U_o_0_1_sva_2 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23296" *) 18'b111111111111111111;
  assign cvt_14_IntSaturation_17U_8U_if_acc_3_nl = { _00186_[10], _00186_[10], _00186_[8:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23312" *) 1'b1;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0, _00235_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23633" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0, _00236_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23656" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0, _00237_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23679" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0, _00238_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23702" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0, _00239_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23725" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0, _00240_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23748" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0, _00241_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23771" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2[4:0] = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0, _00242_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23794" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2[4:0] = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0, _00243_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23817" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0, _00244_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23840" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0, _00245_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23863" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0, _00246_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23886" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0, _00247_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23909" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0, _00248_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23932" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0, _00249_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23955" *) 4'b1101;
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 = { FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0, _00250_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23978" *) 4'b1101;
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7125" *) 5'b11111;
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7134" *) 5'b11111;
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7143" *) 5'b11111;
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7152" *) 5'b11111;
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7161" *) 5'b11111;
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7170" *) 5'b11111;
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7179" *) 5'b11111;
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7188" *) 5'b11111;
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7197" *) 5'b11111;
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7206" *) 5'b11111;
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7215" *) 5'b11111;
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7224" *) 5'b11111;
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7233" *) 5'b11111;
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7242" *) 5'b11111;
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7251" *) 5'b11111;
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg_s[4:0] = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7260" *) 5'b11111;
  assign cvt_2_FpMantRNE_17U_11U_else_acc_1_nl = FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9113" *) FpMantRNE_17U_11U_else_carry_2_sva;
  assign cvt_9_FpMantRNE_17U_11U_else_acc_1_nl = FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9416" *) FpMantRNE_17U_11U_else_carry_9_sva;
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl = _00001_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9509" *) 1'b1;
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = _00003_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9530" *) 1'b1;
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = _00004_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9551" *) 1'b1;
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = _00005_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9578" *) 1'b1;
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = _00006_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9592" *) 1'b1;
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = _00007_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9611" *) 1'b1;
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = _00008_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9624" *) 1'b1;
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = _00009_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9637" *) 1'b1;
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = _00010_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9653" *) 1'b1;
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = _00011_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9669" *) 1'b1;
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = _00012_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9685" *) 1'b1;
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = _00013_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9701" *) 1'b1;
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = _00014_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9718" *) 1'b1;
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = _00015_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9732" *) 1'b1;
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = _00016_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9752" *) 1'b1;
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl = _00017_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9766" *) 1'b1;
  assign cvt_1_FpMantRNE_17U_11U_else_acc_nl = FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[15:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9799" *) FpMantRNE_17U_11U_else_carry_1_sva;
  assign IntSaturation_17U_16U_o_and_21_rgt = cvt_11_IntSaturation_17U_16U_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10000" *) _04174_;
  assign _01433_ = cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10004" *) _04175_;
  assign IntSaturation_17U_16U_and_19_rgt = _01433_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10004" *) _04174_;
  assign IntSaturation_17U_16U_o_and_19_rgt = cvt_10_IntSaturation_17U_16U_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10006" *) _04174_;
  assign _01434_ = cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10010" *) _04176_;
  assign IntSaturation_17U_16U_and_17_rgt = _01434_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10010" *) _04174_;
  assign IntSaturation_17U_16U_o_and_17_rgt = cvt_9_IntSaturation_17U_16U_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10012" *) _04174_;
  assign _01435_ = cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10016" *) _04177_;
  assign IntSaturation_17U_16U_and_15_rgt = _01435_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10016" *) _04174_;
  assign IntSaturation_17U_16U_o_and_15_rgt = cvt_8_IntSaturation_17U_16U_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10018" *) _04174_;
  assign _01436_ = cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10022" *) _04178_;
  assign IntSaturation_17U_16U_and_13_rgt = _01436_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10022" *) _04174_;
  assign IntSaturation_17U_16U_o_and_13_rgt = cvt_7_IntSaturation_17U_16U_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10024" *) _04174_;
  assign _01437_ = cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10028" *) _04179_;
  assign IntSaturation_17U_16U_and_11_rgt = _01437_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10028" *) _04174_;
  assign IntSaturation_17U_16U_o_and_11_rgt = cvt_6_IntSaturation_17U_16U_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10030" *) _04174_;
  assign _01438_ = cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10034" *) _04180_;
  assign IntSaturation_17U_16U_and_9_rgt = _01438_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10034" *) _04174_;
  assign IntSaturation_17U_16U_o_and_9_rgt = cvt_5_IntSaturation_17U_16U_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10036" *) _04174_;
  assign _01439_ = cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10040" *) _04181_;
  assign IntSaturation_17U_16U_and_7_rgt = _01439_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10040" *) _04174_;
  assign IntSaturation_17U_16U_o_and_7_rgt = cvt_4_IntSaturation_17U_16U_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10042" *) _04174_;
  assign _01440_ = cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10046" *) _04182_;
  assign IntSaturation_17U_16U_and_5_rgt = _01440_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10046" *) _04174_;
  assign IntSaturation_17U_16U_o_and_5_rgt = cvt_3_IntSaturation_17U_16U_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10048" *) _04174_;
  assign _01441_ = cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10052" *) _04183_;
  assign IntSaturation_17U_16U_and_3_rgt = _01441_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10052" *) _04174_;
  assign IntSaturation_17U_16U_o_and_3_rgt = cvt_2_IntSaturation_17U_16U_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10054" *) _04174_;
  assign _01442_ = cvt_1_IntSaturation_17U_16U_else_if_acc_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10058" *) _04184_;
  assign IntSaturation_17U_16U_and_1_rgt = _01442_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10058" *) _04174_;
  assign IntSaturation_17U_16U_o_and_1_rgt = cvt_1_IntSaturation_17U_16U_if_acc_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10060" *) _04174_;
  assign IntSaturation_17U_16U_and_33_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10063" *) mux_1626_nl;
  assign and_1386_cse = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10068" *) and_tmp_12;
  assign and_1385_rgt = and_tmp_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10069" *) and_dcpl_114;
  assign _01443_ = or_dcpl_16 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10071" *) or_4862_cse;
  assign _01444_ = _01443_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10071" *) or_4714_cse;
  assign _01445_ = _01444_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10071" *) and_dcpl_401;
  assign _01446_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10075" *) IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse;
  assign IntShiftRightSat_49U_6U_17U_oelse_and_cse = _01446_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10075" *) mux_272_cse;
  assign _01447_ = _01444_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10079" *) or_400_cse_1;
  assign _01448_ = _01447_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10079" *) and_dcpl_401;
  assign _01449_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10084" *) IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse;
  assign IntShiftRightSat_49U_6U_17U_oelse_and_18_cse = _01449_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10084" *) mux_377_nl;
  assign _01450_ = or_dcpl_32 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *) or_4862_cse;
  assign _01451_ = _01450_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *) or_4714_cse;
  assign _01452_ = _01451_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *) or_400_cse_1;
  assign _01453_ = _01452_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10086" *) and_dcpl_401;
  assign IntShiftRightSat_49U_6U_17U_oelse_and_22_cse = _01449_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10089" *) mux_272_cse;
  assign _01454_ = _01444_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *) or_5189_cse;
  assign _01455_ = _01454_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *) and_dcpl_626;
  assign _01456_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *) _05428_;
  assign IntShiftRightSat_49U_6U_17U_oelse_and_25_cse = _01456_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10092" *) mux_320_cse;
  assign _01457_ = _01451_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10094" *) or_5189_cse;
  assign _01458_ = _01457_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10094" *) and_dcpl_626;
  assign and_1467_rgt = and_tmp_11 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10096" *) or_5189_cse;
  assign _01459_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10104" *) FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse;
  assign FpIntToFloat_17U_5U_10U_is_inf_and_28_cse = _01459_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10104" *) _04189_;
  assign _01460_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10110" *) FpIntToFloat_17U_5U_10U_if_nor_10_cse;
  assign FpIntToFloat_17U_5U_10U_if_and_31_cse = _01460_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10110" *) mux_119_nl;
  assign FpIntToFloat_17U_5U_10U_if_and_33_cse = _01460_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10114" *) mux_125_nl;
  assign FpIntToFloat_17U_5U_10U_if_and_36_cse = _01460_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10119" *) mux_134_cse;
  assign _01461_ = and_2186_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10125" *) or_5189_cse;
  assign and_550_cse = _01461_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10125" *) fsm_output[1];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl = _04206_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10403" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl = cvt_1_FpMantRNE_24U_11U_else_and_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10405" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl = _04207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10429" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl = cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10431" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl = _04208_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl = cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10457" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl = _04209_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10481" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl = cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10483" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl = _04210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10507" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl = cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10509" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl = _04211_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10533" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl = cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10535" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl = _04212_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10559" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl = cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10561" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl = _04213_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10585" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl = cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10587" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl = _04214_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10611" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl = cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl = _04215_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10637" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl = cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10639" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl = _04216_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10663" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl = cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10665" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl = _04217_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10689" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl = cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10691" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl = _04218_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10715" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl = cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10717" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl = _04219_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10741" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl = cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10743" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl = _04220_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10767" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl = cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10769" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl = _04221_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10793" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl = cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10795" *) FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c;
  assign _01462_ = IntShiftRightSat_49U_6U_17U_o_0_14_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11235" *) _04286_;
  assign _01463_ = _04287_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11261" *) FpMantRNE_17U_11U_else_mux_7_nl;
  assign _01464_ = _04288_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11261" *) FpIntToFloat_17U_5U_10U_else_mux_10_nl;
  assign _01465_ = _04289_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11281" *) FpMantRNE_17U_11U_else_mux_11_nl;
  assign _01466_ = _04290_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11281" *) FpIntToFloat_17U_5U_10U_else_mux_16_nl;
  assign _01467_ = _04291_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11295" *) FpMantRNE_17U_11U_else_mux_13_nl;
  assign _01468_ = _04292_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11295" *) FpIntToFloat_17U_5U_10U_else_mux_19_nl;
  assign _01469_ = _04293_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11309" *) FpMantRNE_17U_11U_else_mux_15_nl;
  assign _01470_ = _04294_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11309" *) FpIntToFloat_17U_5U_10U_else_mux_22_nl;
  assign _01471_ = _04295_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11323" *) FpMantRNE_17U_11U_else_mux_19_nl;
  assign _01472_ = _04296_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11323" *) FpIntToFloat_17U_5U_10U_else_mux_28_nl;
  assign _01473_ = _04297_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11337" *) FpMantRNE_17U_11U_else_mux_21_nl;
  assign _01474_ = _04298_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11337" *) FpIntToFloat_17U_5U_10U_else_mux_31_nl;
  assign _01475_ = _04299_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11351" *) FpMantRNE_17U_11U_else_mux_23_nl;
  assign _01476_ = _04300_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11351" *) FpIntToFloat_17U_5U_10U_else_mux_34_nl;
  assign _01477_ = _04301_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11365" *) FpMantRNE_17U_11U_else_mux_25_nl;
  assign _01478_ = _04302_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11365" *) FpIntToFloat_17U_5U_10U_else_mux_37_nl;
  assign _01479_ = _04303_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11379" *) FpMantRNE_17U_11U_else_mux_27_nl;
  assign _01480_ = _04304_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11379" *) FpIntToFloat_17U_5U_10U_else_mux_40_nl;
  assign _01481_ = _04305_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11393" *) FpMantRNE_17U_11U_else_mux_29_nl;
  assign _01482_ = _04306_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11393" *) FpIntToFloat_17U_5U_10U_else_mux_43_nl;
  assign _01483_ = _04307_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11407" *) FpMantRNE_17U_11U_else_mux_31_nl;
  assign _01484_ = _04308_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11407" *) FpIntToFloat_17U_5U_10U_else_mux_46_nl;
  assign FpMantRNE_24U_11U_else_carry_1_sva_mx0w0 = chn_in_rsci_d_mxwt[12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *) _05537_;
  assign FpMantRNE_24U_11U_else_carry_2_sva_mx0w0 = chn_in_rsci_d_mxwt[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *) _05549_;
  assign FpMantRNE_24U_11U_else_carry_3_sva_mx0w0 = chn_in_rsci_d_mxwt[76] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *) _05561_;
  assign FpMantRNE_24U_11U_else_carry_4_sva_mx0w0 = chn_in_rsci_d_mxwt[108] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *) _05573_;
  assign FpMantRNE_24U_11U_else_carry_5_sva_mx0w0 = chn_in_rsci_d_mxwt[140] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *) _05585_;
  assign FpMantRNE_24U_11U_else_carry_6_sva_mx0w0 = chn_in_rsci_d_mxwt[172] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *) _05597_;
  assign FpMantRNE_24U_11U_else_carry_7_sva_mx0w0 = chn_in_rsci_d_mxwt[204] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *) _05609_;
  assign FpMantRNE_24U_11U_else_carry_8_sva_mx0w0 = chn_in_rsci_d_mxwt[236] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *) _05621_;
  assign FpMantRNE_24U_11U_else_carry_9_sva_mx0w0 = chn_in_rsci_d_mxwt[268] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *) _05633_;
  assign FpMantRNE_24U_11U_else_carry_10_sva_mx0w0 = chn_in_rsci_d_mxwt[300] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11487" *) _05645_;
  assign FpMantRNE_24U_11U_else_carry_11_sva_mx0w0 = chn_in_rsci_d_mxwt[332] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11493" *) _05657_;
  assign FpMantRNE_24U_11U_else_carry_12_sva_mx0w0 = chn_in_rsci_d_mxwt[364] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11499" *) _05669_;
  assign FpMantRNE_24U_11U_else_carry_13_sva_mx0w0 = chn_in_rsci_d_mxwt[396] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11505" *) _05681_;
  assign FpMantRNE_24U_11U_else_carry_14_sva_mx0w0 = chn_in_rsci_d_mxwt[428] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11511" *) _05693_;
  assign FpMantRNE_24U_11U_else_carry_15_sva_mx0w0 = chn_in_rsci_d_mxwt[460] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11517" *) _05705_;
  assign FpMantRNE_24U_11U_else_carry_sva_mx0w0 = chn_in_rsci_d_mxwt[492] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *) _05717_;
  assign cvt_16_FpMantRNE_24U_11U_else_and_4_tmp = FpMantRNE_24U_11U_else_carry_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11529" *) _03866_;
  assign cvt_15_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_15_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11536" *) _03867_;
  assign cvt_14_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_14_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11543" *) _03868_;
  assign cvt_13_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_13_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11550" *) _03869_;
  assign cvt_12_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_12_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11557" *) _03870_;
  assign cvt_11_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_11_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11564" *) _03871_;
  assign cvt_10_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_10_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11571" *) _03872_;
  assign cvt_9_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_9_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11578" *) _03873_;
  assign cvt_8_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_8_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11585" *) _03874_;
  assign cvt_7_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_7_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11592" *) _03875_;
  assign cvt_6_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_6_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11599" *) _03876_;
  assign cvt_5_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_5_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11604" *) _03877_;
  assign cvt_4_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_4_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11613" *) _03879_;
  assign cvt_3_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11620" *) _03880_;
  assign cvt_2_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11627" *) _03881_;
  assign cvt_1_FpMantRNE_24U_11U_else_and_tmp = FpMantRNE_24U_11U_else_carry_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11634" *) _03882_;
  assign _01485_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_32_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11639" *) _04340_;
  assign _01486_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_33_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11645" *) _04343_;
  assign _01487_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_34_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11651" *) _04346_;
  assign _01488_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_35_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11657" *) _04349_;
  assign _01489_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_36_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11663" *) _04352_;
  assign _01490_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_37_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11669" *) _04355_;
  assign _01491_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_38_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11675" *) _04358_;
  assign _01492_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_39_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11681" *) _04361_;
  assign _01493_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_40_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11687" *) _04364_;
  assign _01494_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_41_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11693" *) _04367_;
  assign _01495_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_42_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11700" *) _04370_;
  assign _01496_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_43_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11707" *) _04373_;
  assign _01497_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_44_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11714" *) _04376_;
  assign _01498_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_45_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11721" *) _04379_;
  assign _01499_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_46_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11728" *) _04382_;
  assign _01500_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_47_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11735" *) _04385_;
  assign _01501_ = IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11738" *) _04388_;
  assign _01502_ = _04054_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11759" *) IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm;
  assign _01503_ = _04055_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11765" *) IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm;
  assign _01504_ = _04056_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11771" *) IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm;
  assign _01505_ = _04057_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11777" *) IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm;
  assign _01506_ = _04058_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11783" *) IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm;
  assign _01507_ = _04059_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11789" *) IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm;
  assign _01508_ = _04060_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11795" *) IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm;
  assign _01509_ = _04061_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11801" *) IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm;
  assign _01510_ = _04062_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11810" *) IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm;
  assign _01511_ = _04063_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11816" *) IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm;
  assign _01512_ = _04064_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11825" *) IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm;
  assign _01513_ = _04065_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11831" *) IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm;
  assign _01514_ = _04066_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11837" *) IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm;
  assign _01515_ = _04067_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11843" *) IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm;
  assign _01516_ = _04068_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11849" *) cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2;
  assign _01517_ = _04069_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11855" *) cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2;
  assign cvt_1_FpMantRNE_17U_11U_else_and_tmp = FpMantRNE_17U_11U_else_carry_1_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11857" *) _03883_;
  assign cvt_2_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_2_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11859" *) _03884_;
  assign cvt_3_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_3_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11861" *) _03885_;
  assign cvt_4_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_4_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11863" *) _03886_;
  assign cvt_5_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_5_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11865" *) _03887_;
  assign cvt_6_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_6_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11867" *) _03888_;
  assign cvt_7_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_7_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11869" *) _03889_;
  assign cvt_8_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_8_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11871" *) _03890_;
  assign cvt_9_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_9_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11873" *) _03891_;
  assign cvt_10_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_10_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11875" *) _03892_;
  assign cvt_11_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_11_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11877" *) _03893_;
  assign cvt_12_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_12_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11879" *) _03894_;
  assign cvt_13_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_13_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11881" *) _03895_;
  assign cvt_14_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_14_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11883" *) _03896_;
  assign cvt_15_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_15_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11885" *) _03897_;
  assign cvt_16_FpMantRNE_17U_11U_else_and_4_tmp = FpMantRNE_17U_11U_else_carry_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11887" *) _03898_;
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11928" *) _05826_;
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11933" *) _04390_;
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11976" *) _05888_;
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11981" *) _04393_;
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12016" *) _05950_;
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12021" *) _04396_;
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12064" *) _06012_;
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12069" *) _04399_;
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12112" *) _06074_;
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12117" *) _04402_;
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12152" *) _06136_;
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12157" *) _04405_;
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12192" *) _06198_;
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12197" *) _04408_;
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12240" *) _06260_;
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12245" *) _04411_;
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12288" *) _06322_;
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12293" *) _04414_;
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12328" *) _06384_;
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12333" *) _04417_;
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12376" *) _06446_;
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12381" *) _04420_;
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_8_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12424" *) _06508_;
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12429" *) _04423_;
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12464" *) _06570_;
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12469" *) _04426_;
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12504" *) _06632_;
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12509" *) _04429_;
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12544" *) _06694_;
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12549" *) _04432_;
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_nl = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[62] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12584" *) _06756_;
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12589" *) _04435_;
  assign cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12608" *) _06786_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12613" *) _04438_;
  assign cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12636" *) _06817_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12641" *) _04441_;
  assign cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12664" *) _06848_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12669" *) _04444_;
  assign cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12692" *) _06879_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12697" *) _04447_;
  assign cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12720" *) _06910_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12725" *) _04450_;
  assign cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12748" *) _06941_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12753" *) _04453_;
  assign cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12776" *) _06972_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12781" *) _04456_;
  assign cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12804" *) _07003_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12809" *) _04459_;
  assign cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12832" *) _07034_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12837" *) _04462_;
  assign cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12860" *) _07065_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12865" *) _04465_;
  assign cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12888" *) _07096_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12893" *) _04468_;
  assign cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12916" *) _07127_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12921" *) _04471_;
  assign cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12944" *) _07158_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12949" *) _04474_;
  assign cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12972" *) _07189_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12977" *) _04477_;
  assign cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13000" *) _07220_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13005" *) _04480_;
  assign cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_8_nl = IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13028" *) _07251_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[44] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13033" *) _04483_;
  assign FpMantRNE_17U_11U_else_carry_1_sva = FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13048" *) _07257_;
  assign FpMantRNE_17U_11U_else_carry_2_sva = FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13057" *) _07262_;
  assign FpMantRNE_17U_11U_else_carry_3_sva = cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13066" *) _07267_;
  assign FpMantRNE_17U_11U_else_carry_4_sva = cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13075" *) _07272_;
  assign FpMantRNE_17U_11U_else_carry_5_sva = cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13084" *) _07277_;
  assign FpMantRNE_17U_11U_else_carry_6_sva = cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13093" *) _07282_;
  assign FpMantRNE_17U_11U_else_carry_7_sva = cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13102" *) _07287_;
  assign FpMantRNE_17U_11U_else_carry_8_sva = cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13111" *) _07292_;
  assign FpMantRNE_17U_11U_else_carry_9_sva = FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13120" *) _07297_;
  assign FpMantRNE_17U_11U_else_carry_10_sva = cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13129" *) _07302_;
  assign FpMantRNE_17U_11U_else_carry_11_sva = cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13138" *) _07307_;
  assign FpMantRNE_17U_11U_else_carry_12_sva = cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13147" *) _07312_;
  assign FpMantRNE_17U_11U_else_carry_13_sva = cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13156" *) _07317_;
  assign FpMantRNE_17U_11U_else_carry_14_sva = cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13165" *) _07322_;
  assign FpMantRNE_17U_11U_else_carry_15_sva = cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13174" *) _07327_;
  assign FpMantRNE_17U_11U_else_carry_sva = cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[5] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13183" *) _07332_;
  assign IntSaturation_17U_8U_and_1_nl = cvt_1_IntSaturation_17U_8U_else_if_acc_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13195" *) _04501_;
  assign IntSaturation_17U_8U_and_3_nl = cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13209" *) _04502_;
  assign IntSaturation_17U_8U_and_5_nl = cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13227" *) _04503_;
  assign IntSaturation_17U_8U_and_7_nl = cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13240" *) _04504_;
  assign IntSaturation_17U_8U_and_9_nl = cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13254" *) _04505_;
  assign IntSaturation_17U_8U_and_11_nl = cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13268" *) _04506_;
  assign IntSaturation_17U_8U_and_13_nl = cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13282" *) _04507_;
  assign IntSaturation_17U_8U_and_15_nl = cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13296" *) _04508_;
  assign IntSaturation_17U_8U_and_17_nl = cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13310" *) _04509_;
  assign IntSaturation_17U_8U_and_19_nl = cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13324" *) _04510_;
  assign IntSaturation_17U_8U_and_21_nl = cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13338" *) _04511_;
  assign IntSaturation_17U_8U_and_23_nl = cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13352" *) _04512_;
  assign IntSaturation_17U_8U_and_25_nl = cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13366" *) _04513_;
  assign IntSaturation_17U_8U_and_27_nl = cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13375" *) _04514_;
  assign IntSaturation_17U_8U_and_29_nl = cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13389" *) _04515_;
  assign IntSaturation_17U_8U_and_31_nl = cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13403" *) _04516_;
  assign cvt_and_147_m1c = _04517_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13412" *) cvt_unequal_tmp_21;
  assign main_stage_en_1 = chn_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13413" *) or_5189_cse;
  assign cvt_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl = _07351_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13530" *) _07353_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva = chn_idata_data_sva_1_27_0_1[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13535" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva = chn_idata_data_sva_1_27_0_1[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13540" *) cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva = chn_idata_data_sva_1_27_0_1[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13542" *) FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva[22:0];
  assign cvt_2_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = _07354_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13546" *) _07356_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva = chn_idata_data_sva_1_59_31_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13551" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva = chn_idata_data_sva_1_59_31_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13556" *) cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva = chn_idata_data_sva_1_59_31_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13558" *) FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva[22:0];
  assign cvt_3_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = _07357_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13562" *) _07359_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva = chn_idata_data_sva_1_91_63_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13567" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva = chn_idata_data_sva_1_91_63_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13572" *) cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva = chn_idata_data_sva_1_91_63_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13574" *) FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva[22:0];
  assign cvt_4_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = _07360_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13578" *) _07362_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_4_sva = chn_idata_data_sva_1_123_95_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13583" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_4_sva = chn_idata_data_sva_1_123_95_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13588" *) cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_4_sva = chn_idata_data_sva_1_123_95_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13590" *) FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva[22:0];
  assign cvt_5_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = _07363_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13594" *) _07365_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_5_sva = chn_idata_data_sva_1_155_127_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13599" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_5_sva = chn_idata_data_sva_1_155_127_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13604" *) cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_5_sva = chn_idata_data_sva_1_155_127_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13606" *) FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva[22:0];
  assign cvt_6_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = _07366_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13610" *) _07368_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_6_sva = chn_idata_data_sva_1_187_159_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13615" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_6_sva = chn_idata_data_sva_1_187_159_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13620" *) cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_6_sva = chn_idata_data_sva_1_187_159_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13622" *) FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva[22:0];
  assign cvt_7_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = _07369_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13626" *) _07371_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_7_sva = chn_idata_data_sva_1_219_191_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13631" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_7_sva = chn_idata_data_sva_1_219_191_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13636" *) cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_7_sva = chn_idata_data_sva_1_219_191_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13638" *) FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva[22:0];
  assign cvt_8_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = _07372_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13642" *) _07374_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_8_sva = chn_idata_data_sva_1_251_223_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13647" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_8_sva = chn_idata_data_sva_1_251_223_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13652" *) cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_8_sva = chn_idata_data_sva_1_251_223_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13654" *) FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva[22:0];
  assign cvt_9_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = _07375_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13658" *) _07377_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_9_sva = chn_idata_data_sva_1_283_255_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13663" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_9_sva = chn_idata_data_sva_1_283_255_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13668" *) cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_9_sva = chn_idata_data_sva_1_283_255_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13670" *) FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva[22:0];
  assign cvt_10_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = _07378_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13674" *) _07380_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_10_sva = chn_idata_data_sva_1_315_287_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13679" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_10_sva = chn_idata_data_sva_1_315_287_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13684" *) cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_10_sva = chn_idata_data_sva_1_315_287_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13686" *) FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva[22:0];
  assign cvt_11_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = _07381_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13690" *) _07383_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_11_sva = chn_idata_data_sva_1_347_319_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13695" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_11_sva = chn_idata_data_sva_1_347_319_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13700" *) cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_11_sva = chn_idata_data_sva_1_347_319_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13702" *) FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva[22:0];
  assign cvt_12_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = _07384_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13706" *) _07386_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_12_sva = chn_idata_data_sva_1_379_351_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13711" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_12_sva = chn_idata_data_sva_1_379_351_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13716" *) cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_12_sva = chn_idata_data_sva_1_379_351_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13718" *) FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva[22:0];
  assign cvt_13_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = _07387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13722" *) _07389_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_13_sva = chn_idata_data_sva_1_411_383_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13727" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_13_sva = chn_idata_data_sva_1_411_383_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13732" *) cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_13_sva = chn_idata_data_sva_1_411_383_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13734" *) FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva[22:0];
  assign cvt_14_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = _07390_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13738" *) _07392_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_14_sva = chn_idata_data_sva_1_443_415_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13743" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_14_sva = chn_idata_data_sva_1_443_415_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13748" *) cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_14_sva = chn_idata_data_sva_1_443_415_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13750" *) FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva[22:0];
  assign cvt_15_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = _07393_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13754" *) _07395_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_15_sva = chn_idata_data_sva_1_475_447_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13759" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_15_sva = chn_idata_data_sva_1_475_447_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13764" *) cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_15_sva = chn_idata_data_sva_1_475_447_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13766" *) FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva[22:0];
  assign cvt_16_FpMantDecShiftRight_23U_8U_10U_carry_and_4_nl = _07396_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13770" *) _07398_;
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva = chn_idata_data_sva_1_507_479_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13775" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva = chn_idata_data_sva_1_507_479_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13780" *) cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl;
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva = chn_idata_data_sva_1_507_479_1[23:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13782" *) FpMantDecShiftRight_23U_8U_10U_least_mask_sva[22:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13784" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13788" *) _03839_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13790" *) _04550_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13792" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13796" *) _03838_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13798" *) _04551_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13800" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13804" *) _03837_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13806" *) _04552_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13808" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13812" *) _03836_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13814" *) _04553_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13816" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13820" *) _03835_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13822" *) _04554_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13824" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13828" *) _03834_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13830" *) _04555_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13832" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13836" *) _03833_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13838" *) _04556_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13840" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13844" *) _03832_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13846" *) _04557_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13848" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13852" *) _03831_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13854" *) _04558_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13856" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13860" *) _03830_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13862" *) _04559_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13864" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13868" *) _03829_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13870" *) _04560_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13872" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13876" *) _03828_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13878" *) _04561_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13880" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13884" *) _03827_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13886" *) _04562_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13888" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13892" *) _03826_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13894" *) _04563_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13896" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13900" *) _03825_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13902" *) _04564_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13904" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13908" *) _03824_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13910" *) _04565_;
  assign _01518_ = cvt_if_unequal_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14072" *) _04517_;
  assign cvt_asn_321 = _01518_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14072" *) _04566_;
  assign _01519_ = cvt_else_nor_dfs & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14073" *) _04517_;
  assign cvt_asn_323 = _01519_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14073" *) cvt_unequal_tmp_21;
  assign _01520_ = cvt_else_equal_tmp_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14074" *) _04517_;
  assign cvt_asn_327 = _01520_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14074" *) cvt_unequal_tmp_21;
  assign _01521_ = cvt_else_nor_dfs_1_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14075" *) _04517_;
  assign cvt_asn_329 = _01521_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14075" *) cvt_unequal_tmp_21;
  assign _01522_ = cvt_else_equal_tmp_4_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14076" *) _04517_;
  assign cvt_asn_333 = _01522_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14076" *) cvt_unequal_tmp_21;
  assign _01523_ = cvt_else_nor_dfs_3_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14077" *) _04517_;
  assign cvt_asn_335 = _01523_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14077" *) cvt_unequal_tmp_21;
  assign _01524_ = cvt_else_equal_tmp_10_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14078" *) _04517_;
  assign cvt_asn_339 = _01524_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14078" *) cvt_unequal_tmp_21;
  assign _01525_ = cvt_else_nor_dfs_13_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14079" *) cvt_unequal_tmp_21;
  assign cvt_asn_341 = _01525_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14079" *) _04517_;
  assign _01526_ = cvt_else_equal_tmp_40_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14080" *) cvt_unequal_tmp_21;
  assign cvt_asn_345 = _01526_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14080" *) _04517_;
  assign _01527_ = cvt_else_nor_dfs_14_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14081" *) _04517_;
  assign cvt_asn_347 = _01527_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14081" *) cvt_unequal_tmp_21;
  assign _01528_ = cvt_else_equal_tmp_43_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14082" *) _04517_;
  assign cvt_asn_351 = _01528_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14082" *) cvt_unequal_tmp_21;
  assign _01529_ = cvt_else_nor_dfs_5_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14083" *) _04517_;
  assign cvt_asn_353 = _01529_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14083" *) cvt_unequal_tmp_21;
  assign _01530_ = cvt_else_equal_tmp_16_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14084" *) _04517_;
  assign cvt_asn_357 = _01530_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14084" *) cvt_unequal_tmp_21;
  assign _01531_ = cvt_else_nor_dfs_13_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14085" *) _04517_;
  assign cvt_asn_359 = _01531_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14085" *) cvt_unequal_tmp_21;
  assign _01532_ = cvt_else_equal_tmp_40_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14086" *) _04517_;
  assign cvt_asn_363 = _01532_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14086" *) cvt_unequal_tmp_21;
  assign _01533_ = cvt_else_nor_dfs_6_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14087" *) _04517_;
  assign cvt_asn_365 = _01533_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14087" *) cvt_unequal_tmp_21;
  assign _01534_ = cvt_else_equal_tmp_19_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14088" *) _04517_;
  assign cvt_asn_369 = _01534_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14088" *) cvt_unequal_tmp_21;
  assign _01535_ = cvt_else_nor_dfs_9_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14089" *) _04517_;
  assign cvt_asn_371 = _01535_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14089" *) cvt_unequal_tmp_21;
  assign _01536_ = cvt_else_equal_tmp_37_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14090" *) _04517_;
  assign cvt_asn_375 = _01536_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14090" *) cvt_unequal_tmp_21;
  assign cvt_asn_377 = cvt_else_nor_dfs_7_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14091" *) cvt_and_147_m1c;
  assign cvt_asn_381 = cvt_else_equal_tmp_22_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14092" *) cvt_and_147_m1c;
  assign _01537_ = cvt_else_nor_dfs_11_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14093" *) _04517_;
  assign cvt_asn_383 = _01537_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14093" *) cvt_unequal_tmp_21;
  assign _01538_ = cvt_else_equal_tmp_34_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14094" *) _04517_;
  assign cvt_asn_387 = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14094" *) cvt_unequal_tmp_21;
  assign _01539_ = cvt_else_nor_dfs_10_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14095" *) _04517_;
  assign cvt_asn_389 = _01539_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14095" *) cvt_unequal_tmp_21;
  assign _01540_ = cvt_else_equal_tmp_31_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14096" *) _04517_;
  assign cvt_asn_393 = _01540_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14096" *) cvt_unequal_tmp_21;
  assign _01541_ = cvt_else_equal_tmp_28_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14097" *) _04517_;
  assign cvt_asn_399 = _01541_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14097" *) cvt_unequal_tmp_21;
  assign and_dcpl_4 = and_dcpl_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14099" *) or_5189_cse;
  assign and_dcpl_70 = chn_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14100" *) cfg_proc_precision_rsci_d[1];
  assign and_dcpl_73 = chn_out_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14102" *) reg_chn_out_rsci_ld_core_psct_cse;
  assign and_tmp_8 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14117" *) mux_110_cse;
  assign and_tmp_11 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14118" *) or_4550_cse;
  assign and_tmp_12 = or_183_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14120" *) or_4550_cse;
  assign and_tmp_16 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14123" *) mux_tmp_117;
  assign and_2487_nl = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14127" *) main_stage_v_1;
  assign _01542_ = and_2487_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14127" *) mux_tmp_120;
  assign and_tmp_18 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14129" *) mux_tmp_120;
  assign and_tmp_19 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14133" *) mux_tmp_123;
  assign and_tmp_33 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14138" *) mux_148_nl;
  assign _01543_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14145" *) _04574_;
  assign _01544_ = cfg_proc_precision_1_sva_st_89[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14156" *) or_4862_cse;
  assign and_tmp_50 = or_4714_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14169" *) or_4862_cse;
  assign _01545_ = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14172" *) _07435_;
  assign and_tmp_52 = _01545_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14172" *) and_tmp_50;
  assign _01546_ = cfg_proc_precision_1_sva_st_64[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14174" *) or_513_cse;
  assign and_152_nl = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14177" *) mux_250_nl;
  assign and_153_nl = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14178" *) mux_tmp_249;
  assign _01547_ = cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14180" *) cfg_out_precision_1_sva_st_154[1];
  assign _01548_ = and_2487_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14200" *) and_tmp_12;
  assign and_tmp_67 = or_510_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14202" *) and_tmp_50;
  assign _01549_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14203" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign and_167_nl = or_510_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14208" *) mux_tmp_298;
  assign _01550_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14209" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign _01551_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14232" *) cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  assign and_tmp_71 = _01551_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14232" *) mux_tmp_120;
  assign _01552_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14241" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign and_176_nl = or_600_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14245" *) mux_tmp_298;
  assign _01553_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14246" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign and_tmp_79 = or_400_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14256" *) mux_1126_cse;
  assign _01554_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14257" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign and_181_nl = or_4536_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14260" *) mux_tmp_298;
  assign _01555_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14261" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign _01556_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14275" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign and_184_nl = or_4535_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14280" *) mux_tmp_298;
  assign _01557_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14281" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign _01558_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14297" *) or_183_cse_1;
  assign _01559_ = _01558_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14298" *) cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  assign and_tmp_93 = _01559_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14298" *) or_4550_cse;
  assign and_tmp_94 = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14301" *) mux_tmp_455;
  assign _01560_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14308" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign and_2218_nl = IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14311" *) mux_tmp_298;
  assign _01561_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14312" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign _01562_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14325" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign and_2214_nl = IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14328" *) mux_tmp_298;
  assign _01563_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14329" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign _01564_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14342" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign and_2210_nl = IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14345" *) mux_tmp_298;
  assign _01565_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14346" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign and_2209_nl = IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14351" *) main_stage_v_2;
  assign _01566_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14364" *) mux_1142_cse;
  assign and_2208_nl = IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14366" *) or_400_cse_1;
  assign and_2206_cse = IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14372" *) main_stage_v_2;
  assign _01567_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14373" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign and_2202_nl = IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14394" *) main_stage_v_2;
  assign and_2199_cse = IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14411" *) main_stage_v_2;
  assign _01568_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14412" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign and_2194_cse = IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14439" *) main_stage_v_2;
  assign _01569_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14440" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign _01570_ = cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14473" *) _03931_;
  assign _01571_ = _01570_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14473" *) mux_tmp_416;
  assign and_tmp_165 = or_3538_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14476" *) or_1159_cse;
  assign and_tmp_166 = or_3542_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14479" *) or_1159_cse;
  assign and_tmp_168 = or_3542_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14482" *) and_tmp_165;
  assign and_tmp_169 = or_3538_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14487" *) mux_969_nl;
  assign _01572_ = cfg_out_precision_1_sva_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14494" *) cfg_out_precision_1_sva_st_144[1];
  assign and_2247_nl = _04633_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14495" *) and_tmp_165;
  assign _01573_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14507" *) _04636_;
  assign and_tmp_171 = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14511" *) mux_tmp_1038;
  assign _01574_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14540" *) _04640_;
  assign and_tmp_175 = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14544" *) mux_tmp_1100;
  assign _01575_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14561" *) mux_tmp_1197;
  assign and_2246_cse = nand_190_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14600" *) or_tmp_2136;
  assign _01576_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14616" *) not_tmp_1709;
  assign and_306_nl = FpIntToFloat_17U_5U_10U_else_unequal_tmp_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14624" *) _04646_;
  assign _01577_ = cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14656" *) main_stage_v_1;
  assign _01578_ = _01577_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14656" *) and_dcpl_3;
  assign and_dcpl_93 = _04648_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14675" *) reg_chn_out_rsci_ld_core_psct_cse;
  assign _01579_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14677" *) _04566_;
  assign and_dcpl_98 = _01579_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14677" *) or_5189_cse;
  assign _01580_ = _04517_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14678" *) main_stage_v_3;
  assign and_dcpl_102 = _01580_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14678" *) or_5189_cse;
  assign and_dcpl_103 = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14679" *) main_stage_v_3;
  assign _01581_ = _04631_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14680" *) chn_out_rsci_bawt;
  assign and_dcpl_105 = _01581_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14680" *) reg_chn_out_rsci_ld_core_psct_cse;
  assign and_dcpl_114 = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14681" *) main_stage_v_1;
  assign _01582_ = _04649_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14684" *) main_stage_v_1;
  assign and_dcpl_204 = or_4550_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14686" *) or_5189_cse;
  assign and_dcpl_209 = _00187_[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14688" *) or_5189_cse;
  assign and_dcpl_217 = _00188_[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14690" *) or_5189_cse;
  assign and_dcpl_224 = _00189_[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14692" *) or_5189_cse;
  assign _01583_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14702" *) and_tmp_12;
  assign and_tmp_225 = or_400_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14706" *) mux_tmp_455;
  assign and_dcpl_301 = _00195_[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14713" *) or_5189_cse;
  assign and_dcpl_363 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14727" *) and_dcpl_228;
  assign and_dcpl_401 = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14735" *) main_stage_v_2;
  assign _01584_ = nor_50_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14736" *) cfg_out_precision_1_sva_st_113[0];
  assign _01585_ = _01584_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14737" *) or_5189_cse;
  assign and_dcpl_407 = _01585_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14737" *) _04650_;
  assign and_dcpl_408 = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14738" *) _04582_;
  assign and_dcpl_409 = or_dcpl_147 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14740" *) and_dcpl_408;
  assign _01586_ = or_4862_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14741" *) cvt_unequal_tmp_20;
  assign and_dcpl_411 = _01586_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14741" *) or_5189_cse;
  assign _01587_ = _04651_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14743" *) _04582_;
  assign and_dcpl_417 = _01587_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14743" *) or_5189_cse;
  assign and_dcpl_420 = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14744" *) cvt_unequal_tmp_20;
  assign and_dcpl_424 = or_4862_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14745" *) or_5189_cse;
  assign and_dcpl_425 = _07615_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14747" *) and_dcpl_420;
  assign _01588_ = nor_50_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14749" *) _03933_;
  assign and_dcpl_433 = _01588_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14749" *) and_dcpl_408;
  assign _01589_ = or_4862_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14750" *) _04652_;
  assign _01590_ = or_4862_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14752" *) and_dcpl_444;
  assign and_dcpl_446 = _01590_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14752" *) and_dcpl_420;
  assign and_dcpl_458 = and_dcpl_444 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14757" *) cvt_unequal_tmp_20;
  assign and_tmp_248 = or_5254_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14758" *) mux_tmp_987;
  assign and_dcpl_473 = and_tmp_225 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14760" *) or_5189_cse;
  assign and_dcpl_481 = and_dcpl_458 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14763" *) or_5189_cse;
  assign and_dcpl_499 = mux_tmp_455 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14766" *) or_5189_cse;
  assign _01591_ = or_1159_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14767" *) _04654_;
  assign _01592_ = _07618_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14778" *) or_1159_cse;
  assign _01593_ = _01592_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14778" *) or_3538_cse;
  assign _01594_ = _01593_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14778" *) or_3542_cse;
  assign and_dcpl_617 = _01594_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14778" *) and_dcpl_103;
  assign and_dcpl_626 = or_400_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14779" *) main_stage_v_2;
  assign _01595_ = _07619_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14781" *) or_1159_cse;
  assign _01596_ = _01595_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14782" *) or_3538_cse;
  assign _01597_ = _01596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14782" *) or_3542_cse;
  assign and_dcpl_631 = _01597_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14782" *) and_dcpl_103;
  assign _01598_ = _07620_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14783" *) or_1159_cse;
  assign _01599_ = _01598_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14784" *) or_3538_cse;
  assign _01600_ = _01599_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14784" *) or_3542_cse;
  assign _01601_ = _01600_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14784" *) or_5254_cse;
  assign and_dcpl_648 = _01601_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14784" *) and_dcpl_103;
  assign or_tmp_3487 = main_stage_en_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14851" *) fsm_output[1];
  assign _01602_ = _00063_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14853" *) main_stage_v_1;
  assign main_stage_v_1_mx0c1 = _01602_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14853" *) or_5189_cse;
  assign _01603_ = cvt_cvt_nand_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14854" *) chn_in_rsci_bawt;
  assign _01604_ = _04688_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14855" *) or_4550_cse;
  assign _01605_ = _01604_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14855" *) or_183_cse_1;
  assign IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 = _01605_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14855" *) and_dcpl_114;
  assign _01606_ = _04185_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14856" *) main_stage_v_2;
  assign main_stage_v_2_mx0c1 = _01606_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14856" *) or_5189_cse;
  assign _01607_ = _00058_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14857" *) main_stage_v_3;
  assign main_stage_v_3_mx0c1 = _01607_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14857" *) or_5189_cse;
  assign cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0 = _07645_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14860" *) and_dcpl_408;
  assign _01608_ = _04690_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14863" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1 = _01608_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14863" *) and_dcpl_417;
  assign and_2158_nl = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14864" *) nor_45_cse;
  assign cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0 = mux_1836_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14867" *) and_dcpl_408;
  assign _01609_ = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14870" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1 = _01609_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14870" *) and_dcpl_417;
  assign and_2157_nl = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14871" *) nor_45_cse;
  assign cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 = mux_1846_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14874" *) and_dcpl_408;
  assign _01610_ = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14877" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1 = _01610_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14877" *) and_dcpl_417;
  assign FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1 = _07646_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14879" *) and_dcpl_420;
  assign _01611_ = mux_tmp_321 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14881" *) _04691_;
  assign _01612_ = _01611_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14881" *) cvt_unequal_tmp_20;
  assign FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2 = _01612_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14881" *) or_5189_cse;
  assign cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0 = _07648_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14884" *) and_dcpl_408;
  assign _01613_ = _04693_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14887" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1 = _01613_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14887" *) and_dcpl_417;
  assign and_2155_nl = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14888" *) nor_45_cse;
  assign cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 = mux_1876_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14891" *) and_dcpl_408;
  assign _01614_ = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14894" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1 = _01614_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14894" *) and_dcpl_417;
  assign and_2152_nl = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14895" *) nor_45_cse;
  assign cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0 = mux_1903_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14898" *) and_dcpl_408;
  assign _01615_ = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14901" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1 = _01615_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14901" *) and_dcpl_417;
  assign and_2150_nl = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14902" *) nor_45_cse;
  assign cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 = mux_1927_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14905" *) and_dcpl_408;
  assign _01616_ = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14908" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1 = _01616_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14908" *) and_dcpl_417;
  assign and_2148_nl = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14909" *) nor_45_cse;
  assign cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0 = mux_1940_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14912" *) and_dcpl_408;
  assign _01617_ = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14915" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1 = _01617_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14915" *) and_dcpl_417;
  assign and_2147_nl = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14916" *) nor_45_cse;
  assign cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0 = mux_1943_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14919" *) and_dcpl_408;
  assign _01618_ = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14922" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1 = _01618_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14922" *) and_dcpl_417;
  assign and_2146_nl = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14923" *) nor_45_cse;
  assign cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 = mux_1953_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14926" *) and_dcpl_408;
  assign _01619_ = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14929" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1 = _01619_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14929" *) and_dcpl_417;
  assign and_2145_nl = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14930" *) nor_45_cse;
  assign cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 = mux_1964_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14933" *) and_dcpl_408;
  assign _01620_ = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14936" *) cfg_proc_precision_1_sva_st_65[1];
  assign cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1 = _01620_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14936" *) and_dcpl_417;
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16 = cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14938" *) IntShiftRightSat_49U_6U_17U_o_16_1_sva_3;
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14940" *) IntShiftRightSat_49U_6U_17U_o_16_2_sva_2;
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14942" *) IntShiftRightSat_49U_6U_17U_o_16_3_sva_3;
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14944" *) IntShiftRightSat_49U_6U_17U_o_16_4_sva_2;
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14946" *) IntShiftRightSat_49U_6U_17U_o_16_5_sva_3;
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14948" *) IntShiftRightSat_49U_6U_17U_o_16_6_sva_2;
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14950" *) IntShiftRightSat_49U_6U_17U_o_16_7_sva_2;
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14952" *) IntShiftRightSat_49U_6U_17U_o_16_8_sva_2;
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14954" *) IntShiftRightSat_49U_6U_17U_o_16_9_sva_3;
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14956" *) IntShiftRightSat_49U_6U_17U_o_16_10_sva_2;
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14958" *) IntShiftRightSat_49U_6U_17U_o_16_11_sva_2;
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14960" *) IntShiftRightSat_49U_6U_17U_o_16_12_sva_2;
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14962" *) IntShiftRightSat_49U_6U_17U_o_16_13_sva_2;
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14964" *) IntShiftRightSat_49U_6U_17U_o_16_14_sva_2;
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14966" *) IntShiftRightSat_49U_6U_17U_o_16_15_sva_2;
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16 = cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14968" *) IntShiftRightSat_49U_6U_17U_o_16_sva_2;
  assign _01621_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14990" *) or_400_cse_1;
  assign and_dcpl_1319 = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14995" *) core_wen;
  assign cvt_and_tmp_1 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14996" *) cvt_unequal_tmp_21;
  assign and_dcpl_1742 = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14997" *) core_wen;
  assign _01622_ = cvt_asn_323 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15057" *) _04699_;
  assign _01623_ = _01622_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15057" *) _04700_;
  assign _01624_ = cvt_asn_329 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15059" *) _04701_;
  assign _01625_ = _01624_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15059" *) _04702_;
  assign _01626_ = cvt_asn_323 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15061" *) _04703_;
  assign _01627_ = _01626_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15061" *) _04704_;
  assign _01628_ = cvt_asn_335 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15063" *) _04705_;
  assign _01629_ = _01628_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15063" *) _04706_;
  assign _01630_ = cvt_asn_323 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15065" *) _04707_;
  assign _01631_ = _01630_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15065" *) _04708_;
  assign _01632_ = cvt_asn_353 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15067" *) _04709_;
  assign _01633_ = _01632_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15067" *) _04710_;
  assign _01634_ = cvt_asn_365 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15069" *) _04711_;
  assign _01635_ = _01634_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15069" *) _04712_;
  assign _01636_ = cvt_asn_377 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15071" *) _04713_;
  assign _01637_ = _01636_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15071" *) _04714_;
  assign _01638_ = cvt_asn_323 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15073" *) _04715_;
  assign _01639_ = _01638_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15073" *) _04716_;
  assign _01640_ = cvt_asn_371 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15075" *) _04717_;
  assign _01641_ = _01640_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15075" *) _04718_;
  assign _01642_ = cvt_asn_389 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15077" *) _04719_;
  assign _01643_ = _01642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15077" *) _04720_;
  assign _01644_ = cvt_asn_383 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15079" *) _04721_;
  assign _01645_ = _01644_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15079" *) _04722_;
  assign _01646_ = cvt_asn_371 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15081" *) _04723_;
  assign _01647_ = _01646_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15081" *) _04724_;
  assign _01648_ = cvt_asn_359 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15083" *) _04725_;
  assign _01649_ = _01648_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15083" *) _04726_;
  assign _01650_ = cvt_asn_347 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15085" *) _04727_;
  assign _01651_ = _01650_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15085" *) _04728_;
  assign _01652_ = cvt_asn_341 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15087" *) _04729_;
  assign _01653_ = _01652_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15087" *) _04730_;
  assign _01654_ = _04731_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15094" *) fsm_output[1];
  assign _01655_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15102" *) chn_in_rsci_ld_core_psct_mx0c0;
  assign _01656_ = cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15332" *) cvt_unequal_tmp_21;
  assign _01657_ = cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15334" *) cvt_unequal_tmp_21;
  assign _01658_ = cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15336" *) cvt_unequal_tmp_21;
  assign _01659_ = cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15338" *) cvt_unequal_tmp_21;
  assign _01660_ = cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15340" *) cvt_unequal_tmp_21;
  assign _01661_ = cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15342" *) cvt_unequal_tmp_21;
  assign _01662_ = cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15344" *) cvt_unequal_tmp_21;
  assign _01663_ = cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15346" *) cvt_unequal_tmp_21;
  assign _01664_ = cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15348" *) cvt_unequal_tmp_21;
  assign _01665_ = cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15350" *) cvt_unequal_tmp_21;
  assign _01666_ = cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15352" *) cvt_unequal_tmp_21;
  assign _01667_ = cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15354" *) cvt_unequal_tmp_21;
  assign _01668_ = cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15356" *) cvt_unequal_tmp_21;
  assign _01669_ = cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15358" *) cvt_unequal_tmp_21;
  assign _01670_ = cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15360" *) cvt_unequal_tmp_21;
  assign _01671_ = cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15362" *) cvt_unequal_tmp_21;
  assign _01672_ = _07672_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15370" *) or_5189_cse;
  assign _01673_ = _01672_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15370" *) and_dcpl_1742;
  assign _01674_ = _07674_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15384" *) or_5189_cse;
  assign _01675_ = _01674_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15384" *) and_dcpl_1742;
  assign _01676_ = _07676_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15397" *) or_5189_cse;
  assign _01677_ = _01676_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15397" *) and_dcpl_1742;
  assign _01678_ = _07678_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15411" *) or_5189_cse;
  assign _01679_ = _01678_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15411" *) and_dcpl_1742;
  assign _01680_ = _07680_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15425" *) or_5189_cse;
  assign _01681_ = _01680_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15425" *) and_dcpl_1742;
  assign _01682_ = _07682_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15439" *) or_5189_cse;
  assign _01683_ = _01682_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15439" *) and_dcpl_1742;
  assign _01684_ = _07684_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15453" *) or_5189_cse;
  assign _01685_ = _01684_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15453" *) and_dcpl_1742;
  assign _01686_ = _07686_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15467" *) or_5189_cse;
  assign _01687_ = _01686_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15467" *) and_dcpl_1742;
  assign _01688_ = _07688_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15481" *) or_5189_cse;
  assign _01689_ = _01688_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15481" *) and_dcpl_1742;
  assign _01690_ = _07690_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15515" *) or_5189_cse;
  assign _01691_ = _01690_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15515" *) and_dcpl_1742;
  assign _01692_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15621" *) _07691_;
  assign _01693_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15629" *) _07692_;
  assign _01694_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15637" *) mux_nl;
  assign _01695_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15645" *) mux_5_nl;
  assign _01696_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15654" *) _04744_;
  assign _01697_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15664" *) _04745_;
  assign _01698_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15673" *) mux_11_nl;
  assign _01699_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15726" *) _04746_;
  assign _01700_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15736" *) _04747_;
  assign _01701_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15745" *) mux_17_nl;
  assign _01702_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15754" *) _04748_;
  assign _01703_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15764" *) _04749_;
  assign _01704_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15773" *) mux_22_nl;
  assign _01705_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15782" *) _04750_;
  assign _01706_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15792" *) _04751_;
  assign _01707_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15801" *) _04752_;
  assign _01708_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15810" *) _04753_;
  assign _01709_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15820" *) _04754_;
  assign _01710_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15829" *) _04755_;
  assign _01711_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15838" *) _04756_;
  assign _01712_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15848" *) _04757_;
  assign _01713_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15857" *) _04758_;
  assign _01714_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15866" *) _04759_;
  assign _01715_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15876" *) _04760_;
  assign _01716_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15885" *) mux_45_nl;
  assign _01717_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15894" *) _04761_;
  assign _01718_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15904" *) _04762_;
  assign _01719_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15913" *) mux_50_nl;
  assign _01720_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15922" *) _04763_;
  assign _01721_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15932" *) _04764_;
  assign _01722_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15941" *) _04765_;
  assign _01723_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15950" *) _04766_;
  assign _01724_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15960" *) _04767_;
  assign _01725_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15969" *) mux_61_nl;
  assign _01726_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15978" *) _04768_;
  assign _01727_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15988" *) _04769_;
  assign _01728_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15997" *) mux_66_nl;
  assign _01729_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16006" *) _04770_;
  assign _01730_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16016" *) _04771_;
  assign _01731_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16025" *) _04772_;
  assign _01732_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16034" *) _04773_;
  assign _01733_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16044" *) _04774_;
  assign _01734_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16053" *) mux_77_nl;
  assign _01735_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16062" *) _04775_;
  assign _01736_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16072" *) _04776_;
  assign _01737_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16081" *) mux_82_nl;
  assign _01738_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16090" *) _04777_;
  assign _01739_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16100" *) _04778_;
  assign _01740_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16109" *) mux_87_nl;
  assign _01741_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16118" *) _04779_;
  assign _01742_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16128" *) _04780_;
  assign _01743_ = _03935_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16304" *) FpMantRNE_24U_11U_else_mux_31_nl;
  assign _01744_ = _01743_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8];
  assign _01745_ = _01744_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *) _04781_;
  assign _01746_ = _03936_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16312" *) FpMantRNE_24U_11U_else_mux_29_nl;
  assign _01747_ = _01746_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _01748_ = _01747_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *) _04783_;
  assign _01749_ = _03937_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16320" *) FpMantRNE_24U_11U_else_mux_27_nl;
  assign _01750_ = _01749_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _01751_ = _01750_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *) _04785_;
  assign _01752_ = _03938_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16328" *) FpMantRNE_24U_11U_else_mux_25_nl;
  assign _01753_ = _01752_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _01754_ = _01753_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *) _04787_;
  assign _01755_ = _03939_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16336" *) FpMantRNE_24U_11U_else_mux_23_nl;
  assign _01756_ = _01755_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _01757_ = _01756_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *) _04789_;
  assign _01758_ = _03940_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16344" *) FpMantRNE_24U_11U_else_mux_21_nl;
  assign _01759_ = _01758_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _01760_ = _01759_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *) _04791_;
  assign _01761_ = _03941_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16352" *) FpMantRNE_24U_11U_else_mux_19_nl;
  assign _01762_ = _01761_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _01763_ = _01762_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *) _04793_;
  assign _01764_ = _03942_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16360" *) FpMantRNE_24U_11U_else_mux_17_nl;
  assign _01765_ = _01764_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _01766_ = _01765_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *) _04795_;
  assign _01767_ = _03943_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16368" *) FpMantRNE_24U_11U_else_mux_15_nl;
  assign _01768_ = _01767_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _01769_ = _01768_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *) _04797_;
  assign _01770_ = _03944_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16376" *) FpMantRNE_24U_11U_else_mux_13_nl;
  assign _01771_ = _01770_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _01772_ = _01771_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *) _04799_;
  assign _01773_ = _03945_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16384" *) FpMantRNE_24U_11U_else_mux_11_nl;
  assign _01774_ = _01773_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _01775_ = _01774_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *) _04801_;
  assign _01776_ = _03946_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16393" *) FpMantRNE_24U_11U_else_mux_9_nl;
  assign _01777_ = _01776_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _01778_ = _01777_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *) _04803_;
  assign _01779_ = _03947_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16401" *) FpMantRNE_24U_11U_else_mux_7_nl;
  assign _01780_ = _01779_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _01781_ = _01780_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *) _04805_;
  assign _01782_ = _03948_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16409" *) FpMantRNE_24U_11U_else_mux_5_nl;
  assign _01783_ = _01782_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _01784_ = _01783_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *) _04807_;
  assign _01785_ = _03949_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16417" *) FpMantRNE_24U_11U_else_mux_3_nl;
  assign _01786_ = _01785_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _01787_ = _01786_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *) _04809_;
  assign _01788_ = _03950_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16425" *) FpMantRNE_24U_11U_else_mux_1_nl;
  assign _01789_ = _01788_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8];
  assign _01790_ = _01789_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *) _04811_;
  assign _01791_ = and_2186_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16448" *) and_dcpl_73;
  assign _01792_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16449" *) _07694_;
  assign _01793_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16494" *) mux_tmp_122;
  assign _01794_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16503" *) mux_159_nl;
  assign _01795_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16522" *) _07695_;
  assign _01796_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *) _03951_;
  assign _01797_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *) _03952_;
  assign _01798_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *) _03953_;
  assign _01799_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *) _03954_;
  assign _01800_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *) _03955_;
  assign _01801_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *) _03956_;
  assign _01802_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *) _03957_;
  assign _01803_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *) _03958_;
  assign _01804_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *) _03959_;
  assign _01805_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *) _03960_;
  assign _01806_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *) _03961_;
  assign _01807_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *) _03962_;
  assign _01808_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *) _03963_;
  assign _01809_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16717" *) IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  assign _01810_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16718" *) _07709_;
  assign _01811_ = _01810_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16718" *) mux_tmp_161;
  assign _01812_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16728" *) mux_162_nl;
  assign _01813_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16736" *) IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  assign _01814_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16737" *) _07710_;
  assign _01815_ = _01814_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16737" *) mux_tmp_161;
  assign _01816_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16759" *) IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  assign _01817_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16760" *) _07711_;
  assign _01818_ = _01817_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16760" *) mux_tmp_161;
  assign _01819_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16770" *) IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  assign _01820_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16771" *) _07712_;
  assign _01821_ = _01820_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16771" *) mux_tmp_161;
  assign _01822_ = nor_1099_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16781" *) or_5189_cse;
  assign _01823_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16781" *) _07713_;
  assign _01824_ = _01823_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16782" *) mux_tmp_161;
  assign _01825_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16792" *) _04853_;
  assign _01826_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16800" *) IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  assign _01827_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16801" *) _07714_;
  assign _01828_ = _01827_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16801" *) mux_tmp_161;
  assign _01829_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16831" *) IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  assign _01830_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16832" *) _07715_;
  assign _01831_ = _01830_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16832" *) mux_tmp_161;
  assign _01832_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16842" *) IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  assign _01833_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16843" *) _07716_;
  assign _01834_ = _01833_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16843" *) mux_tmp_161;
  assign _01835_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16853" *) IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  assign _01836_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16854" *) _07717_;
  assign _01837_ = _01836_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16854" *) mux_tmp_161;
  assign _01838_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16876" *) IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  assign _01839_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16877" *) _07718_;
  assign _01840_ = _01839_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16877" *) mux_tmp_161;
  assign _01841_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16887" *) IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  assign _01842_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16888" *) _07719_;
  assign _01843_ = _01842_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16888" *) mux_tmp_161;
  assign _01844_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16898" *) IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  assign _01845_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16899" *) _07720_;
  assign _01846_ = _01845_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16899" *) mux_tmp_161;
  assign _01847_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16909" *) IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  assign _01848_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16910" *) _07721_;
  assign _01849_ = _01848_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16910" *) mux_tmp_161;
  assign _01850_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16920" *) IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  assign _01851_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16921" *) _07722_;
  assign _01852_ = _01851_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16921" *) mux_tmp_161;
  assign _01853_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16931" *) IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  assign _01854_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16932" *) _07723_;
  assign _01855_ = _01854_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16932" *) mux_tmp_161;
  assign _01856_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16942" *) _04854_;
  assign _01857_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16950" *) IsNaN_8U_23U_land_lpi_1_dfm_3;
  assign _01858_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16951" *) _07724_;
  assign _01859_ = _01858_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16951" *) mux_tmp_161;
  assign _01860_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16961" *) _04855_;
  assign _01861_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16969" *) mux_235_nl;
  assign _01862_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16978" *) IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse;
  assign _01863_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16978" *) mux_243_nl;
  assign _01864_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17000" *) _04856_;
  assign _01865_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17009" *) mux_247_nl;
  assign _01866_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17017" *) mux_248_nl;
  assign _01867_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17026" *) IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse;
  assign _01868_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17026" *) mux_257_nl;
  assign _01869_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17036" *) mux_267_nl;
  assign _01870_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17058" *) not_tmp_249;
  assign _01871_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17068" *) mux_271_nl;
  assign _01872_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17091" *) mux_275_nl;
  assign _01873_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17100" *) mux_285_nl;
  assign _01874_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17122" *) not_tmp_269;
  assign _01875_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17132" *) mux_289_nl;
  assign _01876_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17141" *) mux_291_nl;
  assign _01877_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17150" *) mux_302_nl;
  assign _01878_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17160" *) mux_316_nl;
  assign _01879_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *) _04857_;
  assign _01880_ = _01879_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *) or_dcpl_108;
  assign _01881_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *) _07725_;
  assign _01882_ = _01881_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *) not_tmp_312;
  assign _01883_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17220" *) not_tmp_312;
  assign _01884_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17230" *) mux_322_nl;
  assign _01885_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17239" *) mux_329_nl;
  assign _01886_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17248" *) mux_338_nl;
  assign _01887_ = _04858_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17257" *) core_wen;
  assign _01888_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *) _04859_;
  assign _01889_ = _01888_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *) or_dcpl_110;
  assign _01890_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *) _07727_;
  assign _01891_ = _01890_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *) not_tmp_336;
  assign _01892_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17276" *) not_tmp_336;
  assign _01893_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17286" *) mux_342_nl;
  assign _01894_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17295" *) mux_348_nl;
  assign _01895_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17304" *) mux_359_nl;
  assign _01896_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17314" *) mux_373_nl;
  assign _01897_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *) _04860_;
  assign _01898_ = _01897_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *) or_dcpl_113;
  assign _01899_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *) _07728_;
  assign _01900_ = _01899_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *) not_tmp_388;
  assign _01901_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17344" *) not_tmp_388;
  assign _01902_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17367" *) mux_383_nl;
  assign _01903_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17376" *) mux_394_nl;
  assign _01904_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17386" *) mux_408_nl;
  assign _01905_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *) _04861_;
  assign _01906_ = _01905_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *) or_dcpl_115;
  assign _01907_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *) _07729_;
  assign _01908_ = _01907_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *) not_tmp_436;
  assign _01909_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17406" *) not_tmp_436;
  assign _01910_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17415" *) mux_418_nl;
  assign _01911_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17424" *) mux_431_nl;
  assign _01912_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17434" *) mux_444_nl;
  assign _01913_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *) _04863_;
  assign _01914_ = _01913_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *) or_dcpl_119;
  assign _01915_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *) _07731_;
  assign _01916_ = _01915_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *) not_tmp_497;
  assign _01917_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17462" *) not_tmp_497;
  assign _01918_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17472" *) mux_450_nl;
  assign _01919_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17482" *) mux_453_nl;
  assign _01920_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17491" *) mux_458_nl;
  assign _01921_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17500" *) mux_467_nl;
  assign _01922_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17522" *) not_tmp_520;
  assign _01923_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17532" *) mux_472_nl;
  assign _01924_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17541" *) mux_478_nl;
  assign _01925_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17550" *) mux_490_nl;
  assign _01926_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17560" *) mux_505_nl;
  assign _01927_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *) _04864_;
  assign _01928_ = _01927_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *) or_dcpl_124;
  assign _01929_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *) _07732_;
  assign _01930_ = _01929_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *) not_tmp_580;
  assign _01931_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17580" *) not_tmp_580;
  assign _01932_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17589" *) mux_516_nl;
  assign _01933_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17598" *) mux_528_nl;
  assign _01934_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17608" *) mux_544_nl;
  assign _01935_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *) _04865_;
  assign _01936_ = _01935_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *) or_dcpl_126;
  assign _01937_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *) _07733_;
  assign _01938_ = _01937_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *) not_tmp_638;
  assign _01939_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17628" *) not_tmp_638;
  assign _01940_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17637" *) mux_556_nl;
  assign _01941_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17646" *) mux_569_nl;
  assign _01942_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17656" *) mux_583_nl;
  assign _01943_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *) _04866_;
  assign _01944_ = _01943_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *) or_dcpl_130;
  assign _01945_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *) _07734_;
  assign _01946_ = _01945_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *) _04867_;
  assign _01947_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17686" *) _04867_;
  assign _01948_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17695" *) mux_594_nl;
  assign _01949_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17704" *) mux_605_nl;
  assign _01950_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17714" *) mux_617_nl;
  assign _01951_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *) _04868_;
  assign _01952_ = _01951_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *) or_dcpl_132;
  assign _01953_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *) _07735_;
  assign _01954_ = _01953_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *) not_tmp_757;
  assign _01955_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17734" *) not_tmp_757;
  assign _01956_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17743" *) mux_630_nl;
  assign _01957_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17764" *) mux_644_nl;
  assign and_676_cse = and_tmp_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17773" *) or_5189_cse;
  assign _01958_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17773" *) main_stage_v_1;
  assign _01959_ = _01958_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17774" *) and_dcpl_228;
  assign _01960_ = _01959_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17774" *) core_wen;
  assign _01961_ = _07736_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17782" *) core_wen;
  assign _01962_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *) _04869_;
  assign _01963_ = _01962_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *) or_dcpl_136;
  assign _01964_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *) _07737_;
  assign _01965_ = _01964_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *) not_tmp_811;
  assign _01966_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17801" *) not_tmp_811;
  assign _01967_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17810" *) mux_671_nl;
  assign _01968_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17819" *) mux_684_nl;
  assign _01969_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17829" *) mux_698_nl;
  assign _01970_ = _04870_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17838" *) core_wen;
  assign _01971_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *) _04871_;
  assign _01972_ = _01971_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *) or_dcpl_139;
  assign _01973_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *) _07739_;
  assign _01974_ = _01973_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *) not_tmp_899;
  assign _01975_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17857" *) not_tmp_899;
  assign _01976_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17866" *) mux_715_nl;
  assign _01977_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17875" *) mux_730_nl;
  assign _01978_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17885" *) mux_746_nl;
  assign _01979_ = _04872_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17894" *) core_wen;
  assign _01980_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *) _04873_;
  assign _01981_ = _01980_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *) or_dcpl_143;
  assign _01982_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *) _07741_;
  assign _01983_ = _01982_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *) not_tmp_989;
  assign _01984_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17913" *) not_tmp_989;
  assign _01985_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17922" *) mux_794_nl;
  assign _01986_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17954" *) _07742_;
  assign _01987_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18029" *) _07744_;
  assign _01988_ = _01987_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18030" *) mux_811_nl;
  assign _01989_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18041" *) mux_815_nl;
  assign _01990_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18136" *) _07746_;
  assign _01991_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18149" *) mux_822_nl;
  assign IsNaN_5U_10U_aelse_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18157" *) IsNaN_5U_10U_aelse_or_cse;
  assign _01992_ = IsNaN_5U_10U_aelse_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18157" *) mux_829_nl;
  assign _01993_ = mux_2224_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18166" *) or_5189_cse;
  assign _01994_ = _01993_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18166" *) core_wen;
  assign _01996_ = _07748_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *) or_5189_cse;
  assign _01997_ = _01996_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *) core_wen;
  assign _01998_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18186" *) _07750_;
  assign _01999_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18199" *) mux_833_nl;
  assign _02000_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18283" *) _07752_;
  assign _02001_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18296" *) mux_837_nl;
  assign _02002_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18305" *) _07754_;
  assign _02003_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18340" *) mux_841_nl;
  assign _02004_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18349" *) _07756_;
  assign _02005_ = _02004_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18350" *) mux_849_nl;
  assign _02006_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18361" *) mux_853_nl;
  assign _02007_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18369" *) _07757_;
  assign _02008_ = _02007_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18369" *) mux_859_nl;
  assign _02009_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18381" *) _07759_;
  assign _02010_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18414" *) mux_863_nl;
  assign _02011_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18425" *) _07761_;
  assign _02012_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18438" *) mux_867_nl;
  assign _02013_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18473" *) _07763_;
  assign _02014_ = _02013_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18474" *) mux_875_nl;
  assign _02015_ = _03933_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18485" *) and_2360_cse;
  assign _02016_ = _07764_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18486" *) or_5189_cse;
  assign _02017_ = _02016_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18486" *) core_wen;
  assign _02018_ = _07766_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18495" *) or_5189_cse;
  assign _02019_ = _02018_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18495" *) core_wen;
  assign _02020_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18503" *) mux_879_nl;
  assign _02021_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18512" *) _07768_;
  assign _02022_ = _02021_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18513" *) mux_887_nl;
  assign _02023_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18524" *) mux_891_nl;
  assign IsNaN_5U_10U_aelse_and_1_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18532" *) IsNaN_5U_10U_aelse_or_1_cse;
  assign _02024_ = IsNaN_5U_10U_aelse_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18532" *) _04875_;
  assign _02025_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18544" *) _07770_;
  assign _02026_ = IsNaN_5U_10U_aelse_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18557" *) mux_909_nl;
  assign _02027_ = mux_2237_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18567" *) or_5189_cse;
  assign _02028_ = _02027_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18567" *) core_wen;
  assign _02029_ = _07771_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18575" *) or_5189_cse;
  assign _02030_ = _02029_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18575" *) core_wen;
  assign _02031_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18583" *) mux_913_nl;
  assign _02032_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18592" *) _07773_;
  assign _02033_ = _02032_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18593" *) mux_921_nl;
  assign _02034_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18604" *) mux_925_nl;
  assign _02035_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18615" *) _07775_;
  assign _02036_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18628" *) mux_929_nl;
  assign _02037_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18639" *) _07777_;
  assign _02038_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18652" *) mux_933_nl;
  assign _02039_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18663" *) _07779_;
  assign _02040_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18676" *) mux_937_nl;
  assign _02041_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18687" *) _07781_;
  assign _02042_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18703" *) _07783_;
  assign _02043_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18810" *) mux_943_nl;
  assign _02044_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18883" *) _04892_;
  assign _02045_ = _02044_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18883" *) _04893_;
  assign _02046_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18891" *) mux_959_nl;
  assign _02047_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18900" *) _04894_;
  assign _02048_ = _02047_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18900" *) _04895_;
  assign _02049_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18908" *) mux_982_nl;
  assign _02050_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18938" *) reg_cvt_else_cvt_else_nor_4_cse;
  assign _02051_ = _02050_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18939" *) _04896_;
  assign _02052_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18959" *) _04897_;
  assign _02053_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18967" *) mux_1000_nl;
  assign _02054_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18987" *) mux_1004_nl;
  assign _02055_ = _04898_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18989" *) FpMantRNE_17U_11U_else_mux_1_nl;
  assign _02056_ = _04899_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18989" *) FpIntToFloat_17U_5U_10U_else_mux_1_nl;
  assign _02057_ = mux_2250_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *) or_4862_cse;
  assign _02058_ = _02057_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *) core_wen;
  assign _02059_ = _02058_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *) _04901_;
  assign _02060_ = _02059_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18998" *) main_stage_v_2;
  assign _02061_ = _02060_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18998" *) _03931_;
  assign _02062_ = _02061_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18999" *) _04902_;
  assign _02063_ = _02062_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19000" *) _04903_;
  assign _02064_ = _02063_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19000" *) or_5189_cse;
  assign _02065_ = _02064_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19000" *) cvt_unequal_tmp_20;
  assign _02066_ = mux_2251_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19008" *) core_wen;
  assign _02067_ = _02066_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19008" *) _04901_;
  assign _02068_ = _02067_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19009" *) main_stage_v_2;
  assign _02069_ = _02068_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19009" *) or_5189_cse;
  assign _02070_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19018" *) mux_1011_nl;
  assign _02071_ = and_tmp_50 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19027" *) and_dcpl_401;
  assign _02072_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19027" *) _07804_;
  assign _02073_ = _02072_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19028" *) _04904_;
  assign _02074_ = mux_2252_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19037" *) or_4714_cse;
  assign _02075_ = _02074_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19037" *) or_4862_cse;
  assign _02076_ = _02075_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19037" *) core_wen;
  assign _02077_ = _02076_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *) _04901_;
  assign _02078_ = _02077_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *) main_stage_v_2;
  assign _02079_ = _02078_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *) _03931_;
  assign _02080_ = _02079_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19039" *) _04905_;
  assign _02081_ = _02080_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *) _04906_;
  assign _02082_ = _02081_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *) _03980_;
  assign _02083_ = _02082_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *) or_5189_cse;
  assign _02084_ = _02083_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19041" *) cvt_unequal_tmp_20;
  assign _02085_ = mux_2253_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19049" *) _04901_;
  assign _02086_ = _02085_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19049" *) main_stage_v_2;
  assign _02087_ = _02086_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19050" *) core_wen;
  assign _02088_ = _02087_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19050" *) or_5189_cse;
  assign _02089_ = _04907_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19061" *) FpMantRNE_17U_11U_else_mux_5_nl;
  assign _02090_ = _04908_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19061" *) FpIntToFloat_17U_5U_10U_else_mux_7_nl;
  assign _02091_ = _04910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19064" *) FpMantRNE_17U_11U_else_mux_9_nl;
  assign _02092_ = _04911_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19064" *) FpIntToFloat_17U_5U_10U_else_mux_13_nl;
  assign _02093_ = mux_2254_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19072" *) or_4714_cse;
  assign _02094_ = _02093_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19072" *) or_4862_cse;
  assign _02095_ = _02094_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19072" *) core_wen;
  assign _02096_ = _02095_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *) _04901_;
  assign _02097_ = _02096_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *) main_stage_v_2;
  assign _02098_ = _02097_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *) _03931_;
  assign _02099_ = _02098_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19074" *) _04913_;
  assign _02100_ = _02099_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19075" *) _04914_;
  assign _02101_ = _02100_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19075" *) _03980_;
  assign _02102_ = _02101_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19075" *) or_5189_cse;
  assign _02103_ = _02102_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19076" *) cvt_unequal_tmp_20;
  assign _02104_ = mux_2255_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19084" *) _04901_;
  assign _02105_ = _02104_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19084" *) main_stage_v_2;
  assign _02106_ = _02105_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19085" *) core_wen;
  assign _02107_ = _02106_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19085" *) or_5189_cse;
  assign _02108_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19094" *) mux_1035_nl;
  assign _02109_ = mux_tmp_321 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19103" *) and_dcpl_401;
  assign _02110_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19103" *) _07807_;
  assign _02111_ = _02110_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19104" *) _04915_;
  assign _02112_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19113" *) mux_2256_nl;
  assign _02113_ = _02112_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19113" *) or_400_cse_1;
  assign _02114_ = _02113_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19113" *) or_4714_cse;
  assign _02115_ = _02114_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *) or_4862_cse;
  assign _02116_ = _02115_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *) core_wen;
  assign _02117_ = _02116_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *) _04901_;
  assign _02118_ = _02117_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19114" *) main_stage_v_2;
  assign _02119_ = _02118_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19115" *) _03931_;
  assign _02120_ = _02119_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19116" *) _04916_;
  assign _02121_ = _02120_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19116" *) _04917_;
  assign _02122_ = _02121_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19117" *) _03980_;
  assign _02123_ = _02122_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19117" *) or_5189_cse;
  assign _02124_ = mux_2257_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19125" *) and_dcpl_1319;
  assign _02125_ = _02124_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19125" *) _04901_;
  assign _02126_ = _02125_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19126" *) or_5189_cse;
  assign _02127_ = mux_2258_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19134" *) or_4714_cse;
  assign _02128_ = _02127_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19134" *) or_4862_cse;
  assign _02129_ = _02128_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19134" *) core_wen;
  assign _02130_ = _02129_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *) _04901_;
  assign _02131_ = _02130_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *) main_stage_v_2;
  assign _02132_ = _02131_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *) _03931_;
  assign _02133_ = _02132_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19136" *) _04918_;
  assign _02134_ = _02133_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19137" *) _04647_;
  assign _02135_ = _02134_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19137" *) _03980_;
  assign _02136_ = _02135_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19137" *) or_5189_cse;
  assign _02137_ = _02136_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19138" *) cvt_unequal_tmp_20;
  assign _02138_ = mux_2259_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19146" *) _04901_;
  assign _02139_ = _02138_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19146" *) main_stage_v_2;
  assign _02140_ = _02139_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19147" *) core_wen;
  assign _02141_ = _02140_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19147" *) or_5189_cse;
  assign _02142_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19156" *) mux_1070_nl;
  assign _02143_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19166" *) FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse;
  assign _02144_ = _02143_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19166" *) _04919_;
  assign _02145_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19175" *) mux_2260_nl;
  assign _02146_ = _02145_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19175" *) or_400_cse_1;
  assign _02147_ = _02146_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19175" *) or_4714_cse;
  assign _02148_ = _02147_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *) or_4862_cse;
  assign _02149_ = _02148_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *) core_wen;
  assign _02150_ = _02149_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *) _04901_;
  assign _02151_ = _02150_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19176" *) main_stage_v_2;
  assign _02152_ = _02151_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19177" *) _03931_;
  assign _02153_ = _02152_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19178" *) _04920_;
  assign _02154_ = _02153_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19178" *) _04921_;
  assign _02155_ = _02154_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19179" *) _03980_;
  assign _02156_ = _02155_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19179" *) or_5189_cse;
  assign _02157_ = mux_2261_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19187" *) main_stage_v_2;
  assign _02158_ = _02157_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19187" *) _04901_;
  assign _02159_ = _02158_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19188" *) core_wen;
  assign _02160_ = _02159_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19188" *) or_5189_cse;
  assign _02161_ = _02143_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19197" *) _04922_;
  assign _02162_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19206" *) mux_2262_nl;
  assign _02163_ = _02162_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19206" *) or_400_cse_1;
  assign _02164_ = _02163_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19206" *) or_4714_cse;
  assign _02165_ = _02164_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *) or_4862_cse;
  assign _02166_ = _02165_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *) core_wen;
  assign _02167_ = _02166_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *) _04901_;
  assign _02168_ = _02167_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19207" *) main_stage_v_2;
  assign _02169_ = _02168_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19208" *) _03931_;
  assign _02170_ = _02169_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19209" *) _04923_;
  assign _02171_ = _02170_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19209" *) _04924_;
  assign _02172_ = _02171_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19210" *) _03980_;
  assign _02173_ = _02172_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19210" *) or_5189_cse;
  assign _02174_ = mux_2263_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19218" *) main_stage_v_2;
  assign _02175_ = _02174_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19218" *) _04901_;
  assign _02176_ = _02175_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19219" *) core_wen;
  assign _02177_ = _02176_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19219" *) or_5189_cse;
  assign _02178_ = _02143_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19228" *) _04925_;
  assign _02179_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19237" *) mux_2264_nl;
  assign _02180_ = _02179_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19237" *) or_400_cse_1;
  assign _02181_ = _02180_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19237" *) or_4714_cse;
  assign _02182_ = _02181_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *) or_4862_cse;
  assign _02183_ = _02182_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *) core_wen;
  assign _02184_ = _02183_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *) _04901_;
  assign _02185_ = _02184_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19238" *) main_stage_v_2;
  assign _02186_ = _02185_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19239" *) _03931_;
  assign _02187_ = _02186_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19240" *) _04926_;
  assign _02188_ = _02187_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19240" *) _04927_;
  assign _02189_ = _02188_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19241" *) _03980_;
  assign _02190_ = _02189_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19241" *) or_5189_cse;
  assign _02191_ = mux_2265_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19249" *) _04901_;
  assign _02192_ = _02191_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19249" *) core_wen;
  assign _02193_ = _02192_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19250" *) main_stage_v_2;
  assign _02194_ = _02193_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19250" *) or_5189_cse;
  assign _02195_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19258" *) mux_1127_nl;
  assign _02196_ = _04928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19260" *) FpMantRNE_17U_11U_else_mux_17_nl;
  assign _02197_ = _04929_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19260" *) FpIntToFloat_17U_5U_10U_else_mux_25_nl;
  assign _02198_ = mux_2266_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19268" *) or_4714_cse;
  assign _02199_ = _02198_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19268" *) or_4862_cse;
  assign _02200_ = _02199_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19268" *) core_wen;
  assign _02201_ = _02200_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *) _04901_;
  assign _02202_ = _02201_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *) main_stage_v_2;
  assign _02203_ = _02202_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *) _03931_;
  assign _02204_ = _02203_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19270" *) _04931_;
  assign _02205_ = _02204_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19271" *) _04932_;
  assign _02206_ = _02205_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19271" *) _03980_;
  assign _02207_ = _02206_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19271" *) or_5189_cse;
  assign _02208_ = _02207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19272" *) cvt_unequal_tmp_20;
  assign _02209_ = mux_2267_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19280" *) _04901_;
  assign _02210_ = _02209_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19280" *) main_stage_v_2;
  assign _02211_ = _02210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19281" *) core_wen;
  assign _02212_ = _02211_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19281" *) or_5189_cse;
  assign _02213_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19290" *) mux_1134_nl;
  assign _02214_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19299" *) FpIntToFloat_17U_5U_10U_is_inf_or_cse;
  assign _02215_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19308" *) mux_2268_nl;
  assign _02216_ = _02215_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19308" *) or_400_cse_1;
  assign _02217_ = _02216_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19308" *) or_4714_cse;
  assign _02218_ = _02217_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *) or_4862_cse;
  assign _02219_ = _02218_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *) core_wen;
  assign _02220_ = _02219_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *) _04901_;
  assign _02221_ = _02220_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19309" *) main_stage_v_2;
  assign _02222_ = _02221_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19310" *) _03931_;
  assign _02223_ = _02222_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19311" *) _04933_;
  assign _02224_ = _02223_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19311" *) _04934_;
  assign _02225_ = _02224_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19312" *) _03980_;
  assign _02226_ = _02225_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19312" *) or_5189_cse;
  assign _02227_ = mux_2269_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19320" *) main_stage_v_2;
  assign _02228_ = _02227_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19320" *) _04901_;
  assign _02229_ = _02228_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19321" *) core_wen;
  assign _02230_ = _02229_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19321" *) or_5189_cse;
  assign _02231_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19329" *) FpIntToFloat_17U_5U_10U_is_inf_or_cse;
  assign _02232_ = _02231_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19330" *) _04935_;
  assign _02233_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19339" *) mux_2270_nl;
  assign _02234_ = _02233_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19339" *) or_4714_cse;
  assign _02235_ = _02234_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19339" *) or_400_cse_1;
  assign _02236_ = _02235_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *) or_4862_cse;
  assign _02237_ = _02236_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *) core_wen;
  assign _02238_ = _02237_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *) _04901_;
  assign _02239_ = _02238_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19340" *) main_stage_v_2;
  assign _02240_ = _02239_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19341" *) _03931_;
  assign _02241_ = _02240_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19342" *) _04936_;
  assign _02242_ = _02241_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19342" *) _04937_;
  assign _02243_ = _02242_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19343" *) _03980_;
  assign _02244_ = _02243_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19343" *) or_5189_cse;
  assign _02245_ = mux_2271_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19351" *) main_stage_v_2;
  assign _02246_ = _02245_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19351" *) _04901_;
  assign _02247_ = _02246_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19352" *) core_wen;
  assign _02248_ = _02247_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19352" *) or_5189_cse;
  assign _02249_ = _02231_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19361" *) _04938_;
  assign _02250_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19370" *) mux_2272_nl;
  assign _02251_ = _02250_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19370" *) or_4714_cse;
  assign _02252_ = _02251_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19370" *) or_400_cse_1;
  assign _02253_ = _02252_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *) or_4862_cse;
  assign _02254_ = _02253_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *) core_wen;
  assign _02255_ = _02254_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *) _04901_;
  assign _02256_ = _02255_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19371" *) main_stage_v_2;
  assign _02257_ = _02256_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19372" *) _03931_;
  assign _02258_ = _02257_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19373" *) _04939_;
  assign _02259_ = _02258_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19373" *) _04940_;
  assign _02260_ = _02259_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19374" *) _03980_;
  assign _02261_ = _02260_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19374" *) or_5189_cse;
  assign _02262_ = mux_2273_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19382" *) main_stage_v_2;
  assign _02263_ = _02262_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19382" *) _04901_;
  assign _02264_ = _02263_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19383" *) core_wen;
  assign _02265_ = _02264_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19383" *) or_5189_cse;
  assign _02266_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19403" *) mux_2274_nl;
  assign _02267_ = _02266_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19403" *) or_4714_cse;
  assign _02268_ = _02267_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19403" *) or_400_cse_1;
  assign _02269_ = _02268_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *) or_4862_cse;
  assign _02270_ = _02269_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *) core_wen;
  assign _02271_ = _02270_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *) _04901_;
  assign _02272_ = _02271_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19404" *) main_stage_v_2;
  assign _02273_ = _02272_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19405" *) _03931_;
  assign _02274_ = _02273_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19406" *) _04941_;
  assign _02275_ = _02274_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19406" *) _04942_;
  assign _02276_ = _02275_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19407" *) _03980_;
  assign _02277_ = _02276_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19407" *) or_5189_cse;
  assign _02278_ = mux_2275_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19415" *) main_stage_v_2;
  assign _02279_ = _02278_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19415" *) _04901_;
  assign _02280_ = _02279_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19416" *) core_wen;
  assign _02281_ = _02280_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19416" *) or_5189_cse;
  assign _02282_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19424" *) _04943_;
  assign _02283_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19432" *) _04944_;
  assign _02284_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19440" *) mux_2276_nl;
  assign _02285_ = _02284_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19440" *) or_4714_cse;
  assign _02286_ = _02285_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19440" *) or_400_cse_1;
  assign _02287_ = _02286_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *) or_4862_cse;
  assign _02288_ = _02287_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *) core_wen;
  assign _02289_ = _02288_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *) _04901_;
  assign _02290_ = _02289_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19441" *) main_stage_v_2;
  assign _02291_ = _02290_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19442" *) _03931_;
  assign _02292_ = _02291_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19443" *) _04945_;
  assign _02293_ = _02292_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19443" *) _04946_;
  assign _02294_ = _02293_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19444" *) _03980_;
  assign _02295_ = _02294_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19444" *) or_5189_cse;
  assign _02296_ = mux_2277_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19452" *) and_dcpl_1319;
  assign _02297_ = _02296_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19452" *) _04901_;
  assign _02298_ = _02297_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19453" *) or_5189_cse;
  assign _02299_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19461" *) core_wen;
  assign _02300_ = _02299_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19461" *) _04947_;
  assign _02301_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19490" *) mux_2278_nl;
  assign _02302_ = _02301_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19490" *) or_4714_cse;
  assign _02303_ = _02302_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19490" *) or_400_cse_1;
  assign _02304_ = _02303_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *) or_4862_cse;
  assign _02305_ = _02304_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *) core_wen;
  assign _02306_ = _02305_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *) _04901_;
  assign _02307_ = _02306_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19491" *) main_stage_v_2;
  assign _02308_ = _02307_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19492" *) _03931_;
  assign _02309_ = _02308_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19493" *) _04948_;
  assign _02310_ = _02309_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19493" *) _04949_;
  assign _02311_ = _02310_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19494" *) _03980_;
  assign _02312_ = _02311_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19494" *) or_5189_cse;
  assign _02313_ = mux_2279_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19502" *) and_dcpl_1319;
  assign _02314_ = _02313_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19502" *) _04901_;
  assign _02315_ = _02314_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19503" *) or_5189_cse;
  assign _02316_ = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19511" *) mux_2280_nl;
  assign _02317_ = _02316_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19511" *) or_4714_cse;
  assign _02318_ = _02317_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19511" *) or_400_cse_1;
  assign _02319_ = _02318_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *) or_4862_cse;
  assign _02320_ = _02319_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *) core_wen;
  assign _02321_ = _02320_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *) _04901_;
  assign _02322_ = _02321_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19512" *) main_stage_v_2;
  assign _02323_ = _02322_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19513" *) _03931_;
  assign _02324_ = _02323_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19514" *) _04950_;
  assign _02325_ = _02324_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19514" *) _04951_;
  assign _02326_ = _02325_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19515" *) _03980_;
  assign _02327_ = _02326_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19515" *) or_5189_cse;
  assign _02328_ = mux_2281_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19523" *) _04901_;
  assign _02329_ = _02328_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19523" *) core_wen;
  assign _02330_ = _02329_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19524" *) main_stage_v_2;
  assign _02331_ = _02330_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19524" *) or_5189_cse;
  assign _02332_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19532" *) mux_1262_nl;
  assign _02333_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19540" *) mux_1266_nl;
  assign and_1179_nl = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19568" *) cfg_mode_eql_1_sva_5;
  assign _02334_ = and_1179_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19568" *) core_wen;
  assign _02335_ = _07811_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19578" *) or_5189_cse;
  assign _02336_ = _02335_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19578" *) core_wen;
  assign _02337_ = _07812_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19586" *) or_5189_cse;
  assign _02338_ = _02337_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19587" *) core_wen;
  assign _02339_ = or_tmp_3032 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19607" *) or_4862_cse;
  assign _02340_ = _02339_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19607" *) or_4714_cse;
  assign _02341_ = _02340_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *) or_5189_cse;
  assign _02342_ = _02341_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *) _03980_;
  assign _02343_ = _02342_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *) main_stage_v_2;
  assign _02344_ = _02343_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19608" *) or_400_cse_1;
  assign _02345_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19609" *) _07813_;
  assign _02346_ = _02345_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19609" *) mux_1429_nl;
  assign _02347_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19663" *) _07814_;
  assign _02348_ = _02347_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19663" *) mux_1472_nl;
  assign _02351_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19805" *) _04955_;
  assign _02352_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19813" *) mux_1534_nl;
  assign _02353_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19821" *) mux_1535_nl;
  assign _02354_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19829" *) mux_1536_nl;
  assign _02355_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19837" *) mux_1537_nl;
  assign _02356_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19845" *) mux_1538_nl;
  assign _02357_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19853" *) mux_1539_nl;
  assign _02358_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19861" *) mux_1540_nl;
  assign _02359_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19869" *) mux_1541_nl;
  assign _02360_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19877" *) mux_1542_nl;
  assign _02361_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19885" *) mux_1543_nl;
  assign _02362_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19893" *) mux_1544_nl;
  assign _02363_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19901" *) mux_1545_nl;
  assign _02364_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19909" *) mux_1546_nl;
  assign _02365_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19917" *) mux_1547_nl;
  assign _02366_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19925" *) mux_1548_nl;
  assign _02367_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19933" *) mux_1549_nl;
  assign _02368_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19941" *) mux_1550_nl;
  assign _02369_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19949" *) mux_1551_nl;
  assign _02370_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19957" *) mux_1552_nl;
  assign _02371_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19965" *) mux_1553_nl;
  assign _02372_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19973" *) mux_1554_nl;
  assign _02373_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19981" *) mux_1555_nl;
  assign _02374_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19989" *) mux_1556_nl;
  assign _02375_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19997" *) mux_1557_nl;
  assign _02376_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20005" *) mux_1558_nl;
  assign _02377_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20013" *) mux_1559_nl;
  assign _02378_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20021" *) mux_1560_nl;
  assign _02379_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20029" *) mux_1561_nl;
  assign _02380_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20037" *) mux_1562_nl;
  assign _02381_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20045" *) mux_1563_nl;
  assign _02382_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20053" *) mux_1564_nl;
  assign _02383_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20061" *) mux_1565_nl;
  assign _02384_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20069" *) _04956_;
  assign _02385_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20078" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl[8];
  assign _02386_ = _02385_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20078" *) _04781_;
  assign _02387_ = _02386_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20078" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8];
  assign _02388_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *) _07815_;
  assign _02389_ = _02388_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *) _04957_;
  assign _02390_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20088" *) _04958_;
  assign _02391_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20097" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _02392_ = _02391_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20097" *) _04783_;
  assign _02393_ = _02392_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20097" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _02394_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20098" *) _07816_;
  assign _02395_ = _02394_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20098" *) _04957_;
  assign _02396_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20107" *) _04959_;
  assign _02397_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20116" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _02398_ = _02397_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20116" *) _04785_;
  assign _02399_ = _02398_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20116" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _02400_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20117" *) _07817_;
  assign _02401_ = _02400_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20117" *) _04957_;
  assign _02402_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20126" *) _04960_;
  assign _02403_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20135" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _02404_ = _02403_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20135" *) _04787_;
  assign _02405_ = _02404_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20135" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _02406_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20136" *) _07818_;
  assign _02407_ = _02406_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20136" *) _04957_;
  assign _02408_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20145" *) _04961_;
  assign _02409_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20154" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _02410_ = _02409_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20154" *) _04789_;
  assign _02411_ = _02410_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20154" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _02412_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20155" *) _07819_;
  assign _02413_ = _02412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20155" *) _04957_;
  assign _02414_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20164" *) _04962_;
  assign _02415_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20173" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _02416_ = _02415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20173" *) _04791_;
  assign _02417_ = _02416_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20173" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _02418_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20174" *) _07820_;
  assign _02419_ = _02418_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20174" *) _04957_;
  assign _02420_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20183" *) mux_1591_nl;
  assign _02421_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20192" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _02422_ = _02421_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20192" *) _04793_;
  assign _02423_ = _02422_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20192" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _02424_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20193" *) _07821_;
  assign _02425_ = _02424_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20193" *) _04957_;
  assign _02426_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20202" *) _04963_;
  assign _02427_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20211" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _02428_ = _02427_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20211" *) _04795_;
  assign _02429_ = _02428_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20211" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _02430_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20212" *) _07822_;
  assign _02431_ = _02430_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20212" *) _04957_;
  assign _02432_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20221" *) _04964_;
  assign _02433_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20230" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _02434_ = _02433_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20230" *) _04797_;
  assign _02435_ = _02434_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20230" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _02436_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20231" *) _07823_;
  assign _02437_ = _02436_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20231" *) _04957_;
  assign _02438_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20240" *) _04965_;
  assign _02439_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20249" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _02440_ = _02439_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20249" *) _04799_;
  assign _02441_ = _02440_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20249" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _02442_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20250" *) _07824_;
  assign _02443_ = _02442_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20250" *) _04957_;
  assign _02444_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20259" *) mux_1605_nl;
  assign _02445_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20268" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _02446_ = _02445_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20268" *) _04801_;
  assign _02447_ = _02446_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20268" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _02448_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20269" *) _07825_;
  assign _02449_ = _02448_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20269" *) _04957_;
  assign _02450_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20278" *) _04966_;
  assign _02451_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20287" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _02452_ = _02451_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20287" *) _04803_;
  assign _02453_ = _02452_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20287" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _02454_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20288" *) _07826_;
  assign _02455_ = _02454_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20288" *) _04957_;
  assign _02456_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20297" *) _04967_;
  assign _02457_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20306" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _02458_ = _02457_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20306" *) _04805_;
  assign _02459_ = _02458_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20306" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _02460_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20307" *) _07827_;
  assign _02461_ = _02460_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20307" *) _04957_;
  assign _02462_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20316" *) _04968_;
  assign _02463_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20325" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _02464_ = _02463_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20325" *) _04807_;
  assign _02465_ = _02464_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20325" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _02466_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20326" *) _07828_;
  assign _02467_ = _02466_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20326" *) _04957_;
  assign _02468_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20335" *) _04969_;
  assign _02469_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20344" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _02470_ = _02469_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20344" *) _04809_;
  assign _02471_ = _02470_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20344" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _02472_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20345" *) _07829_;
  assign _02473_ = _02472_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20345" *) _04957_;
  assign _02474_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20354" *) _04970_;
  assign _02475_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20363" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8];
  assign _02476_ = _02475_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20363" *) _04811_;
  assign _02477_ = _02476_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20363" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8];
  assign _02478_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20364" *) _07830_;
  assign _02479_ = _02478_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20364" *) _04957_;
  assign _02480_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20375" *) _07832_;
  assign _02481_ = _02480_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20375" *) mux_tmp_161;
  assign _02482_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20387" *) _07834_;
  assign _02483_ = _02482_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20387" *) mux_tmp_161;
  assign _02484_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20399" *) _07836_;
  assign _02485_ = _02484_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20399" *) mux_tmp_161;
  assign _02486_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20411" *) _07838_;
  assign _02487_ = _02486_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20411" *) mux_tmp_161;
  assign _02488_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20423" *) _07840_;
  assign _02489_ = _02488_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20423" *) mux_tmp_161;
  assign _02490_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20435" *) _07842_;
  assign _02491_ = _02490_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20435" *) mux_tmp_161;
  assign _02492_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20447" *) _07844_;
  assign _02493_ = _02492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20447" *) mux_tmp_161;
  assign _02494_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20459" *) _07846_;
  assign _02495_ = _02494_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20459" *) mux_tmp_161;
  assign _02496_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20471" *) _07848_;
  assign _02497_ = _02496_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20471" *) mux_tmp_161;
  assign _02498_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20483" *) _07850_;
  assign _02499_ = _02498_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20483" *) mux_tmp_161;
  assign _02500_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20495" *) _07852_;
  assign _02501_ = _02500_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20495" *) mux_tmp_161;
  assign _02502_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20506" *) _07854_;
  assign _02503_ = _02502_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20507" *) mux_tmp_161;
  assign _02504_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20518" *) _07856_;
  assign _02505_ = _02504_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20519" *) mux_tmp_161;
  assign _02506_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20530" *) _07858_;
  assign _02507_ = _02506_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20531" *) mux_tmp_161;
  assign _02508_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20542" *) _07860_;
  assign _02509_ = _02508_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20543" *) mux_tmp_161;
  assign _02510_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20554" *) _07862_;
  assign _02511_ = _02510_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20555" *) mux_tmp_161;
  assign _02512_ = IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20581" *) _04971_;
  assign _02513_ = IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20583" *) _04972_;
  assign _02514_ = IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20585" *) _04973_;
  assign _02515_ = IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20587" *) _04974_;
  assign _02516_ = IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20589" *) _04975_;
  assign _02517_ = IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20591" *) _04976_;
  assign _02518_ = IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20593" *) _04977_;
  assign _02519_ = IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20595" *) _04978_;
  assign _02520_ = IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20597" *) _04979_;
  assign _02521_ = IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20599" *) _04980_;
  assign _02522_ = IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20601" *) _04981_;
  assign _02523_ = IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20603" *) _04982_;
  assign _02524_ = IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20605" *) _04983_;
  assign _02525_ = IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20607" *) _04984_;
  assign _02526_ = IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20609" *) _04985_;
  assign _02527_ = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20616" *) mux_1627_nl;
  assign _02528_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20625" *) mux_1640_nl;
  assign _02529_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20635" *) mux_1649_nl;
  assign _02530_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20646" *) mux_1660_nl;
  assign _02531_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20656" *) mux_1663_nl;
  assign _02532_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20666" *) mux_1674_nl;
  assign _02533_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20676" *) mux_1685_nl;
  assign _02534_ = _01449_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20701" *) mux_320_cse;
  assign _02535_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20726" *) IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_15_cse;
  assign _02536_ = _02535_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20726" *) mux_449_nl;
  assign _02537_ = _01446_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20737" *) mux_454_nl;
  assign _02538_ = _02535_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20762" *) mux_272_cse;
  assign _02539_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20787" *) IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_8_cse;
  assign _02540_ = _02539_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20787" *) mux_770_nl;
  assign _02541_ = _02539_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20798" *) mux_789_nl;
  assign _02542_ = _01446_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20809" *) mux_799_nl;
  assign _02543_ = or_dcpl_386 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20819" *) or_4862_cse;
  assign _02544_ = _02543_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20819" *) and_dcpl_401;
  assign _02545_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20820" *) _07878_;
  assign _02546_ = _02545_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20820" *) mux_803_nl;
  assign _02547_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *) _04986_;
  assign _02548_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *) _04987_;
  assign _02549_ = _02548_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *) mux_tmp_245;
  assign _02550_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *) _04988_;
  assign _02551_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *) _04989_;
  assign _02552_ = _02551_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *) mux_1687_nl;
  assign _02553_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *) _04990_;
  assign _02554_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *) _04991_;
  assign _02555_ = _02554_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *) mux_1689_nl;
  assign _02556_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *) _04992_;
  assign _02557_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *) _04993_;
  assign _02558_ = _02557_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *) mux_1692_nl;
  assign _02559_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20904" *) _04994_;
  assign _02560_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20914" *) _04995_;
  assign _02561_ = _02560_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20914" *) mux_1694_nl;
  assign _02562_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *) _04996_;
  assign _02563_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *) _04997_;
  assign _02564_ = _02563_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *) mux_1697_nl;
  assign _02565_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *) _04998_;
  assign _02566_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *) _04999_;
  assign _02567_ = _02566_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *) mux_1700_nl;
  assign _02568_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *) _05000_;
  assign _02569_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *) _05001_;
  assign _02570_ = _02569_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *) mux_1704_nl;
  assign _02571_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20979" *) _05002_;
  assign _02572_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20989" *) _05003_;
  assign _02573_ = _02572_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20989" *) mux_1707_nl;
  assign _02574_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *) _05004_;
  assign _02575_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *) _05005_;
  assign _02576_ = _02575_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21007" *) mux_1711_nl;
  assign _02577_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *) _05006_;
  assign _02578_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *) _05007_;
  assign _02579_ = _02578_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *) mux_1715_nl;
  assign _02580_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *) _05008_;
  assign _02581_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *) _05009_;
  assign _02582_ = _02581_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21045" *) mux_tmp_585;
  assign _02583_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21055" *) _05010_;
  assign _02584_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21065" *) _05011_;
  assign _02585_ = _02584_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21065" *) mux_1720_nl;
  assign _02586_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21075" *) _05012_;
  assign _02587_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *) _05013_;
  assign _02588_ = _02587_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *) mux_1727_nl;
  assign _02589_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21094" *) _05014_;
  assign _02590_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *) _05015_;
  assign _02591_ = _02590_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *) mux_1734_nl;
  assign _02592_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *) _05016_;
  assign _02593_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *) _05017_;
  assign _02594_ = _02593_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21122" *) mux_1743_nl;
  assign _02595_ = _01459_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21152" *) _05018_;
  assign _02596_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *) _05019_;
  assign _02597_ = _02596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *) _05020_;
  assign _02598_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21180" *) _05021_;
  assign _02599_ = _02598_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21180" *) mux_121_nl;
  assign _02601_ = _02600_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *) _05023_;
  assign _02602_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21206" *) FpIntToFloat_17U_5U_10U_if_nor_6_cse;
  assign _02603_ = _02602_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21207" *) mux_131_nl;
  assign _02604_ = _02602_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21226" *) mux_134_cse;
  assign _02605_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21234" *) nor_1992_nl;
  assign _02606_ = _02605_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21234" *) mux_143_nl;
  assign _02607_ = _02602_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21243" *) mux_150_nl;
  assign _02608_ = _01460_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21252" *) mux_153_nl;
  assign _02609_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *) _05024_;
  assign _02610_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *) _05025_;
  assign _02611_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *) _05026_;
  assign _02612_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *) _05027_;
  assign _02613_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *) _05028_;
  assign _02614_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *) _05029_;
  assign _02615_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *) _05030_;
  assign _02616_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *) _05031_;
  assign _02617_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *) _05032_;
  assign _02618_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *) _05033_;
  assign _02619_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *) _05034_;
  assign _02620_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *) _05035_;
  assign _02621_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *) _05036_;
  assign _02622_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *) _05037_;
  assign _02623_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *) _05038_;
  assign _02624_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *) _05039_;
  assign cvt_and_261_nl = _01622_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21417" *) _05040_;
  assign cvt_and_262_nl = FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21418" *) cvt_asn_323;
  assign cvt_and_257_nl = _01626_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21420" *) _05041_;
  assign cvt_and_258_nl = FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21421" *) cvt_asn_323;
  assign cvt_and_253_nl = _01630_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21423" *) _05042_;
  assign cvt_and_254_nl = FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21424" *) cvt_asn_323;
  assign cvt_and_245_nl = _01638_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21426" *) _05043_;
  assign cvt_and_246_nl = FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21427" *) cvt_asn_323;
  assign _02625_ = reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21429" *) _04700_;
  assign _02626_ = reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21431" *) _04702_;
  assign _02627_ = reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21433" *) _04704_;
  assign _02628_ = reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21435" *) _04706_;
  assign _02629_ = reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21437" *) _04708_;
  assign _02630_ = reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21439" *) _04710_;
  assign _02631_ = reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21441" *) _04712_;
  assign _02632_ = reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21443" *) _04714_;
  assign _02633_ = reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21445" *) _04716_;
  assign _02634_ = reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21447" *) _04718_;
  assign _02635_ = reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21449" *) _04720_;
  assign _02636_ = reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21451" *) _04722_;
  assign _02637_ = reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21453" *) _04724_;
  assign _02638_ = reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21455" *) _04726_;
  assign _02639_ = reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21457" *) _04728_;
  assign _02640_ = reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21459" *) _04730_;
  assign cvt_and_259_nl = _01624_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21462" *) _05044_;
  assign cvt_and_260_nl = FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21463" *) cvt_asn_329;
  assign and_3148_nl = cvt_asn_333 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21464" *) _05044_;
  assign and_3140_nl = cvt_or_6_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21467" *) _05045_;
  assign cvt_and_255_nl = _01628_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21469" *) _05045_;
  assign cvt_and_256_nl = FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21470" *) cvt_asn_335;
  assign cvt_and_251_nl = _01632_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21474" *) _05046_;
  assign cvt_and_252_nl = FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21475" *) cvt_asn_353;
  assign and_3136_nl = cvt_asn_357 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21476" *) _05046_;
  assign cvt_and_249_nl = _01634_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21480" *) _05047_;
  assign cvt_and_250_nl = FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21481" *) cvt_asn_365;
  assign and_3133_nl = cvt_asn_369 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21482" *) _05047_;
  assign and_3128_nl = cvt_or_14_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21485" *) _05048_;
  assign cvt_and_247_nl = _01636_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21487" *) _05048_;
  assign cvt_and_248_nl = FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21488" *) cvt_asn_377;
  assign and_3130_nl = cvt_asn_381 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21489" *) _05048_;
  assign cvt_and_243_nl = _01640_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21493" *) _05049_;
  assign cvt_and_244_nl = FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21494" *) cvt_asn_371;
  assign and_3124_nl = cvt_asn_399 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21495" *) _05049_;
  assign cvt_and_241_nl = _01642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21499" *) _05050_;
  assign cvt_and_242_nl = FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21500" *) cvt_asn_389;
  assign and_3121_nl = cvt_asn_393 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21501" *) _05050_;
  assign and_3116_nl = cvt_or_22_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21504" *) _05051_;
  assign cvt_and_239_nl = _01644_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21506" *) _05051_;
  assign cvt_and_240_nl = FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21507" *) cvt_asn_383;
  assign and_3118_nl = cvt_asn_387 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21508" *) _05051_;
  assign cvt_and_237_nl = _01646_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21512" *) _05052_;
  assign cvt_and_238_nl = FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21513" *) cvt_asn_371;
  assign and_3115_nl = cvt_asn_375 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21514" *) _05052_;
  assign and_3110_nl = cvt_or_26_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21517" *) _05053_;
  assign cvt_and_235_nl = _01648_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21519" *) _05053_;
  assign cvt_and_236_nl = FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21520" *) cvt_asn_359;
  assign and_3112_nl = cvt_asn_363 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21521" *) _05053_;
  assign and_3104_nl = cvt_or_30_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21522" *) _05054_;
  assign cvt_and_231_nl = _01652_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21524" *) _05054_;
  assign cvt_and_232_nl = FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21525" *) cvt_asn_341;
  assign and_3105_nl = cvt_asn_345 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21526" *) _05054_;
  assign cvt_and_233_nl = _01650_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21528" *) _05055_;
  assign cvt_and_234_nl = FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21529" *) cvt_asn_347;
  assign and_3109_nl = cvt_asn_351 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21530" *) _05055_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_nl = FpFloatToInt_16U_5U_10U_mux_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21541" *) _04718_;
  assign _02641_ = cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21547" *) _05056_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_1_nl = FpFloatToInt_16U_5U_10U_mux_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21568" *) _04700_;
  assign _02642_ = IntShiftRightSat_49U_6U_17U_o_0_2_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21574" *) _05057_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_2_nl = FpFloatToInt_16U_5U_10U_mux_18_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21594" *) _04702_;
  assign _02643_ = IntShiftRightSat_49U_6U_17U_o_0_3_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21600" *) _05058_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_3_nl = FpFloatToInt_16U_5U_10U_mux_25_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21621" *) _04704_;
  assign _02644_ = IntShiftRightSat_49U_6U_17U_o_0_4_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21627" *) _05059_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_4_nl = FpFloatToInt_16U_5U_10U_mux_32_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21648" *) _04706_;
  assign _02645_ = IntShiftRightSat_49U_6U_17U_o_0_5_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21654" *) _05060_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_5_nl = FpFloatToInt_16U_5U_10U_mux_39_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21675" *) _04708_;
  assign _02646_ = IntShiftRightSat_49U_6U_17U_o_0_6_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21681" *) _05061_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_6_nl = FpFloatToInt_16U_5U_10U_mux_46_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21702" *) _04710_;
  assign _02647_ = IntShiftRightSat_49U_6U_17U_o_0_7_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21708" *) _05062_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_7_nl = FpFloatToInt_16U_5U_10U_mux_53_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21729" *) _04712_;
  assign _02648_ = IntShiftRightSat_49U_6U_17U_o_0_8_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21735" *) _05063_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_8_nl = FpFloatToInt_16U_5U_10U_mux_60_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21756" *) _04714_;
  assign _02649_ = IntShiftRightSat_49U_6U_17U_o_0_9_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21762" *) _05064_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_9_nl = FpFloatToInt_16U_5U_10U_mux_67_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21783" *) _04720_;
  assign _02650_ = cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21789" *) _05065_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_10_nl = FpFloatToInt_16U_5U_10U_mux_74_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21810" *) _04722_;
  assign _02651_ = IntShiftRightSat_49U_6U_17U_o_0_11_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21816" *) _05066_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_11_nl = FpFloatToInt_16U_5U_10U_mux_81_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21837" *) _04724_;
  assign _02652_ = IntShiftRightSat_49U_6U_17U_o_0_12_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21843" *) _05067_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_12_nl = FpFloatToInt_16U_5U_10U_mux_88_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21864" *) _04726_;
  assign _02653_ = IntShiftRightSat_49U_6U_17U_o_0_13_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21870" *) _05068_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_13_nl = FpFloatToInt_16U_5U_10U_mux_95_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21891" *) _04728_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_14_nl = FpFloatToInt_16U_5U_10U_mux_102_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21914" *) _04730_;
  assign _02654_ = IntShiftRightSat_49U_6U_17U_o_0_15_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21920" *) _05069_;
  assign _02655_ = IntShiftRightSat_49U_6U_17U_o_0_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21935" *) _05070_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_15_nl = FpFloatToInt_16U_5U_10U_mux_109_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21947" *) _04716_;
  assign _02656_ = cvt_1_FpMantRNE_24U_11U_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21969" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8];
  assign _02657_ = _02656_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21969" *) _03950_;
  assign and_98_nl = chn_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21977" *) mux_2_nl;
  assign _02658_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2;
  assign _02659_ = _02658_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2;
  assign _02660_ = _05075_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2;
  assign and_2240_nl = _08073_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21982" *) main_stage_v_1;
  assign and_2242_nl = _08074_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21986" *) main_stage_v_1;
  assign _02661_ = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22096" *) main_stage_v_1;
  assign _02662_ = _02661_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22096" *) and_dcpl_3;
  assign _02663_ = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22125" *) main_stage_v_1;
  assign _02664_ = _02663_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22125" *) and_dcpl_3;
  assign _02665_ = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22147" *) main_stage_v_1;
  assign _02666_ = _02665_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22147" *) and_dcpl_3;
  assign _02667_ = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22224" *) main_stage_v_1;
  assign _02668_ = _02667_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22224" *) and_dcpl_3;
  assign _02669_ = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22301" *) main_stage_v_1;
  assign _02670_ = _02669_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22301" *) and_dcpl_3;
  assign and_132_nl = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22477" *) mux_155_nl;
  assign _02671_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22538" *) cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp;
  assign and_143_nl = _02671_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22538" *) or_4550_cse;
  assign _02672_ = and_dcpl_114 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22541" *) cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp;
  assign and_145_nl = _02672_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22541" *) or_4550_cse;
  assign and_2857_nl = mux_tmp_239 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22546" *) and_dcpl_444;
  assign _02673_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22556" *) cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  assign and_147_nl = _02673_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22556" *) and_tmp_12;
  assign and_2234_nl = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22560" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign and_2233_nl = IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22565" *) mux_tmp_263;
  assign _02674_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22573" *) cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  assign and_156_nl = _02674_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22573" *) and_tmp_12;
  assign _02675_ = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22575" *) cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  assign and_160_nl = _02675_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22575" *) and_tmp_50;
  assign and_161_nl = _08304_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22580" *) mux_tmp_263;
  assign _02676_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22589" *) cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  assign and_164_nl = _02676_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22589" *) mux_tmp_117;
  assign and_166_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22592" *) mux_290_nl;
  assign and_168_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22606" *) mux_tmp_321;
  assign _02677_ = cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22610" *) main_stage_v_2;
  assign and_171_nl = _02677_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22610" *) mux_1126_cse;
  assign and_172_nl = _08310_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22616" *) mux_tmp_263;
  assign and_2265_nl = _08311_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22621" *) or_tmp_3768;
  assign _02678_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22629" *) cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  assign and_173_nl = _02678_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22629" *) mux_344_cse;
  assign _02679_ = IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22631" *) main_stage_v_2;
  assign and_2229_nl = _02679_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22631" *) mux_382_cse;
  assign _02680_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22647" *) cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  assign and_179_nl = _02680_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22647" *) mux_344_cse;
  assign _02681_ = or_4536_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22648" *) main_stage_v_2;
  assign and_180_nl = _02681_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22648" *) mux_382_cse;
  assign _02682_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22663" *) cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  assign and_182_nl = _02682_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22663" *) mux_344_cse;
  assign _02683_ = or_4535_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22664" *) main_stage_v_2;
  assign and_183_nl = _02683_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22664" *) mux_417_cse;
  assign and_185_nl = or_4535_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22675" *) mux_tmp_441;
  assign and_2856_nl = and_tmp_93 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22685" *) or_5189_cse;
  assign and_194_nl = cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22690" *) mux_tmp_263;
  assign _02684_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22697" *) cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  assign and_195_nl = _02684_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22697" *) mux_474_cse;
  assign _02685_ = IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22699" *) main_stage_v_2;
  assign and_2221_nl = _02685_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22699" *) mux_382_cse;
  assign _02686_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22715" *) cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  assign and_199_nl = _02686_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22715" *) mux_474_cse;
  assign _02687_ = IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22717" *) main_stage_v_2;
  assign and_2217_nl = _02687_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22717" *) mux_382_cse;
  assign _02688_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22733" *) cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  assign and_203_nl = _02688_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22733" *) mux_474_cse;
  assign and_2213_nl = IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22734" *) mux_417_cse;
  assign and_205_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22736" *) mux_555_nl;
  assign _02689_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22752" *) cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  assign and_210_nl = _02689_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22752" *) mux_474_cse;
  assign and_212_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22755" *) mux_593_nl;
  assign _02690_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22757" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign _02691_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22773" *) cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  assign and_213_nl = _02691_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22773" *) mux_474_cse;
  assign and_2203_nl = IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22774" *) mux_417_cse;
  assign and_215_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22776" *) mux_629_nl;
  assign _02692_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22792" *) cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  assign and_216_nl = _02692_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22792" *) mux_474_cse;
  assign and_2201_nl = IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22793" *) mux_417_cse;
  assign and_218_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22795" *) mux_670_nl;
  assign _02693_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22797" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign _02694_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22817" *) cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp;
  assign and_219_nl = _02694_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22817" *) mux_344_cse;
  assign and_2196_nl = IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22818" *) mux_417_cse;
  assign and_221_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22820" *) mux_714_nl;
  assign _02695_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22822" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp;
  assign and_136_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22843" *) or_tmp_389;
  assign _02696_ = _08350_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22887" *) or_1159_cse;
  assign and_227_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22899" *) _08355_;
  assign _02697_ = cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22901" *) _05125_;
  assign and_228_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22903" *) mux_814_nl;
  assign and_229_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22909" *) _08359_;
  assign _02698_ = cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22911" *) _05125_;
  assign and_230_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22913" *) mux_821_nl;
  assign _02699_ = or_1202_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *) _05130_;
  assign and_2191_nl = IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22920" *) cvt_unequal_tmp_20;
  assign and_2357_nl = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22929" *) _08368_;
  assign and_233_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22935" *) _08372_;
  assign _02700_ = cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22937" *) _05125_;
  assign and_234_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22939" *) mux_832_nl;
  assign and_235_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22951" *) _08376_;
  assign _02701_ = cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22953" *) _05125_;
  assign and_236_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22955" *) mux_836_nl;
  assign _02702_ = _05135_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22958" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c;
  assign FpFloatToInt_16U_5U_10U_and_37_nl = _02702_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22958" *) and_dcpl_408;
  assign _02703_ = chn_idata_data_sva_2_143_127_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22960" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c;
  assign FpFloatToInt_16U_5U_10U_and_38_nl = _02703_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22960" *) and_dcpl_408;
  assign _02704_ = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22962" *) _05136_;
  assign FpFloatToInt_16U_5U_10U_and_7_nl = _02704_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22962" *) and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_o_int_and_28_nl = IsNaN_5U_10U_land_4_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22964" *) and_dcpl_408;
  assign and_237_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22969" *) _08380_;
  assign _02705_ = cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22971" *) _05125_;
  assign and_238_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22973" *) mux_840_nl;
  assign _02706_ = _08390_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22986" *) or_1159_cse;
  assign and_240_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22998" *) _08395_;
  assign _02707_ = cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23000" *) _05125_;
  assign and_241_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23002" *) mux_852_nl;
  assign and_242_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23020" *) _08406_;
  assign _02708_ = cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23022" *) _05125_;
  assign and_243_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23024" *) mux_862_nl;
  assign and_244_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23030" *) _08410_;
  assign _02709_ = cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23032" *) _05125_;
  assign and_245_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23034" *) mux_866_nl;
  assign _02710_ = _08420_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23047" *) or_1159_cse;
  assign and_247_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23059" *) _08425_;
  assign _02711_ = cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23061" *) _05125_;
  assign and_248_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23063" *) mux_878_nl;
  assign _02712_ = _08435_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23076" *) or_1159_cse;
  assign and_250_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23088" *) _08440_;
  assign _02713_ = cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23090" *) _05125_;
  assign and_251_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23092" *) mux_890_nl;
  assign _02714_ = nor_63_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23094" *) nor_1048_cse;
  assign _02715_ = _05159_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *) nor_1048_cse;
  assign _02716_ = _05163_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *) nor_1048_cse;
  assign and_2190_nl = cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23102" *) cvt_unequal_tmp_20;
  assign and_2189_nl = nor_1666_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23124" *) mux_906_nl;
  assign and_252_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23138" *) _08462_;
  assign _02717_ = cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23140" *) _05125_;
  assign and_253_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23142" *) mux_912_nl;
  assign _02718_ = _08474_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23160" *) mux_1832_nl;
  assign and_255_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23168" *) _08479_;
  assign _02719_ = cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23170" *) _05125_;
  assign and_256_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23172" *) mux_924_nl;
  assign and_257_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23178" *) _08483_;
  assign _02720_ = cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23180" *) _05125_;
  assign and_258_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23182" *) mux_928_nl;
  assign and_259_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23188" *) _08487_;
  assign _02721_ = cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23190" *) _05125_;
  assign and_260_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23192" *) mux_932_nl;
  assign and_261_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23198" *) _08491_;
  assign _02722_ = cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23200" *) _05125_;
  assign and_262_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23202" *) mux_936_nl;
  assign and_2811_nl = _05198_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23361" *) or_1202_cse;
  assign _02723_ = _04898_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23364" *) _03981_;
  assign _02724_ = _05200_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23380" *) FpMantRNE_17U_11U_else_mux_3_nl;
  assign _02725_ = _05201_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23381" *) FpIntToFloat_17U_5U_10U_else_mux_4_nl;
  assign and_2809_nl = _05203_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23388" *) or_1596_cse;
  assign _02726_ = _05200_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23393" *) _03982_;
  assign _02727_ = or_1596_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *) _05204_;
  assign and_2807_nl = _05206_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23407" *) or_1625_cse;
  assign _02728_ = _04907_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23412" *) _03983_;
  assign _02729_ = or_1625_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *) _05207_;
  assign and_2805_nl = _05209_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23421" *) or_1659_cse_1;
  assign _02730_ = _04287_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23426" *) _03984_;
  assign _02731_ = or_1659_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *) _05210_;
  assign and_2803_nl = _05212_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23430" *) or_1693_cse;
  assign _02732_ = _04910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23435" *) _03985_;
  assign _02733_ = or_1693_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *) _05213_;
  assign and_2801_nl = _05215_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23448" *) or_1720_cse_1;
  assign _02734_ = _04289_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23453" *) _03986_;
  assign _02735_ = or_1720_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *) _05216_;
  assign and_2799_nl = _05218_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23460" *) or_1752_cse_1;
  assign _02736_ = _04291_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23465" *) _03987_;
  assign _02737_ = or_1752_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *) _05219_;
  assign and_2797_nl = _05221_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23476" *) or_1789_cse_1;
  assign _02738_ = _04293_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23481" *) _03988_;
  assign _02739_ = or_1789_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *) _05222_;
  assign and_2795_nl = _05224_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23494" *) or_1829_cse;
  assign _02740_ = _04928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23499" *) _03989_;
  assign _02741_ = or_1829_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *) _05225_;
  assign and_2793_nl = _05227_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23505" *) or_1851_cse_1;
  assign _02742_ = or_400_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23509" *) or_1851_cse_1;
  assign _02743_ = _04295_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23510" *) _03990_;
  assign _02744_ = _02742_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *) _05228_;
  assign and_2791_nl = _05230_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23517" *) or_1892_cse_1;
  assign _02745_ = _04297_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23522" *) _03991_;
  assign _02746_ = or_1892_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *) _05231_;
  assign and_2789_nl = or_400_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *) _05233_;
  assign and_3372_nl = mux_1142_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23525" *) _04947_;
  assign _02747_ = cfg_proc_precision_1_sva_st_108[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23530" *) mux_tmp_987;
  assign and_2788_nl = _05235_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23538" *) or_1925_cse_1;
  assign _02748_ = _04299_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23543" *) _03992_;
  assign _02749_ = or_1925_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *) _05236_;
  assign and_3373_nl = or_400_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *) _05238_;
  assign and_2786_nl = _05239_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23547" *) or_5038_cse;
  assign _02750_ = _04301_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23550" *) _03993_;
  assign _02751_ = or_5038_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23551" *) or_400_cse_1;
  assign _02752_ = _02751_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *) _05240_;
  assign _02753_ = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23556" *) _05242_;
  assign _02754_ = cvt_else_equal_tmp_46 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23557" *) main_stage_v_3;
  assign _02755_ = _02754_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23557" *) mux_tmp_1197;
  assign _02756_ = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23562" *) _05243_;
  assign _02757_ = cvt_else_equal_tmp_45 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23563" *) main_stage_v_3;
  assign _02758_ = _02757_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23563" *) mux_tmp_1197;
  assign and_2784_nl = _05244_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23568" *) or_5053_cse;
  assign _02759_ = _04303_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23571" *) _03994_;
  assign _02760_ = or_5053_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23572" *) or_400_cse_1;
  assign _02761_ = _02760_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *) _05245_;
  assign and_2782_nl = _05247_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23577" *) or_5069_cse;
  assign _02762_ = _04305_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23580" *) _03995_;
  assign _02763_ = or_5069_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23581" *) or_400_cse_1;
  assign _02764_ = _02763_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *) _05248_;
  assign and_2780_nl = _05250_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23586" *) or_5086_cse;
  assign _02765_ = _04307_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23589" *) _03996_;
  assign _02766_ = or_5086_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *) _05251_;
  assign and_223_nl = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23594" *) mux_417_cse;
  assign _02767_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23620" *) mux_1466_cse;
  assign _02768_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23625" *) mux_1470_nl;
  assign _02769_ = cvt_1_FpMantRNE_24U_11U_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23644" *) _03950_;
  assign _02770_ = cvt_2_FpMantRNE_24U_11U_else_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23667" *) _03949_;
  assign _02771_ = cvt_3_FpMantRNE_24U_11U_else_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23690" *) _03948_;
  assign _02772_ = cvt_4_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23713" *) _03947_;
  assign _02773_ = cvt_5_FpMantRNE_24U_11U_else_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23736" *) _03946_;
  assign _02774_ = or_tmp_2466 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23738" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _02775_ = _02774_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23738" *) _04803_;
  assign _02776_ = _02775_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _02777_ = _02776_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *) _03865_;
  assign _02778_ = _02777_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *) chn_in_rsci_bawt;
  assign _02779_ = cvt_6_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23759" *) _03945_;
  assign _02780_ = cvt_7_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23782" *) _03944_;
  assign _02781_ = cvt_8_FpMantRNE_24U_11U_else_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23805" *) _03943_;
  assign _02782_ = cvt_9_FpMantRNE_24U_11U_else_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23828" *) _03942_;
  assign _02783_ = cvt_10_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23851" *) _03941_;
  assign _02784_ = cvt_11_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23874" *) _03940_;
  assign _02785_ = cvt_12_FpMantRNE_24U_11U_else_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23897" *) _03939_;
  assign _02786_ = cvt_13_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23920" *) _03938_;
  assign _02787_ = cvt_14_FpMantRNE_24U_11U_else_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23943" *) _03937_;
  assign _02788_ = cvt_15_FpMantRNE_24U_11U_else_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23966" *) _03936_;
  assign _02789_ = cvt_16_FpMantRNE_24U_11U_else_and_4_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23989" *) _03935_;
  assign _02790_ = cvt_10_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24031" *) _03865_;
  assign and_2243_nl = _02790_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24031" *) chn_in_rsci_bawt;
  assign _02791_ = cvt_10_FpMantRNE_24U_11U_else_and_2_svs & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24033" *) _03865_;
  assign and_2162_nl = _02791_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24033" *) chn_in_rsci_bawt;
  assign _02792_ = cfg_proc_precision_1_sva_st_64[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *) cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign _02793_ = cvt_6_FpMantRNE_24U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24056" *) _03865_;
  assign and_nl = _02793_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24056" *) chn_in_rsci_bawt;
  assign _02794_ = cvt_6_FpMantRNE_24U_11U_else_and_2_svs & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24058" *) _03865_;
  assign and_2161_nl = _02794_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24058" *) chn_in_rsci_bawt;
  assign _02795_ = cfg_proc_precision_1_sva_st_64[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24063" *) cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign and_2160_nl = cfg_mode_eql_1_sva_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24090" *) main_stage_v_2;
  assign _02796_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24099" *) _03997_;
  assign _02797_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24110" *) _03998_;
  assign _02798_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24119" *) _03999_;
  assign _02799_ = cfg_proc_precision_1_sva_st_101[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24132" *) mux_tmp_455;
  assign _02800_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24229" *) and_tmp_16;
  assign _02801_ = cvt_10_IntSaturation_17U_8U_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02802_ = cvt_2_IntSaturation_17U_8U_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02803_ = cvt_3_IntSaturation_17U_8U_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02804_ = cvt_4_IntSaturation_17U_8U_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02805_ = cvt_5_IntSaturation_17U_8U_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02806_ = cvt_6_IntSaturation_17U_8U_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02807_ = cvt_1_IntSaturation_17U_8U_if_acc_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02808_ = cvt_7_IntSaturation_17U_8U_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02809_ = cvt_16_IntSaturation_17U_8U_if_acc_4_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02810_ = cvt_8_IntSaturation_17U_8U_if_acc_3_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02811_ = cvt_15_IntSaturation_17U_8U_if_acc_3_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02812_ = cvt_9_IntSaturation_17U_8U_if_acc_1_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02813_ = cvt_13_IntSaturation_17U_8U_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02814_ = cvt_11_IntSaturation_17U_8U_if_acc_2_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02815_ = cvt_12_IntSaturation_17U_8U_if_acc_3_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_411;
  assign _02816_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02817_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02818_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02819_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02820_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02821_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02822_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02823_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02824_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02825_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02826_ = IntShiftRightSat_49U_6U_17U_o_0_1_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02827_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02828_ = IntShiftRightSat_49U_6U_17U_o_0_10_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02829_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02830_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02831_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) and_dcpl_420;
  assign _02832_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_13_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_mux_59_nl;
  assign _02833_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02834_ = IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02835_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_1_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_4_mx1;
  assign _02836_ = IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_4_mx1;
  assign _02837_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02838_ = IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02839_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_10_mx0;
  assign _02840_ = IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_10_mx0;
  assign _02841_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02842_ = IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02843_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_16_mx1;
  assign _02844_ = IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_16_mx1;
  assign _02845_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_19_mx0;
  assign _02846_ = IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_19_mx0;
  assign _02847_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_22_mx1;
  assign _02848_ = IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_22_mx1;
  assign _02849_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_8_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02850_ = IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_1;
  assign _02851_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_9_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_28_mx1;
  assign _02852_ = IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_28_mx1;
  assign _02853_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_10_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_31_mx0;
  assign _02854_ = IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_31_mx0;
  assign _02855_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_34_mx1;
  assign _02856_ = IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_34_mx1;
  assign _02857_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_12_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_37_mx0;
  assign _02858_ = IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_37_mx0;
  assign _02859_ = IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_40_mx1;
  assign _02860_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_14_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_43_mx0;
  assign _02861_ = IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_43_mx0;
  assign _02862_ = IntSaturation_17U_8U_IntSaturation_17U_8U_or_15_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_40_mx1;
  assign _02863_ = IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24251" *) cvt_else_equal_tmp_40_mx1;
  assign _02864_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02865_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02866_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02867_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02868_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02869_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02870_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02871_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02872_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02873_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02874_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02875_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02876_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02877_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02878_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_dcpl_409;
  assign _02879_ = FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_900_rgt;
  assign _02880_ = FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  assign _02881_ = FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  assign _02882_ = FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _02883_ = FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_956_rgt;
  assign _02884_ = FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1;
  assign _02885_ = FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _02886_ = FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_986_rgt;
  assign _02887_ = FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_989_rgt;
  assign _02888_ = FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  assign _02889_ = FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) and_1011_rgt;
  assign _02890_ = FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _02891_ = FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  assign _02892_ = FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  assign _02893_ = FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _02894_ = FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _02895_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_mux_62_nl;
  assign _02896_ = cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02897_ = reg_chn_idata_data_sva_3_15_0_1_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02898_ = IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_3_mx0;
  assign _02899_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_3_mx0;
  assign _02900_ = cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02901_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02902_ = cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_9_mx1;
  assign _02903_ = FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[14] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_9_mx1;
  assign _02904_ = cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02905_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02906_ = cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_15_mx0;
  assign _02907_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_15_mx0;
  assign _02908_ = cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_18_mx0;
  assign _02909_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_18_mx0;
  assign _02910_ = cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_21_mx1;
  assign _02911_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_21_mx1;
  assign _02912_ = cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02913_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp;
  assign _02914_ = cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_27_mx0;
  assign _02915_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_27_mx0;
  assign _02916_ = cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_30_mx0;
  assign _02917_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_30_mx0;
  assign _02918_ = cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_33_mx1;
  assign _02919_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_33_mx1;
  assign _02920_ = cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_36_mx0;
  assign _02921_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_36_mx0;
  assign _02922_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_39_mx1;
  assign _02923_ = cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_42_mx0;
  assign _02924_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_42_mx0;
  assign _02925_ = cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_39_mx1;
  assign _02926_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) cvt_else_equal_tmp_39_mx1;
  assign _02927_ = FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02928_ = FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02929_ = FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02930_ = FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02931_ = FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02932_ = FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02933_ = FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02934_ = FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02935_ = FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02936_ = FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02937_ = FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02938_ = FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02939_ = FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02940_ = FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02941_ = FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_dcpl_407;
  assign _02942_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_896_rgt;
  assign _02943_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  assign _02944_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  assign _02945_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  assign _02946_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_954_rgt;
  assign _02947_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0;
  assign _02948_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  assign _02949_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_984_rgt;
  assign _02950_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_987_rgt;
  assign _02951_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0;
  assign _02952_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) and_1009_rgt;
  assign _02953_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  assign _02954_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  assign _02955_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0;
  assign _02956_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  assign _02957_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  assign _02958_ = FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_mux_56_nl;
  assign _02959_ = FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02960_ = IntShiftRightSat_49U_6U_17U_o_16_1_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02961_ = FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_1_mx1;
  assign _02962_ = IntShiftRightSat_49U_6U_17U_o_16_2_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_1_mx1;
  assign _02963_ = FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02964_ = IntShiftRightSat_49U_6U_17U_o_16_3_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02965_ = FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_3_mx1;
  assign _02966_ = IntShiftRightSat_49U_6U_17U_o_16_4_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_3_mx1;
  assign _02967_ = FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02968_ = IntShiftRightSat_49U_6U_17U_o_16_5_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02969_ = FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_5_mx1;
  assign _02970_ = IntShiftRightSat_49U_6U_17U_o_16_6_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_5_mx1;
  assign _02971_ = FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_6_mx1;
  assign _02972_ = IntShiftRightSat_49U_6U_17U_o_16_7_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_6_mx1;
  assign _02973_ = FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_7_mx1;
  assign _02974_ = IntShiftRightSat_49U_6U_17U_o_16_8_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_7_mx1;
  assign _02975_ = FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02976_ = IntShiftRightSat_49U_6U_17U_o_16_9_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs;
  assign _02977_ = FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_9_mx1;
  assign _02978_ = IntShiftRightSat_49U_6U_17U_o_16_10_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_9_mx1;
  assign _02979_ = FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_10_mx1;
  assign _02980_ = IntShiftRightSat_49U_6U_17U_o_16_11_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_10_mx1;
  assign _02981_ = FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_11_mx1;
  assign _02982_ = IntShiftRightSat_49U_6U_17U_o_16_12_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_11_mx1;
  assign _02983_ = FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_9_mx1;
  assign _02984_ = IntShiftRightSat_49U_6U_17U_o_16_13_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_9_mx1;
  assign _02985_ = IntShiftRightSat_49U_6U_17U_o_16_14_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_13_mx1;
  assign _02986_ = FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_14_mx1;
  assign _02987_ = IntShiftRightSat_49U_6U_17U_o_16_15_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_14_mx1;
  assign _02988_ = FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_13_mx1;
  assign _02989_ = IntShiftRightSat_49U_6U_17U_o_16_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) cvt_else_nor_dfs_13_mx1;
  assign _02990_ = IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_327;
  assign _02991_ = IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_333;
  assign _02992_ = IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_327;
  assign _02993_ = IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_339;
  assign _02994_ = IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_327;
  assign _02995_ = IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_357;
  assign _02996_ = IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_369;
  assign _02997_ = IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_381;
  assign _02998_ = IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_327;
  assign _02999_ = IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_399;
  assign _03000_ = IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_393;
  assign _03001_ = IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_387;
  assign _03002_ = IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_375;
  assign _03003_ = IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_363;
  assign _03004_ = IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cvt_asn_351;
  assign _03005_ = chn_idata_data_sva_3_495_479_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24266" *) cfg_mode_eql_1_sva_6;
  assign _03006_ = SetToInf_5U_10U_SetToInf_5U_10U_or_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_323;
  assign _03007_ = SetToInf_5U_10U_SetToInf_5U_10U_or_1_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_329;
  assign _03008_ = SetToInf_5U_10U_SetToInf_5U_10U_or_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_323;
  assign _03009_ = SetToInf_5U_10U_SetToInf_5U_10U_or_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_335;
  assign _03010_ = SetToInf_5U_10U_SetToInf_5U_10U_or_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_323;
  assign _03011_ = SetToInf_5U_10U_SetToInf_5U_10U_or_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_353;
  assign _03012_ = SetToInf_5U_10U_SetToInf_5U_10U_or_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_365;
  assign _03013_ = SetToInf_5U_10U_SetToInf_5U_10U_or_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_377;
  assign _03014_ = SetToInf_5U_10U_SetToInf_5U_10U_or_8_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_323;
  assign _03015_ = SetToInf_5U_10U_SetToInf_5U_10U_or_9_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_371;
  assign _03016_ = SetToInf_5U_10U_SetToInf_5U_10U_or_10_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_389;
  assign _03017_ = SetToInf_5U_10U_SetToInf_5U_10U_or_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_383;
  assign _03018_ = SetToInf_5U_10U_SetToInf_5U_10U_or_12_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_371;
  assign _03019_ = SetToInf_5U_10U_SetToInf_5U_10U_or_13_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_359;
  assign _03020_ = SetToInf_5U_10U_SetToInf_5U_10U_or_14_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_347;
  assign _03021_ = IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) cvt_asn_345;
  assign _03022_ = reg_chn_idata_data_sva_3_15_0_1_reg[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03023_ = chn_idata_data_sva_3_47_31_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03024_ = chn_idata_data_sva_3_79_63_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03025_ = chn_idata_data_sva_3_111_95_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03026_ = chn_idata_data_sva_3_143_127_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03027_ = chn_idata_data_sva_3_175_159_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03028_ = chn_idata_data_sva_3_207_191_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03029_ = chn_idata_data_sva_3_239_223_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03030_ = chn_idata_data_sva_3_271_255_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03031_ = chn_idata_data_sva_3_303_287_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03032_ = chn_idata_data_sva_3_335_319_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03033_ = chn_idata_data_sva_3_367_351_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03034_ = chn_idata_data_sva_3_399_383_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03035_ = chn_idata_data_sva_3_431_415_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03036_ = chn_idata_data_sva_3_463_447_1[15] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cfg_mode_eql_1_sva_6;
  assign _03037_ = SetToInf_5U_10U_SetToInf_5U_10U_or_15_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) cvt_asn_341;
  assign _03038_ = FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03039_ = FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03040_ = FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03041_ = FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03042_ = FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03043_ = FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03044_ = FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03045_ = FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03046_ = FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03047_ = FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03048_ = FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03049_ = FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03050_ = FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03051_ = FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03052_ = FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03053_ = FpFloatToInt_16U_5U_10U_internal_int_0_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) cvt_asn_321;
  assign _03054_ = reg_chn_idata_data_sva_3_15_0_1_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_cse;
  assign _03055_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_2_cse;
  assign _03056_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_cse;
  assign _03057_ = FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[13] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_6_cse;
  assign _03058_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_cse;
  assign _03059_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_10_cse;
  assign _03060_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_12_cse;
  assign _03061_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_14_cse;
  assign _03062_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_cse;
  assign _03063_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_18_cse;
  assign _03064_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_20_cse;
  assign _03065_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_22_cse;
  assign _03066_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_24_cse;
  assign _03067_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_26_cse;
  assign _03068_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_28_cse;
  assign _03069_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) cvt_or_30_cse;
  assign _03070_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt, IntSaturation_17U_16U_o_and_31_rgt };
  assign _03071_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt, IntSaturation_17U_16U_o_and_29_rgt };
  assign _03072_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt, IntSaturation_17U_16U_o_and_27_rgt };
  assign _03073_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt, IntSaturation_17U_16U_o_and_25_rgt };
  assign _03074_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt, IntSaturation_17U_16U_o_and_23_rgt };
  assign _03075_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt, IntSaturation_17U_16U_o_and_21_rgt };
  assign _03076_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt, IntSaturation_17U_16U_o_and_19_rgt };
  assign _03077_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt, IntSaturation_17U_16U_o_and_17_rgt };
  assign _03078_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt, IntSaturation_17U_16U_o_and_15_rgt };
  assign _03079_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt, IntSaturation_17U_16U_o_and_13_rgt };
  assign _03080_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt, IntSaturation_17U_16U_o_and_11_rgt };
  assign _03081_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt, IntSaturation_17U_16U_o_and_9_rgt };
  assign _03082_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt, IntSaturation_17U_16U_o_and_7_rgt };
  assign _03083_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt, IntSaturation_17U_16U_o_and_5_rgt };
  assign _03084_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt, IntSaturation_17U_16U_o_and_3_rgt };
  assign _03085_ = 14'b11111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt, IntSaturation_17U_16U_o_and_1_rgt };
  assign _03086_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl, mux_1752_nl };
  assign _03087_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl, mux_1758_nl };
  assign _03088_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse };
  assign _03089_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse };
  assign _03090_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse, mux_1762_cse };
  assign _03091_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl };
  assign _03092_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl, mux_1780_nl };
  assign _03093_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl, mux_1788_nl };
  assign _03094_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl, mux_1791_nl };
  assign _03095_ = IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl, and_843_nl };
  assign _03096_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl, mux_1808_nl };
  assign _03097_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24281" *) { mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl, mux_1817_nl };
  assign _03098_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt, IntSaturation_17U_16U_and_31_rgt };
  assign _03099_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt, IntSaturation_17U_16U_and_29_rgt };
  assign _03100_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt, IntSaturation_17U_16U_and_27_rgt };
  assign _03101_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt, IntSaturation_17U_16U_and_25_rgt };
  assign _03102_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt, IntSaturation_17U_16U_and_23_rgt };
  assign _03103_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt, IntSaturation_17U_16U_and_21_rgt };
  assign _03104_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt, IntSaturation_17U_16U_and_19_rgt };
  assign _03105_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt, IntSaturation_17U_16U_and_17_rgt };
  assign _03106_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt, IntSaturation_17U_16U_and_15_rgt };
  assign _03107_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt, IntSaturation_17U_16U_and_13_rgt };
  assign _03108_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt, IntSaturation_17U_16U_and_11_rgt };
  assign _03109_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt, IntSaturation_17U_16U_and_9_rgt };
  assign _03110_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt, IntSaturation_17U_16U_and_7_rgt };
  assign _03111_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt, IntSaturation_17U_16U_and_5_rgt };
  assign _03112_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt, IntSaturation_17U_16U_and_3_rgt };
  assign _03113_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt, IntSaturation_17U_16U_and_1_rgt };
  assign _03114_ = IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl, and_699_nl };
  assign _03115_ = IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl, and_714_nl };
  assign _03116_ = IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl, and_729_nl };
  assign _03117_ = IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl, and_744_nl };
  assign _03118_ = IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl, and_759_nl };
  assign _03119_ = IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl, and_783_nl };
  assign _03120_ = IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl, and_797_nl };
  assign _03121_ = IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl, and_811_nl };
  assign _03122_ = IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl, and_826_nl };
  assign _03123_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl, and_840_nl };
  assign _03124_ = IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl, and_859_nl };
  assign _03125_ = IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) { and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl, and_876_nl };
  assign _03126_ = IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt };
  assign _03127_ = IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt };
  assign _03128_ = IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt };
  assign _03129_ = IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt };
  assign _03130_ = IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt };
  assign _03131_ = IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt };
  assign _03132_ = IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt };
  assign _03133_ = IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt };
  assign _03134_ = IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt };
  assign _03135_ = IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt };
  assign _03136_ = IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt };
  assign _03137_ = IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt };
  assign _03138_ = IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt };
  assign _03139_ = IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt };
  assign _03140_ = IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt };
  assign _03141_ = IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt, IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt };
  assign _03142_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl, and_696_nl };
  assign _03143_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl, and_711_nl };
  assign _03144_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl, and_726_nl };
  assign _03145_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl, and_741_nl };
  assign _03146_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl, and_756_nl };
  assign _03147_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl, and_780_nl };
  assign _03148_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl, and_794_nl };
  assign _03149_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl, and_808_nl };
  assign _03150_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl, and_823_nl };
  assign _03151_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_63_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl, or_4348_nl };
  assign _03152_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl, and_856_nl };
  assign _03153_ = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) { and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl, and_873_nl };
  assign _03154_ = IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24297" *) { FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2 };
  assign _03155_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24297" *) { mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl, mux_1889_nl };
  assign _03156_ = IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24297" *) { and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl, and_908_nl };
  assign _03157_ = IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *) { FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1, FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1 };
  assign _03158_ = IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *) { and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420, and_dcpl_420 };
  assign _03159_ = IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *) { and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425 };
  assign _03160_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *) { FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl, FpFloatToInt_16U_5U_10U_o_int_and_28_nl };
  assign _03161_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *) { FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl, FpFloatToInt_16U_5U_10U_o_int_and_23_nl };
  assign _03162_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *) { FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl, FpFloatToInt_16U_5U_10U_o_int_and_15_nl };
  assign _03163_ = FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *) { FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl, FpFloatToInt_16U_5U_10U_and_7_nl };
  assign _03164_ = FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *) { FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl, FpFloatToInt_16U_5U_10U_and_27_nl };
  assign _03165_ = FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *) { FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl, FpFloatToInt_16U_5U_10U_and_1_nl };
  assign _03166_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *) { FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl, FpFloatToInt_16U_5U_10U_and_38_nl };
  assign _03167_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *) { FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl, FpFloatToInt_16U_5U_10U_and_58_nl };
  assign _03168_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *) { FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl, FpFloatToInt_16U_5U_10U_and_32_nl };
  assign _03169_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *) { FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl, FpFloatToInt_16U_5U_10U_and_37_nl };
  assign _03170_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *) { FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl, FpFloatToInt_16U_5U_10U_and_57_nl };
  assign _03171_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *) { FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl, FpFloatToInt_16U_5U_10U_and_nl };
  assign _03172_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_1_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl, mux_1831_nl };
  assign _03173_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422 };
  assign _03174_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse };
  assign _03175_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422 };
  assign _03176_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl, mux_1867_nl };
  assign _03177_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse };
  assign _03178_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse };
  assign _03179_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_8_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl, mux_1909_nl };
  assign _03180_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_9_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse, mux_1852_cse };
  assign _03181_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_10_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl, mux_1933_nl };
  assign _03182_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422, not_tmp_2422 };
  assign _03183_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_12_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse };
  assign _03184_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_13_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24317" *) { mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse, mux_1882_cse };
  assign _03185_ = IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl, and_921_nl };
  assign _03186_ = IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446 };
  assign _03187_ = IntShiftRightSat_49U_6U_17U_o_15_1_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl, and_949_nl };
  assign _03188_ = IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446 };
  assign _03189_ = IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl, and_966_nl };
  assign _03190_ = IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse };
  assign _03191_ = IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse };
  assign _03192_ = IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl, and_1004_nl };
  assign _03193_ = IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse, and_978_cse };
  assign _03194_ = IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl, and_1027_nl };
  assign _03195_ = IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446, and_dcpl_446 };
  assign _03196_ = IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse };
  assign _03197_ = IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) { and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse, and_1039_cse };
  assign _03198_ = IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl, and_916_nl };
  assign _03199_ = IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425 };
  assign _03200_ = IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl, and_945_nl };
  assign _03201_ = IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425 };
  assign _03202_ = IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl, and_961_nl };
  assign _03203_ = IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl };
  assign _03204_ = IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl };
  assign _03205_ = IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl, and_999_nl };
  assign _03206_ = IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl, and_1013_nl };
  assign _03207_ = IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl };
  assign _03208_ = IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425, and_dcpl_425 };
  assign _03209_ = IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl };
  assign _03210_ = IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) { and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl, and_1023_nl };
  assign _03211_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl, FpFloatToInt_16U_5U_10U_o_int_and_nl };
  assign _03212_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl, FpFloatToInt_16U_5U_10U_o_int_and_29_nl };
  assign _03213_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl, FpFloatToInt_16U_5U_10U_o_int_and_27_nl };
  assign _03214_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl, FpFloatToInt_16U_5U_10U_o_int_and_26_nl };
  assign _03215_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl, FpFloatToInt_16U_5U_10U_o_int_and_25_nl };
  assign _03216_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl, FpFloatToInt_16U_5U_10U_o_int_and_24_nl };
  assign _03217_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl, FpFloatToInt_16U_5U_10U_o_int_and_22_nl };
  assign _03218_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl, FpFloatToInt_16U_5U_10U_o_int_and_21_nl };
  assign _03219_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl, FpFloatToInt_16U_5U_10U_o_int_and_20_nl };
  assign _03220_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl, FpFloatToInt_16U_5U_10U_o_int_and_19_nl };
  assign _03221_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl, FpFloatToInt_16U_5U_10U_o_int_and_18_nl };
  assign _03222_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl, FpFloatToInt_16U_5U_10U_o_int_and_17_nl };
  assign _03223_ = 15'b100000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) { FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl, FpFloatToInt_16U_5U_10U_o_int_and_16_nl };
  assign _03224_ = FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl, FpFloatToInt_16U_5U_10U_and_3_nl };
  assign _03225_ = FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl, FpFloatToInt_16U_5U_10U_and_5_nl };
  assign _03226_ = FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl, FpFloatToInt_16U_5U_10U_and_31_nl };
  assign _03227_ = FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl, FpFloatToInt_16U_5U_10U_and_9_nl };
  assign _03228_ = FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl, FpFloatToInt_16U_5U_10U_and_29_nl };
  assign _03229_ = FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl, FpFloatToInt_16U_5U_10U_and_11_nl };
  assign _03230_ = FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl, FpFloatToInt_16U_5U_10U_and_13_nl };
  assign _03231_ = FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl, FpFloatToInt_16U_5U_10U_and_25_nl };
  assign _03232_ = FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl, FpFloatToInt_16U_5U_10U_and_15_nl };
  assign _03233_ = FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl, FpFloatToInt_16U_5U_10U_and_23_nl };
  assign _03234_ = FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl, FpFloatToInt_16U_5U_10U_and_17_nl };
  assign _03235_ = FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl, FpFloatToInt_16U_5U_10U_and_21_nl };
  assign _03236_ = FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) { FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl, FpFloatToInt_16U_5U_10U_and_19_nl };
  assign _03237_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl, FpFloatToInt_16U_5U_10U_and_34_nl };
  assign _03238_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl, FpFloatToInt_16U_5U_10U_and_36_nl };
  assign _03239_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl, FpFloatToInt_16U_5U_10U_and_62_nl };
  assign _03240_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl, FpFloatToInt_16U_5U_10U_and_40_nl };
  assign _03241_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl, FpFloatToInt_16U_5U_10U_and_60_nl };
  assign _03242_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl, FpFloatToInt_16U_5U_10U_and_42_nl };
  assign _03243_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl, FpFloatToInt_16U_5U_10U_and_44_nl };
  assign _03244_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl, FpFloatToInt_16U_5U_10U_and_56_nl };
  assign _03245_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl, FpFloatToInt_16U_5U_10U_and_46_nl };
  assign _03246_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl, FpFloatToInt_16U_5U_10U_and_54_nl };
  assign _03247_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl, FpFloatToInt_16U_5U_10U_and_48_nl };
  assign _03248_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl, FpFloatToInt_16U_5U_10U_and_52_nl };
  assign _03249_ = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva[15:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) { FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl, FpFloatToInt_16U_5U_10U_and_50_nl };
  assign _03250_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl, FpFloatToInt_16U_5U_10U_and_33_nl };
  assign _03251_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl, FpFloatToInt_16U_5U_10U_and_35_nl };
  assign _03252_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl, FpFloatToInt_16U_5U_10U_and_61_nl };
  assign _03253_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl, FpFloatToInt_16U_5U_10U_and_39_nl };
  assign _03254_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl, FpFloatToInt_16U_5U_10U_and_59_nl };
  assign _03255_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl, FpFloatToInt_16U_5U_10U_and_41_nl };
  assign _03256_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl, FpFloatToInt_16U_5U_10U_and_43_nl };
  assign _03257_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl, FpFloatToInt_16U_5U_10U_and_55_nl };
  assign _03258_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl, FpFloatToInt_16U_5U_10U_and_45_nl };
  assign _03259_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl, FpFloatToInt_16U_5U_10U_and_53_nl };
  assign _03260_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl, FpFloatToInt_16U_5U_10U_and_47_nl };
  assign _03261_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl, FpFloatToInt_16U_5U_10U_and_51_nl };
  assign _03262_ = FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva[14:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) { FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl, FpFloatToInt_16U_5U_10U_and_49_nl };
  assign _03263_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_14_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24334" *) { _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0], _00000_[0] };
  assign _03264_ = FpFloatToInt_16U_5U_10U_o_int_mux1h_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24335" *) { _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1], _00000_[1] };
  assign _03265_ = chn_idata_data_sva_2_15_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24336" *) { and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl, and_1179_nl };
  assign _03266_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_164_cse, nand_164_cse, nand_164_cse, nand_164_cse };
  assign _03267_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_162_cse, nand_162_cse, nand_162_cse, nand_162_cse };
  assign _03268_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_160_cse, nand_160_cse, nand_160_cse, nand_160_cse };
  assign _03269_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_158_cse, nand_158_cse, nand_158_cse, nand_158_cse };
  assign _03270_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_156_cse, nand_156_cse, nand_156_cse, nand_156_cse };
  assign _03271_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_153_cse, nand_153_cse, nand_153_cse, nand_153_cse };
  assign _03272_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_151_cse, nand_151_cse, nand_151_cse, nand_151_cse };
  assign _03273_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_149_cse, nand_149_cse, nand_149_cse, nand_149_cse };
  assign _03274_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_147_cse, nand_147_cse, nand_147_cse, nand_147_cse };
  assign _03275_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_145_cse, nand_145_cse, nand_145_cse, nand_145_cse };
  assign _03276_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_143_cse, nand_143_cse, nand_143_cse, nand_143_cse };
  assign _03277_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_141_cse, nand_141_cse, nand_141_cse, nand_141_cse };
  assign _03278_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_139_cse, nand_139_cse, nand_139_cse, nand_139_cse };
  assign _03279_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_137_cse, nand_137_cse, nand_137_cse, nand_137_cse };
  assign _03280_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_135_cse, nand_135_cse, nand_135_cse, nand_135_cse };
  assign _03281_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24348" *) { nand_133_cse, nand_133_cse, nand_133_cse, nand_133_cse };
  assign _03282_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl };
  assign _03283_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl };
  assign _03284_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl };
  assign _03285_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl };
  assign _03286_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl };
  assign _03287_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl };
  assign _03288_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl };
  assign _03289_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl };
  assign _03290_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl };
  assign _03291_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl };
  assign _03292_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl };
  assign _03293_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl };
  assign _03294_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl };
  assign _03295_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl };
  assign _03296_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl };
  assign _03297_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl };
  assign _03298_ = chn_idata_data_sva_1_27_0_1[26:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl };
  assign _03299_ = chn_idata_data_sva_1_59_31_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl };
  assign _03300_ = chn_idata_data_sva_1_91_63_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl };
  assign _03301_ = chn_idata_data_sva_1_123_95_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl };
  assign _03302_ = chn_idata_data_sva_1_155_127_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl };
  assign _03303_ = chn_idata_data_sva_1_187_159_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl };
  assign _03304_ = chn_idata_data_sva_1_219_191_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl };
  assign _03305_ = chn_idata_data_sva_1_251_223_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl };
  assign _03306_ = chn_idata_data_sva_1_283_255_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl };
  assign _03307_ = chn_idata_data_sva_1_315_287_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl };
  assign _03308_ = chn_idata_data_sva_1_347_319_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl };
  assign _03309_ = chn_idata_data_sva_1_379_351_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl };
  assign _03310_ = chn_idata_data_sva_1_411_383_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl };
  assign _03311_ = chn_idata_data_sva_1_443_415_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl };
  assign _03312_ = chn_idata_data_sva_1_475_447_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl };
  assign _03313_ = chn_idata_data_sva_1_507_479_1[27:24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl, FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl };
  assign _03314_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc };
  assign _03315_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc };
  assign _03316_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc };
  assign _03317_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc };
  assign _03318_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc };
  assign _03319_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc };
  assign _03320_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc };
  assign _03321_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc };
  assign _03322_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc };
  assign _03323_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc };
  assign _03324_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc };
  assign _03325_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc };
  assign _03326_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc };
  assign _03327_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc };
  assign _03328_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc };
  assign _03329_ = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) { FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc, FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc };
  assign _03330_ = reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_tmp_4102, or_tmp_4102, or_tmp_4102, or_tmp_4102 };
  assign _03331_ = reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5175_tmp, or_5175_tmp, or_5175_tmp, or_5175_tmp };
  assign _03332_ = reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5177_tmp, or_5177_tmp, or_5177_tmp, or_5177_tmp };
  assign _03333_ = reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5181_tmp, or_5181_tmp, or_5181_tmp, or_5181_tmp };
  assign _03334_ = reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5174_tmp, or_5174_tmp, or_5174_tmp, or_5174_tmp };
  assign _03335_ = reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5176_tmp, or_5176_tmp, or_5176_tmp, or_5176_tmp };
  assign _03336_ = reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5178_tmp, or_5178_tmp, or_5178_tmp, or_5178_tmp };
  assign _03337_ = reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5179_tmp, or_5179_tmp, or_5179_tmp, or_5179_tmp };
  assign _03338_ = reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5180_tmp, or_5180_tmp, or_5180_tmp, or_5180_tmp };
  assign _03339_ = reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5182_tmp, or_5182_tmp, or_5182_tmp, or_5182_tmp };
  assign _03340_ = reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5183_tmp, or_5183_tmp, or_5183_tmp, or_5183_tmp };
  assign _03341_ = reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5184_tmp, or_5184_tmp, or_5184_tmp, or_5184_tmp };
  assign _03342_ = reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5185_tmp, or_5185_tmp, or_5185_tmp, or_5185_tmp };
  assign _03343_ = reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5186_tmp, or_5186_tmp, or_5186_tmp, or_5186_tmp };
  assign _03344_ = reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5188_tmp, or_5188_tmp, or_5188_tmp, or_5188_tmp };
  assign _03345_ = reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24365" *) { or_5187_tmp, or_5187_tmp, or_5187_tmp, or_5187_tmp };
  assign _03346_ = { IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03347_ = { IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03348_ = { IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03349_ = { IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03350_ = { IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3148_nl, and_3148_nl, and_3148_nl, and_3148_nl };
  assign _03351_ = { IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { cvt_asn_339, cvt_asn_339, cvt_asn_339, cvt_asn_339 };
  assign _03352_ = { IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3136_nl, and_3136_nl, and_3136_nl, and_3136_nl };
  assign _03353_ = { IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3133_nl, and_3133_nl, and_3133_nl, and_3133_nl };
  assign _03354_ = { IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3130_nl, and_3130_nl, and_3130_nl, and_3130_nl };
  assign _03355_ = { IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3124_nl, and_3124_nl, and_3124_nl, and_3124_nl };
  assign _03356_ = { IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3121_nl, and_3121_nl, and_3121_nl, and_3121_nl };
  assign _03357_ = { IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3118_nl, and_3118_nl, and_3118_nl, and_3118_nl };
  assign _03358_ = { IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3115_nl, and_3115_nl, and_3115_nl, and_3115_nl };
  assign _03359_ = { IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3112_nl, and_3112_nl, and_3112_nl, and_3112_nl };
  assign _03360_ = chn_idata_data_sva_3_495_479_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03361_ = { IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) { and_3109_nl, and_3109_nl, and_3109_nl, and_3109_nl };
  assign _03362_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_262_nl, cvt_and_262_nl, cvt_and_262_nl, cvt_and_262_nl };
  assign _03363_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_258_nl, cvt_and_258_nl, cvt_and_258_nl, cvt_and_258_nl };
  assign _03364_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_254_nl, cvt_and_254_nl, cvt_and_254_nl, cvt_and_254_nl };
  assign _03365_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_246_nl, cvt_and_246_nl, cvt_and_246_nl, cvt_and_246_nl };
  assign _03366_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_260_nl, cvt_and_260_nl, cvt_and_260_nl, cvt_and_260_nl };
  assign _03367_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_256_nl, cvt_and_256_nl, cvt_and_256_nl, cvt_and_256_nl };
  assign _03368_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_252_nl, cvt_and_252_nl, cvt_and_252_nl, cvt_and_252_nl };
  assign _03369_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_250_nl, cvt_and_250_nl, cvt_and_250_nl, cvt_and_250_nl };
  assign _03370_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_248_nl, cvt_and_248_nl, cvt_and_248_nl, cvt_and_248_nl };
  assign _03371_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_244_nl, cvt_and_244_nl, cvt_and_244_nl, cvt_and_244_nl };
  assign _03372_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_242_nl, cvt_and_242_nl, cvt_and_242_nl, cvt_and_242_nl };
  assign _03373_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_240_nl, cvt_and_240_nl, cvt_and_240_nl, cvt_and_240_nl };
  assign _03374_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_238_nl, cvt_and_238_nl, cvt_and_238_nl, cvt_and_238_nl };
  assign _03375_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_236_nl, cvt_and_236_nl, cvt_and_236_nl, cvt_and_236_nl };
  assign _03376_ = { IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { and_3105_nl, and_3105_nl, and_3105_nl, and_3105_nl };
  assign _03377_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) { cvt_and_234_nl, cvt_and_234_nl, cvt_and_234_nl, cvt_and_234_nl };
  assign _03378_ = { _04700_, _04700_, _04700_, _04700_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_261_nl, cvt_and_261_nl, cvt_and_261_nl, cvt_and_261_nl };
  assign _03379_ = { _04704_, _04704_, _04704_, _04704_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_257_nl, cvt_and_257_nl, cvt_and_257_nl, cvt_and_257_nl };
  assign _03380_ = { _04708_, _04708_, _04708_, _04708_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_253_nl, cvt_and_253_nl, cvt_and_253_nl, cvt_and_253_nl };
  assign _03381_ = { _04716_, _04716_, _04716_, _04716_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_245_nl, cvt_and_245_nl, cvt_and_245_nl, cvt_and_245_nl };
  assign _03382_ = { _04702_, _04702_, _04702_, _04702_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_259_nl, cvt_and_259_nl, cvt_and_259_nl, cvt_and_259_nl };
  assign _03383_ = { _04706_, _04706_, _04706_, _04706_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_255_nl, cvt_and_255_nl, cvt_and_255_nl, cvt_and_255_nl };
  assign _03384_ = { _04710_, _04710_, _04710_, _04710_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_251_nl, cvt_and_251_nl, cvt_and_251_nl, cvt_and_251_nl };
  assign _03385_ = { _04712_, _04712_, _04712_, _04712_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_249_nl, cvt_and_249_nl, cvt_and_249_nl, cvt_and_249_nl };
  assign _03386_ = { _04714_, _04714_, _04714_, _04714_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_247_nl, cvt_and_247_nl, cvt_and_247_nl, cvt_and_247_nl };
  assign _03387_ = { _04718_, _04718_, _04718_, _04718_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_243_nl, cvt_and_243_nl, cvt_and_243_nl, cvt_and_243_nl };
  assign _03388_ = { _04720_, _04720_, _04720_, _04720_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_241_nl, cvt_and_241_nl, cvt_and_241_nl, cvt_and_241_nl };
  assign _03389_ = { _04722_, _04722_, _04722_, _04722_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_239_nl, cvt_and_239_nl, cvt_and_239_nl, cvt_and_239_nl };
  assign _03390_ = { _04724_, _04724_, _04724_, _04724_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_237_nl, cvt_and_237_nl, cvt_and_237_nl, cvt_and_237_nl };
  assign _03391_ = { _04726_, _04726_, _04726_, _04726_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_235_nl, cvt_and_235_nl, cvt_and_235_nl, cvt_and_235_nl };
  assign _03392_ = 4'b1110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_232_nl, cvt_and_232_nl, cvt_and_232_nl, cvt_and_232_nl };
  assign _03393_ = { _04728_, _04728_, _04728_, _04728_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) { cvt_and_233_nl, cvt_and_233_nl, cvt_and_233_nl, cvt_and_233_nl };
  assign _03394_ = reg_chn_idata_data_sva_3_15_0_1_reg[3:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03395_ = chn_idata_data_sva_3_79_63_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03396_ = chn_idata_data_sva_3_143_127_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03397_ = chn_idata_data_sva_3_271_255_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03398_ = chn_idata_data_sva_3_47_31_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03399_ = chn_idata_data_sva_3_111_95_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03400_ = chn_idata_data_sva_3_175_159_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03401_ = chn_idata_data_sva_3_207_191_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03402_ = chn_idata_data_sva_3_239_223_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03403_ = chn_idata_data_sva_3_303_287_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03404_ = chn_idata_data_sva_3_335_319_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03405_ = chn_idata_data_sva_3_367_351_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03406_ = chn_idata_data_sva_3_399_383_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03407_ = chn_idata_data_sva_3_431_415_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03408_ = { _04730_, _04730_, _04730_, _04730_ } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cvt_and_231_nl, cvt_and_231_nl, cvt_and_231_nl, cvt_and_231_nl };
  assign _03409_ = chn_idata_data_sva_3_463_447_1[14:11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03410_ = { reg_chn_idata_data_sva_3_15_0_1_reg[2:0], reg_chn_idata_data_sva_3_15_0_2_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03411_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03412_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03413_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03414_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse };
  assign _03415_ = FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[12:9] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { and_3140_nl, and_3140_nl, and_3140_nl, and_3140_nl };
  assign _03416_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse };
  assign _03417_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse };
  assign _03418_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { and_3128_nl, and_3128_nl, and_3128_nl, and_3128_nl };
  assign _03419_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse };
  assign _03420_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse };
  assign _03421_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { and_3116_nl, and_3116_nl, and_3116_nl, and_3116_nl };
  assign _03422_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse };
  assign _03423_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { and_3110_nl, and_3110_nl, and_3110_nl, and_3110_nl };
  assign _03424_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { and_3104_nl, and_3104_nl, and_3104_nl, and_3104_nl };
  assign _03425_ = { reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[2:0], reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[9] } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) { cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse };
  assign _03426_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03427_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03428_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03429_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03430_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03431_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03432_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03433_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03434_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03435_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03436_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03437_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03438_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03439_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03440_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03441_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24381" *) { _00002_[0], _00002_[0], _00002_[0], _00002_[0], _00002_[0] };
  assign _03442_ = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_31_nl, FpIntToFloat_17U_5U_10U_o_expo_and_31_nl, FpIntToFloat_17U_5U_10U_o_expo_and_31_nl, FpIntToFloat_17U_5U_10U_o_expo_and_31_nl, FpIntToFloat_17U_5U_10U_o_expo_and_31_nl };
  assign _03443_ = cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_29_nl, FpIntToFloat_17U_5U_10U_o_expo_and_29_nl, FpIntToFloat_17U_5U_10U_o_expo_and_29_nl, FpIntToFloat_17U_5U_10U_o_expo_and_29_nl, FpIntToFloat_17U_5U_10U_o_expo_and_29_nl };
  assign _03444_ = cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_27_nl, FpIntToFloat_17U_5U_10U_o_expo_and_27_nl, FpIntToFloat_17U_5U_10U_o_expo_and_27_nl, FpIntToFloat_17U_5U_10U_o_expo_and_27_nl, FpIntToFloat_17U_5U_10U_o_expo_and_27_nl };
  assign _03445_ = cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_25_nl, FpIntToFloat_17U_5U_10U_o_expo_and_25_nl, FpIntToFloat_17U_5U_10U_o_expo_and_25_nl, FpIntToFloat_17U_5U_10U_o_expo_and_25_nl, FpIntToFloat_17U_5U_10U_o_expo_and_25_nl };
  assign _03446_ = cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_23_nl, FpIntToFloat_17U_5U_10U_o_expo_and_23_nl, FpIntToFloat_17U_5U_10U_o_expo_and_23_nl, FpIntToFloat_17U_5U_10U_o_expo_and_23_nl, FpIntToFloat_17U_5U_10U_o_expo_and_23_nl };
  assign _03447_ = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_21_nl, FpIntToFloat_17U_5U_10U_o_expo_and_21_nl, FpIntToFloat_17U_5U_10U_o_expo_and_21_nl, FpIntToFloat_17U_5U_10U_o_expo_and_21_nl, FpIntToFloat_17U_5U_10U_o_expo_and_21_nl };
  assign _03448_ = cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_19_nl, FpIntToFloat_17U_5U_10U_o_expo_and_19_nl, FpIntToFloat_17U_5U_10U_o_expo_and_19_nl, FpIntToFloat_17U_5U_10U_o_expo_and_19_nl, FpIntToFloat_17U_5U_10U_o_expo_and_19_nl };
  assign _03449_ = cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_17_nl, FpIntToFloat_17U_5U_10U_o_expo_and_17_nl, FpIntToFloat_17U_5U_10U_o_expo_and_17_nl, FpIntToFloat_17U_5U_10U_o_expo_and_17_nl, FpIntToFloat_17U_5U_10U_o_expo_and_17_nl };
  assign _03450_ = cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_15_nl, FpIntToFloat_17U_5U_10U_o_expo_and_15_nl, FpIntToFloat_17U_5U_10U_o_expo_and_15_nl, FpIntToFloat_17U_5U_10U_o_expo_and_15_nl, FpIntToFloat_17U_5U_10U_o_expo_and_15_nl };
  assign _03451_ = cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_13_nl, FpIntToFloat_17U_5U_10U_o_expo_and_13_nl, FpIntToFloat_17U_5U_10U_o_expo_and_13_nl, FpIntToFloat_17U_5U_10U_o_expo_and_13_nl, FpIntToFloat_17U_5U_10U_o_expo_and_13_nl };
  assign _03452_ = cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_11_nl, FpIntToFloat_17U_5U_10U_o_expo_and_11_nl, FpIntToFloat_17U_5U_10U_o_expo_and_11_nl, FpIntToFloat_17U_5U_10U_o_expo_and_11_nl, FpIntToFloat_17U_5U_10U_o_expo_and_11_nl };
  assign _03453_ = cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_9_nl, FpIntToFloat_17U_5U_10U_o_expo_and_9_nl, FpIntToFloat_17U_5U_10U_o_expo_and_9_nl, FpIntToFloat_17U_5U_10U_o_expo_and_9_nl, FpIntToFloat_17U_5U_10U_o_expo_and_9_nl };
  assign _03454_ = cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_7_nl, FpIntToFloat_17U_5U_10U_o_expo_and_7_nl, FpIntToFloat_17U_5U_10U_o_expo_and_7_nl, FpIntToFloat_17U_5U_10U_o_expo_and_7_nl, FpIntToFloat_17U_5U_10U_o_expo_and_7_nl };
  assign _03455_ = cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_5_nl, FpIntToFloat_17U_5U_10U_o_expo_and_5_nl, FpIntToFloat_17U_5U_10U_o_expo_and_5_nl, FpIntToFloat_17U_5U_10U_o_expo_and_5_nl, FpIntToFloat_17U_5U_10U_o_expo_and_5_nl };
  assign _03456_ = cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_3_nl, FpIntToFloat_17U_5U_10U_o_expo_and_3_nl, FpIntToFloat_17U_5U_10U_o_expo_and_3_nl, FpIntToFloat_17U_5U_10U_o_expo_and_3_nl, FpIntToFloat_17U_5U_10U_o_expo_and_3_nl };
  assign _03457_ = cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) { FpIntToFloat_17U_5U_10U_o_expo_and_1_nl, FpIntToFloat_17U_5U_10U_o_expo_and_1_nl, FpIntToFloat_17U_5U_10U_o_expo_and_1_nl, FpIntToFloat_17U_5U_10U_o_expo_and_1_nl, FpIntToFloat_17U_5U_10U_o_expo_and_1_nl };
  assign _03458_ = _00001_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_15_nl, FpIntToFloat_17U_5U_10U_o_expo_or_15_nl, FpIntToFloat_17U_5U_10U_o_expo_or_15_nl, FpIntToFloat_17U_5U_10U_o_expo_or_15_nl, FpIntToFloat_17U_5U_10U_o_expo_or_15_nl };
  assign _03459_ = _00003_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_14_nl, FpIntToFloat_17U_5U_10U_o_expo_or_14_nl, FpIntToFloat_17U_5U_10U_o_expo_or_14_nl, FpIntToFloat_17U_5U_10U_o_expo_or_14_nl, FpIntToFloat_17U_5U_10U_o_expo_or_14_nl };
  assign _03460_ = _00004_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_13_nl, FpIntToFloat_17U_5U_10U_o_expo_or_13_nl, FpIntToFloat_17U_5U_10U_o_expo_or_13_nl, FpIntToFloat_17U_5U_10U_o_expo_or_13_nl, FpIntToFloat_17U_5U_10U_o_expo_or_13_nl };
  assign _03461_ = _00005_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_12_nl, FpIntToFloat_17U_5U_10U_o_expo_or_12_nl, FpIntToFloat_17U_5U_10U_o_expo_or_12_nl, FpIntToFloat_17U_5U_10U_o_expo_or_12_nl, FpIntToFloat_17U_5U_10U_o_expo_or_12_nl };
  assign _03462_ = _00006_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_11_nl, FpIntToFloat_17U_5U_10U_o_expo_or_11_nl, FpIntToFloat_17U_5U_10U_o_expo_or_11_nl, FpIntToFloat_17U_5U_10U_o_expo_or_11_nl, FpIntToFloat_17U_5U_10U_o_expo_or_11_nl };
  assign _03463_ = _00007_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_10_nl, FpIntToFloat_17U_5U_10U_o_expo_or_10_nl, FpIntToFloat_17U_5U_10U_o_expo_or_10_nl, FpIntToFloat_17U_5U_10U_o_expo_or_10_nl, FpIntToFloat_17U_5U_10U_o_expo_or_10_nl };
  assign _03464_ = _00008_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_9_nl, FpIntToFloat_17U_5U_10U_o_expo_or_9_nl, FpIntToFloat_17U_5U_10U_o_expo_or_9_nl, FpIntToFloat_17U_5U_10U_o_expo_or_9_nl, FpIntToFloat_17U_5U_10U_o_expo_or_9_nl };
  assign _03465_ = _00009_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_8_nl, FpIntToFloat_17U_5U_10U_o_expo_or_8_nl, FpIntToFloat_17U_5U_10U_o_expo_or_8_nl, FpIntToFloat_17U_5U_10U_o_expo_or_8_nl, FpIntToFloat_17U_5U_10U_o_expo_or_8_nl };
  assign _03466_ = _00010_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_7_nl, FpIntToFloat_17U_5U_10U_o_expo_or_7_nl, FpIntToFloat_17U_5U_10U_o_expo_or_7_nl, FpIntToFloat_17U_5U_10U_o_expo_or_7_nl, FpIntToFloat_17U_5U_10U_o_expo_or_7_nl };
  assign _03467_ = _00011_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_6_nl, FpIntToFloat_17U_5U_10U_o_expo_or_6_nl, FpIntToFloat_17U_5U_10U_o_expo_or_6_nl, FpIntToFloat_17U_5U_10U_o_expo_or_6_nl, FpIntToFloat_17U_5U_10U_o_expo_or_6_nl };
  assign _03468_ = _00012_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_5_nl, FpIntToFloat_17U_5U_10U_o_expo_or_5_nl, FpIntToFloat_17U_5U_10U_o_expo_or_5_nl, FpIntToFloat_17U_5U_10U_o_expo_or_5_nl, FpIntToFloat_17U_5U_10U_o_expo_or_5_nl };
  assign _03469_ = _00013_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_4_nl, FpIntToFloat_17U_5U_10U_o_expo_or_4_nl, FpIntToFloat_17U_5U_10U_o_expo_or_4_nl, FpIntToFloat_17U_5U_10U_o_expo_or_4_nl, FpIntToFloat_17U_5U_10U_o_expo_or_4_nl };
  assign _03470_ = _00014_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_3_nl, FpIntToFloat_17U_5U_10U_o_expo_or_3_nl, FpIntToFloat_17U_5U_10U_o_expo_or_3_nl, FpIntToFloat_17U_5U_10U_o_expo_or_3_nl, FpIntToFloat_17U_5U_10U_o_expo_or_3_nl };
  assign _03471_ = _00015_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_2_nl, FpIntToFloat_17U_5U_10U_o_expo_or_2_nl, FpIntToFloat_17U_5U_10U_o_expo_or_2_nl, FpIntToFloat_17U_5U_10U_o_expo_or_2_nl, FpIntToFloat_17U_5U_10U_o_expo_or_2_nl };
  assign _03472_ = _00016_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_1_nl, FpIntToFloat_17U_5U_10U_o_expo_or_1_nl, FpIntToFloat_17U_5U_10U_o_expo_or_1_nl, FpIntToFloat_17U_5U_10U_o_expo_or_1_nl, FpIntToFloat_17U_5U_10U_o_expo_or_1_nl };
  assign _03473_ = _00017_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) { FpIntToFloat_17U_5U_10U_o_expo_or_nl, FpIntToFloat_17U_5U_10U_o_expo_or_nl, FpIntToFloat_17U_5U_10U_o_expo_or_nl, FpIntToFloat_17U_5U_10U_o_expo_or_nl, FpIntToFloat_17U_5U_10U_o_expo_or_nl };
  assign _03474_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2 };
  assign _03475_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2 };
  assign _03476_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2 };
  assign _03477_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2 };
  assign _03478_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2 };
  assign _03479_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2 };
  assign _03480_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2 };
  assign _03481_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2 };
  assign _03482_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2 };
  assign _03483_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2 };
  assign _03484_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2 };
  assign _03485_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2 };
  assign _03486_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2 };
  assign _03487_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1, cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1, cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1, cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1, cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1, cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1, cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1 };
  assign _03488_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2 };
  assign _03489_ = 6'b111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24394" *) { FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2, FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2 };
  assign _03490_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_1_nl, IntSaturation_17U_8U_and_1_nl, IntSaturation_17U_8U_and_1_nl, IntSaturation_17U_8U_and_1_nl, IntSaturation_17U_8U_and_1_nl, IntSaturation_17U_8U_and_1_nl, IntSaturation_17U_8U_and_1_nl };
  assign _03491_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_3_nl, IntSaturation_17U_8U_and_3_nl, IntSaturation_17U_8U_and_3_nl, IntSaturation_17U_8U_and_3_nl, IntSaturation_17U_8U_and_3_nl, IntSaturation_17U_8U_and_3_nl, IntSaturation_17U_8U_and_3_nl };
  assign _03492_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_5_nl, IntSaturation_17U_8U_and_5_nl, IntSaturation_17U_8U_and_5_nl, IntSaturation_17U_8U_and_5_nl, IntSaturation_17U_8U_and_5_nl, IntSaturation_17U_8U_and_5_nl, IntSaturation_17U_8U_and_5_nl };
  assign _03493_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_7_nl, IntSaturation_17U_8U_and_7_nl, IntSaturation_17U_8U_and_7_nl, IntSaturation_17U_8U_and_7_nl, IntSaturation_17U_8U_and_7_nl, IntSaturation_17U_8U_and_7_nl, IntSaturation_17U_8U_and_7_nl };
  assign _03494_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_9_nl, IntSaturation_17U_8U_and_9_nl, IntSaturation_17U_8U_and_9_nl, IntSaturation_17U_8U_and_9_nl, IntSaturation_17U_8U_and_9_nl, IntSaturation_17U_8U_and_9_nl, IntSaturation_17U_8U_and_9_nl };
  assign _03495_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_11_nl, IntSaturation_17U_8U_and_11_nl, IntSaturation_17U_8U_and_11_nl, IntSaturation_17U_8U_and_11_nl, IntSaturation_17U_8U_and_11_nl, IntSaturation_17U_8U_and_11_nl, IntSaturation_17U_8U_and_11_nl };
  assign _03496_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_13_nl, IntSaturation_17U_8U_and_13_nl, IntSaturation_17U_8U_and_13_nl, IntSaturation_17U_8U_and_13_nl, IntSaturation_17U_8U_and_13_nl, IntSaturation_17U_8U_and_13_nl, IntSaturation_17U_8U_and_13_nl };
  assign _03497_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_15_nl, IntSaturation_17U_8U_and_15_nl, IntSaturation_17U_8U_and_15_nl, IntSaturation_17U_8U_and_15_nl, IntSaturation_17U_8U_and_15_nl, IntSaturation_17U_8U_and_15_nl, IntSaturation_17U_8U_and_15_nl };
  assign _03498_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_17_nl, IntSaturation_17U_8U_and_17_nl, IntSaturation_17U_8U_and_17_nl, IntSaturation_17U_8U_and_17_nl, IntSaturation_17U_8U_and_17_nl, IntSaturation_17U_8U_and_17_nl, IntSaturation_17U_8U_and_17_nl };
  assign _03499_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_19_nl, IntSaturation_17U_8U_and_19_nl, IntSaturation_17U_8U_and_19_nl, IntSaturation_17U_8U_and_19_nl, IntSaturation_17U_8U_and_19_nl, IntSaturation_17U_8U_and_19_nl, IntSaturation_17U_8U_and_19_nl };
  assign _03500_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_21_nl, IntSaturation_17U_8U_and_21_nl, IntSaturation_17U_8U_and_21_nl, IntSaturation_17U_8U_and_21_nl, IntSaturation_17U_8U_and_21_nl, IntSaturation_17U_8U_and_21_nl, IntSaturation_17U_8U_and_21_nl };
  assign _03501_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_23_nl, IntSaturation_17U_8U_and_23_nl, IntSaturation_17U_8U_and_23_nl, IntSaturation_17U_8U_and_23_nl, IntSaturation_17U_8U_and_23_nl, IntSaturation_17U_8U_and_23_nl, IntSaturation_17U_8U_and_23_nl };
  assign _03502_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_25_nl, IntSaturation_17U_8U_and_25_nl, IntSaturation_17U_8U_and_25_nl, IntSaturation_17U_8U_and_25_nl, IntSaturation_17U_8U_and_25_nl, IntSaturation_17U_8U_and_25_nl, IntSaturation_17U_8U_and_25_nl };
  assign _03503_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_27_nl, IntSaturation_17U_8U_and_27_nl, IntSaturation_17U_8U_and_27_nl, IntSaturation_17U_8U_and_27_nl, IntSaturation_17U_8U_and_27_nl, IntSaturation_17U_8U_and_27_nl, IntSaturation_17U_8U_and_27_nl };
  assign _03504_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_29_nl, IntSaturation_17U_8U_and_29_nl, IntSaturation_17U_8U_and_29_nl, IntSaturation_17U_8U_and_29_nl, IntSaturation_17U_8U_and_29_nl, IntSaturation_17U_8U_and_29_nl, IntSaturation_17U_8U_and_29_nl };
  assign _03505_ = 7'b1000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) { IntSaturation_17U_8U_and_31_nl, IntSaturation_17U_8U_and_31_nl, IntSaturation_17U_8U_and_31_nl, IntSaturation_17U_8U_and_31_nl, IntSaturation_17U_8U_and_31_nl, IntSaturation_17U_8U_and_31_nl, IntSaturation_17U_8U_and_31_nl };
  assign _03506_ = reg_chn_idata_data_sva_3_15_0_2_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl };
  assign _03507_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl };
  assign _03508_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl };
  assign _03509_ = FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl };
  assign _03510_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl };
  assign _03511_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl };
  assign _03512_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl };
  assign _03513_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl };
  assign _03514_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl };
  assign _03515_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl };
  assign _03516_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl };
  assign _03517_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl };
  assign _03518_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl };
  assign _03519_ = reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl };
  assign _03520_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl };
  assign { _03846_[6:2], _03521_ } = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[6:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl, IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl };
  assign _03522_ = { IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24408" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03523_ = FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24409" *) { cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323 };
  assign _03524_ = reg_chn_idata_data_sva_3_15_0_2_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24410" *) { cvt_or_48_nl, cvt_or_48_nl, cvt_or_48_nl, cvt_or_48_nl, cvt_or_48_nl, cvt_or_48_nl, cvt_or_48_nl, cvt_or_48_nl, cvt_or_48_nl };
  assign _03525_ = reg_chn_idata_data_sva_3_15_0_2_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24411" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03526_ = { IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_333, cvt_asn_333, cvt_asn_333, cvt_asn_333, cvt_asn_333, cvt_asn_333, cvt_asn_333, cvt_asn_333, cvt_asn_333 };
  assign _03527_ = { IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03528_ = { IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_339, cvt_asn_339, cvt_asn_339, cvt_asn_339, cvt_asn_339, cvt_asn_339, cvt_asn_339, cvt_asn_339, cvt_asn_339 };
  assign _03529_ = { IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03530_ = { IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_357, cvt_asn_357, cvt_asn_357, cvt_asn_357, cvt_asn_357, cvt_asn_357, cvt_asn_357, cvt_asn_357, cvt_asn_357 };
  assign _03531_ = { IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_369, cvt_asn_369, cvt_asn_369, cvt_asn_369, cvt_asn_369, cvt_asn_369, cvt_asn_369, cvt_asn_369, cvt_asn_369 };
  assign _03532_ = { IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_381, cvt_asn_381, cvt_asn_381, cvt_asn_381, cvt_asn_381, cvt_asn_381, cvt_asn_381, cvt_asn_381, cvt_asn_381 };
  assign _03533_ = { IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327, cvt_asn_327 };
  assign _03534_ = { IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_399, cvt_asn_399, cvt_asn_399, cvt_asn_399, cvt_asn_399, cvt_asn_399, cvt_asn_399, cvt_asn_399, cvt_asn_399 };
  assign _03535_ = { IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_393, cvt_asn_393, cvt_asn_393, cvt_asn_393, cvt_asn_393, cvt_asn_393, cvt_asn_393, cvt_asn_393, cvt_asn_393 };
  assign _03536_ = { IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_387, cvt_asn_387, cvt_asn_387, cvt_asn_387, cvt_asn_387, cvt_asn_387, cvt_asn_387, cvt_asn_387, cvt_asn_387 };
  assign _03537_ = { IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_375, cvt_asn_375, cvt_asn_375, cvt_asn_375, cvt_asn_375, cvt_asn_375, cvt_asn_375, cvt_asn_375, cvt_asn_375 };
  assign _03538_ = { IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_363, cvt_asn_363, cvt_asn_363, cvt_asn_363, cvt_asn_363, cvt_asn_363, cvt_asn_363, cvt_asn_363, cvt_asn_363 };
  assign _03539_ = { IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cvt_asn_351, cvt_asn_351, cvt_asn_351, cvt_asn_351, cvt_asn_351, cvt_asn_351, cvt_asn_351, cvt_asn_351, cvt_asn_351 };
  assign _03540_ = chn_idata_data_sva_3_495_479_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24424" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03541_ = FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_329, cvt_asn_329, cvt_asn_329, cvt_asn_329, cvt_asn_329, cvt_asn_329, cvt_asn_329, cvt_asn_329, cvt_asn_329 };
  assign _03542_ = FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323 };
  assign _03543_ = FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_335, cvt_asn_335, cvt_asn_335, cvt_asn_335, cvt_asn_335, cvt_asn_335, cvt_asn_335, cvt_asn_335, cvt_asn_335 };
  assign _03544_ = FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323 };
  assign _03545_ = FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_353, cvt_asn_353, cvt_asn_353, cvt_asn_353, cvt_asn_353, cvt_asn_353, cvt_asn_353, cvt_asn_353, cvt_asn_353 };
  assign _03546_ = FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_365, cvt_asn_365, cvt_asn_365, cvt_asn_365, cvt_asn_365, cvt_asn_365, cvt_asn_365, cvt_asn_365, cvt_asn_365 };
  assign _03547_ = FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_377, cvt_asn_377, cvt_asn_377, cvt_asn_377, cvt_asn_377, cvt_asn_377, cvt_asn_377, cvt_asn_377, cvt_asn_377 };
  assign _03548_ = FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323, cvt_asn_323 };
  assign _03549_ = FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371 };
  assign _03550_ = FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_389, cvt_asn_389, cvt_asn_389, cvt_asn_389, cvt_asn_389, cvt_asn_389, cvt_asn_389, cvt_asn_389, cvt_asn_389 };
  assign _03551_ = FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_383, cvt_asn_383, cvt_asn_383, cvt_asn_383, cvt_asn_383, cvt_asn_383, cvt_asn_383, cvt_asn_383, cvt_asn_383 };
  assign _03552_ = FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371, cvt_asn_371 };
  assign _03553_ = FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_359, cvt_asn_359, cvt_asn_359, cvt_asn_359, cvt_asn_359, cvt_asn_359, cvt_asn_359, cvt_asn_359, cvt_asn_359 };
  assign _03554_ = FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_347, cvt_asn_347, cvt_asn_347, cvt_asn_347, cvt_asn_347, cvt_asn_347, cvt_asn_347, cvt_asn_347, cvt_asn_347 };
  assign _03555_ = { IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6], IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) { cvt_asn_345, cvt_asn_345, cvt_asn_345, cvt_asn_345, cvt_asn_345, cvt_asn_345, cvt_asn_345, cvt_asn_345, cvt_asn_345 };
  assign _03556_ = chn_idata_data_sva_3_47_31_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03557_ = chn_idata_data_sva_3_79_63_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03558_ = chn_idata_data_sva_3_111_95_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03559_ = chn_idata_data_sva_3_143_127_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03560_ = chn_idata_data_sva_3_175_159_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03561_ = chn_idata_data_sva_3_207_191_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03562_ = chn_idata_data_sva_3_239_223_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03563_ = chn_idata_data_sva_3_271_255_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03564_ = chn_idata_data_sva_3_303_287_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03565_ = chn_idata_data_sva_3_335_319_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03566_ = chn_idata_data_sva_3_367_351_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03567_ = chn_idata_data_sva_3_399_383_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03568_ = chn_idata_data_sva_3_431_415_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03569_ = chn_idata_data_sva_3_463_447_1[10:2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6, cfg_mode_eql_1_sva_6 };
  assign _03570_ = FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) { cvt_asn_341, cvt_asn_341, cvt_asn_341, cvt_asn_341, cvt_asn_341, cvt_asn_341, cvt_asn_341, cvt_asn_341, cvt_asn_341 };
  assign _03571_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03572_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03573_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03574_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03575_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03576_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03577_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03578_ = FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03579_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03580_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03581_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03582_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03583_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03584_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03585_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[9:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) { cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321, cvt_asn_321 };
  assign _03586_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse, cvt_or_2_cse };
  assign _03587_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03588_ = FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_6_cse, cvt_or_6_cse, cvt_or_6_cse, cvt_or_6_cse, cvt_or_6_cse, cvt_or_6_cse, cvt_or_6_cse, cvt_or_6_cse, cvt_or_6_cse };
  assign _03589_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03590_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse, cvt_or_10_cse };
  assign _03591_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse, cvt_or_12_cse };
  assign _03592_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_14_cse, cvt_or_14_cse, cvt_or_14_cse, cvt_or_14_cse, cvt_or_14_cse, cvt_or_14_cse, cvt_or_14_cse, cvt_or_14_cse, cvt_or_14_cse };
  assign _03593_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse, cvt_or_cse };
  assign _03594_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse, cvt_or_18_cse };
  assign _03595_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse, cvt_or_20_cse };
  assign _03596_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_22_cse, cvt_or_22_cse, cvt_or_22_cse, cvt_or_22_cse, cvt_or_22_cse, cvt_or_22_cse, cvt_or_22_cse, cvt_or_22_cse, cvt_or_22_cse };
  assign _03597_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse, cvt_or_24_cse };
  assign _03598_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_26_cse, cvt_or_26_cse, cvt_or_26_cse, cvt_or_26_cse, cvt_or_26_cse, cvt_or_26_cse, cvt_or_26_cse, cvt_or_26_cse, cvt_or_26_cse };
  assign _03599_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse, cvt_or_28_cse };
  assign _03600_ = reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[8:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) { cvt_or_30_cse, cvt_or_30_cse, cvt_or_30_cse, cvt_or_30_cse, cvt_or_30_cse, cvt_or_30_cse, cvt_or_30_cse, cvt_or_30_cse, cvt_or_30_cse };
  assign _03601_ = cvt_else_equal_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8773" *) _04517_;
  assign _03602_ = _03601_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8773" *) cvt_unequal_tmp_21;
  assign chn_out_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8774" *) _05299_;
  assign _03603_ = _09452_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8777" *) or_5189_cse;
  assign and_3024_cse = _03603_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8777" *) and_dcpl_1742;
  assign _03604_ = cvt_else_equal_tmp_3_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8779" *) _04517_;
  assign _03605_ = _03604_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8779" *) cvt_unequal_tmp_21;
  assign _03606_ = cvt_else_equal_tmp_9_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8781" *) _04517_;
  assign _03607_ = _03606_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8781" *) cvt_unequal_tmp_21;
  assign _03608_ = cvt_else_equal_tmp_15_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8783" *) _04517_;
  assign _03609_ = _03608_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8783" *) cvt_unequal_tmp_21;
  assign _03610_ = cvt_else_equal_tmp_18_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8785" *) _04517_;
  assign _03611_ = _03610_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8785" *) cvt_unequal_tmp_21;
  assign _03612_ = cvt_else_equal_tmp_21_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8786" *) cvt_and_147_m1c;
  assign _03613_ = cvt_else_equal_tmp_27_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8788" *) _04517_;
  assign _03614_ = _03613_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8788" *) cvt_unequal_tmp_21;
  assign _03615_ = cvt_else_equal_tmp_30_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8790" *) _04517_;
  assign _03616_ = _03615_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8790" *) cvt_unequal_tmp_21;
  assign _03617_ = cvt_else_equal_tmp_33_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8792" *) _04517_;
  assign _03618_ = _03617_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8792" *) cvt_unequal_tmp_21;
  assign _03619_ = cvt_else_equal_tmp_36_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8794" *) _04517_;
  assign _03620_ = _03619_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8794" *) cvt_unequal_tmp_21;
  assign _03621_ = cvt_else_equal_tmp_39_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8796" *) _04517_;
  assign _03622_ = _03621_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8796" *) cvt_unequal_tmp_21;
  assign _03623_ = _09454_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8800" *) or_5189_cse;
  assign and_3063_cse = _03623_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8800" *) and_dcpl_1742;
  assign _03624_ = cvt_else_equal_tmp_42_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8802" *) _04517_;
  assign _03625_ = _03624_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8802" *) cvt_unequal_tmp_21;
  assign _03626_ = cvt_else_equal_tmp_39_mx1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8805" *) cvt_unequal_tmp_21;
  assign _03627_ = _03626_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8805" *) _04517_;
  assign _03628_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8806" *) cvt_unequal_tmp_21;
  assign _03629_ = _03628_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8807" *) or_5189_cse;
  assign chn_out_and_32_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8807" *) _09455_;
  assign _03630_ = cfg_mode_eql_1_sva_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8809" *) main_stage_v_3;
  assign _03631_ = _03630_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8809" *) or_5189_cse;
  assign chn_out_and_77_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8809" *) _09456_;
  assign and_2239_cse = cfg_mode_eql_1_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8811" *) main_stage_v_1;
  assign IntShiftRightSat_49U_6U_17U_o_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8813" *) _04174_;
  assign chn_idata_data_and_1_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8813" *) mux_12_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8816" *) _04957_;
  assign IntMulExt_33U_16U_49U_and_11_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8817" *) mux_133_cse;
  assign IntMulExt_33U_16U_49U_and_1_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8818" *) _09457_;
  assign cfg_proc_precision_and_11_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8819" *) mux_tmp_114;
  assign chn_idata_data_and_16_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8820" *) mux_tmp_161;
  assign and_637_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8821" *) _05301_;
  assign _03632_ = cfg_proc_precision_1_sva_st_65[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8822" *) cfg_out_precision_1_sva_st_149[0];
  assign and_639_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8825" *) _05302_;
  assign FpFloatToInt_16U_5U_10U_shift_and_1_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8829" *) mux_163_nl;
  assign and_641_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8830" *) _05303_;
  assign and_643_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8831" *) _05304_;
  assign and_646_rgt = or_tmp_2469 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8833" *) or_5189_cse;
  assign and_648_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8841" *) _05305_;
  assign FpFloatToInt_16U_5U_10U_shift_and_5_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8845" *) _05306_;
  assign and_650_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8846" *) _05307_;
  assign and_652_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8847" *) _05308_;
  assign and_654_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8848" *) _05309_;
  assign and_656_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8853" *) _05310_;
  assign and_658_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8854" *) _05311_;
  assign and_660_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8855" *) _05312_;
  assign and_662_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8856" *) _05313_;
  assign and_664_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8857" *) _05314_;
  assign and_666_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8858" *) _05315_;
  assign and_668_rgt = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8859" *) _05316_;
  assign and_2237_cse = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8864" *) or_4862_cse;
  assign _03633_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8871" *) _05318_;
  assign _03634_ = _03633_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8872" *) _05431_;
  assign _03635_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8872" *) _09461_;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_cse = _03635_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8873" *) _04856_;
  assign _03636_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8882" *) _05319_;
  assign _03637_ = _03636_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8883" *) _05435_;
  assign _03638_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8883" *) _09463_;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_13_cse = _03638_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8884" *) not_tmp_249;
  assign IntShiftRightSat_49U_6U_17U_if_and_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8890" *) mux_273_nl;
  assign and_685_rgt = or_dcpl_15 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8891" *) or_5189_cse;
  assign _03639_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8893" *) _05320_;
  assign _03640_ = _03639_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8894" *) _05439_;
  assign _03641_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8895" *) _09465_;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_15_cse = _03641_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8895" *) not_tmp_269;
  assign _03642_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8899" *) and_dcpl_228;
  assign _03643_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8900" *) _04857_;
  assign and_696_nl = _03643_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8900" *) or_dcpl_108;
  assign _03644_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8901" *) or_dcpl_109;
  assign and_699_nl = _03644_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8901" *) and_dcpl_228;
  assign and_2257_cse = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8910" *) core_wen;
  assign and_2259_cse = _04862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8917" *) core_wen;
  assign and_704_rgt = or_dcpl_109 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8918" *) or_5189_cse;
  assign and_2230_cse = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8919" *) mux_1126_cse;
  assign _03645_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8921" *) _04859_;
  assign and_711_nl = _03645_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8921" *) or_dcpl_110;
  assign _03646_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8922" *) or_dcpl_111;
  assign and_714_nl = _03646_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8922" *) and_dcpl_228;
  assign and_719_rgt = or_dcpl_111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8930" *) or_5189_cse;
  assign and_174_cse = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8934" *) mux_382_cse;
  assign _03647_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8939" *) _04860_;
  assign and_726_nl = _03647_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8939" *) or_dcpl_113;
  assign _03648_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8940" *) or_dcpl_114;
  assign and_729_nl = _03648_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8940" *) and_dcpl_228;
  assign and_2275_cse = _05321_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8947" *) core_wen;
  assign and_734_rgt = or_dcpl_114 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8948" *) or_5189_cse;
  assign and_178_itm = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8949" *) and_tmp_79;
  assign IntShiftRightSat_49U_6U_17U_if_and_3_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8952" *) mux_378_nl;
  assign _03649_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8957" *) _04861_;
  assign and_741_nl = _03649_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8957" *) or_dcpl_115;
  assign _03650_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8958" *) or_dcpl_116;
  assign and_744_nl = _03650_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8958" *) and_dcpl_228;
  assign and_749_rgt = or_dcpl_116 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8962" *) or_5189_cse;
  assign _03651_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8968" *) _04863_;
  assign and_756_nl = _03651_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8968" *) or_dcpl_119;
  assign _03652_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8969" *) or_dcpl_120;
  assign and_759_nl = _03652_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8969" *) and_dcpl_228;
  assign and_766_rgt = or_dcpl_120 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8974" *) or_5189_cse;
  assign _03653_ = or_5189_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8976" *) _05324_;
  assign _03654_ = _03653_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8977" *) _05450_;
  assign _03655_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8977" *) _09475_;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_22_cse = _03655_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8978" *) not_tmp_520;
  assign _03656_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8984" *) _04864_;
  assign and_780_nl = _03656_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8984" *) or_dcpl_124;
  assign _03657_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8985" *) or_dcpl_125;
  assign and_783_nl = _03657_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8985" *) and_dcpl_228;
  assign and_787_rgt = or_dcpl_125 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8990" *) or_5189_cse;
  assign _03658_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8992" *) _04865_;
  assign and_794_nl = _03658_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8992" *) or_dcpl_126;
  assign _03659_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8993" *) or_dcpl_127;
  assign and_797_nl = _03659_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8993" *) and_dcpl_228;
  assign and_801_rgt = or_dcpl_127 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8998" *) or_5189_cse;
  assign _03660_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9001" *) _04866_;
  assign and_808_nl = _03660_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9001" *) or_dcpl_130;
  assign _03661_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9002" *) or_dcpl_131;
  assign and_811_nl = _03661_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9002" *) and_dcpl_228;
  assign and_2317_cse = _05327_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9011" *) core_wen;
  assign and_816_rgt = or_dcpl_131 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9012" *) or_5189_cse;
  assign _03662_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9014" *) _04868_;
  assign and_823_nl = _03662_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9014" *) or_dcpl_132;
  assign _03663_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9015" *) or_dcpl_133;
  assign and_826_nl = _03663_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9015" *) and_dcpl_228;
  assign _03664_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9016" *) _05328_;
  assign and_830_rgt = or_dcpl_133 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9022" *) or_5189_cse;
  assign IntShiftRightSat_49U_6U_17U_o_and_90_cse = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9024" *) mux_tmp_161;
  assign _03665_ = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9032" *) _03980_;
  assign _03666_ = _03665_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9032" *) mux_1142_cse;
  assign _03667_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9038" *) and_dcpl_363;
  assign _03668_ = _03667_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9038" *) or_dcpl_136;
  assign and_840_nl = _03668_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9038" *) _04869_;
  assign and_843_nl = _03667_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9039" *) or_dcpl_137;
  assign and_849_rgt = or_dcpl_137 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9044" *) or_5189_cse;
  assign _03669_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9048" *) _04871_;
  assign and_856_nl = _03669_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9048" *) or_dcpl_139;
  assign _03670_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9049" *) or_dcpl_140;
  assign and_859_nl = _03670_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9049" *) and_dcpl_228;
  assign _03671_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9051" *) and_tmp_225;
  assign and_866_rgt = or_dcpl_140 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9057" *) or_5189_cse;
  assign _03672_ = _03642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9059" *) _04873_;
  assign and_873_nl = _03672_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9059" *) or_dcpl_143;
  assign _03673_ = and_676_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9060" *) or_dcpl_144;
  assign and_876_nl = _03673_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9060" *) and_dcpl_228;
  assign and_881_rgt = or_dcpl_144 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9070" *) or_5189_cse;
  assign cfg_proc_precision_and_24_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9077" *) mux_796_nl;
  assign cfg_proc_precision_and_27_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9079" *) mux_800_nl;
  assign FpFloatToInt_16U_5U_10U_internal_int_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9081" *) _09486_;
  assign and_896_rgt = _09492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9090" *) and_dcpl_408;
  assign _03674_ = nor_1056_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9091" *) cfg_proc_precision_1_sva_st_65[1];
  assign and_900_rgt = _03674_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9091" *) and_dcpl_417;
  assign FpFloatToInt_16U_5U_10U_if_and_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9102" *) mux_818_nl;
  assign _03675_ = nor_50_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9103" *) or_5189_cse;
  assign _03676_ = cfg_out_precision_1_sva_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9107" *) or_1159_cse;
  assign _03677_ = _05332_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9121" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c;
  assign FpFloatToInt_16U_5U_10U_and_33_nl = _03677_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9121" *) and_dcpl_433;
  assign _03678_ = chn_idata_data_sva_2_79_63_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9123" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c;
  assign FpFloatToInt_16U_5U_10U_and_34_nl = _03678_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9123" *) and_dcpl_433;
  assign _03679_ = cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9125" *) _05333_;
  assign FpFloatToInt_16U_5U_10U_and_3_nl = _03679_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9125" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_nl = IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9127" *) and_dcpl_433;
  assign and_916_nl = _09498_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9128" *) and_dcpl_420;
  assign _03680_ = and_tmp_50 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9129" *) _04000_;
  assign _03681_ = _03680_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9130" *) cvt_unequal_tmp_20;
  assign and_921_nl = _03681_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9130" *) or_5189_cse;
  assign _03682_ = _05334_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9152" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c;
  assign FpFloatToInt_16U_5U_10U_and_35_nl = _03682_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9152" *) and_dcpl_433;
  assign _03683_ = chn_idata_data_sva_2_111_95_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9154" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c;
  assign FpFloatToInt_16U_5U_10U_and_36_nl = _03683_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9154" *) and_dcpl_433;
  assign _03684_ = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9156" *) _05335_;
  assign FpFloatToInt_16U_5U_10U_and_5_nl = _03684_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9156" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_29_nl = IsNaN_5U_10U_land_3_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9158" *) and_dcpl_433;
  assign _03685_ = cfg_proc_precision_1_sva_st_65[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9167" *) cvt_unequal_tmp_20;
  assign _03686_ = mux_2226_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9172" *) or_5189_cse;
  assign and_2365_cse = _03686_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9172" *) core_wen;
  assign _03687_ = _09504_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9174" *) or_5189_cse;
  assign and_2369_cse = _03687_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9174" *) core_wen;
  assign _03688_ = _05338_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9184" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c;
  assign FpFloatToInt_16U_5U_10U_and_61_nl = _03688_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9184" *) and_dcpl_433;
  assign _03689_ = chn_idata_data_sva_2_511_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9186" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c;
  assign FpFloatToInt_16U_5U_10U_and_62_nl = _03689_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9186" *) and_dcpl_433;
  assign _03690_ = cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9188" *) _05339_;
  assign FpFloatToInt_16U_5U_10U_and_31_nl = _03690_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9188" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_27_nl = IsNaN_5U_10U_land_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9190" *) and_dcpl_433;
  assign and_945_nl = _09510_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9191" *) and_dcpl_420;
  assign _03691_ = mux_tmp_1813 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9192" *) or_5189_cse;
  assign and_949_nl = _03691_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9192" *) and_dcpl_458;
  assign and_2371_nl = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9200" *) _09509_;
  assign _03692_ = mux_2227_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9202" *) or_5189_cse;
  assign and_2372_cse = _03692_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9202" *) core_wen;
  assign _01995_ = or_4714_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9203" *) _03931_;
  assign _03693_ = _01995_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *) or_400_cse_1;
  assign _03694_ = _09512_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *) or_5189_cse;
  assign and_2380_cse = _03694_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *) core_wen;
  assign and_2156_nl = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9205" *) nor_2285_cse;
  assign and_954_rgt = mux_1859_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9207" *) and_dcpl_408;
  assign _03695_ = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9209" *) cfg_proc_precision_1_sva_st_65[1];
  assign and_956_rgt = _03695_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9209" *) and_dcpl_417;
  assign _03696_ = _05139_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9213" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c;
  assign FpFloatToInt_16U_5U_10U_and_39_nl = _03696_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9213" *) and_dcpl_433;
  assign _03697_ = chn_idata_data_sva_2_175_159_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9215" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c;
  assign FpFloatToInt_16U_5U_10U_and_40_nl = _03697_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9215" *) and_dcpl_433;
  assign _03698_ = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9217" *) _05340_;
  assign FpFloatToInt_16U_5U_10U_and_9_nl = _03698_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9217" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_26_nl = IsNaN_5U_10U_land_5_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9219" *) and_dcpl_433;
  assign and_957_rgt = or_dcpl_147 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9232" *) or_5189_cse;
  assign _03699_ = _05148_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9239" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c;
  assign FpFloatToInt_16U_5U_10U_and_59_nl = _03699_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9239" *) and_dcpl_433;
  assign _03700_ = chn_idata_data_sva_2_495_479_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9241" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c;
  assign FpFloatToInt_16U_5U_10U_and_60_nl = _03700_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9241" *) and_dcpl_433;
  assign _03701_ = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9243" *) _05341_;
  assign FpFloatToInt_16U_5U_10U_and_29_nl = _03701_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9243" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_25_nl = IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9245" *) and_dcpl_433;
  assign and_961_nl = _09522_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9246" *) and_dcpl_420;
  assign _03702_ = and_dcpl_473 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9247" *) _04947_;
  assign _03703_ = _03702_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9248" *) _04691_;
  assign and_966_nl = _03703_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9248" *) cvt_unequal_tmp_20;
  assign and_2388_cse = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9261" *) or_4749_cse;
  assign _03704_ = mux_2231_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9263" *) or_5189_cse;
  assign and_2389_cse = _03704_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9263" *) core_wen;
  assign _03705_ = _09523_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9266" *) or_5189_cse;
  assign and_2393_cse = _03705_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9266" *) core_wen;
  assign and_1013_nl = _09524_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9268" *) and_dcpl_420;
  assign and_978_cse = and_tmp_225 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9269" *) and_dcpl_481;
  assign _03706_ = _05343_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9277" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c;
  assign FpFloatToInt_16U_5U_10U_and_41_nl = _03706_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9277" *) and_dcpl_433;
  assign _03707_ = chn_idata_data_sva_2_207_191_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9279" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c;
  assign FpFloatToInt_16U_5U_10U_and_42_nl = _03707_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9279" *) and_dcpl_433;
  assign _03708_ = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9281" *) _05344_;
  assign FpFloatToInt_16U_5U_10U_and_11_nl = _03708_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9281" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_24_nl = IsNaN_5U_10U_land_6_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9283" *) and_dcpl_433;
  assign _03709_ = or_4714_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *) _05345_;
  assign and_2395_nl = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *) _05346_;
  assign _03710_ = mux_2233_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9292" *) or_5189_cse;
  assign and_2396_cse = _03710_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9292" *) core_wen;
  assign _03711_ = or_400_cse_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9293" *) cfg_out_precision_1_sva_st_113[1];
  assign _03712_ = _03711_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *) _05347_;
  assign _03713_ = _09531_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9295" *) or_5189_cse;
  assign and_2402_cse = _03713_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9295" *) core_wen;
  assign and_2154_nl = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9296" *) nor_45_cse;
  assign and_984_rgt = mux_1886_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9298" *) and_dcpl_408;
  assign _03714_ = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9300" *) cfg_proc_precision_1_sva_st_65[1];
  assign and_986_rgt = _03714_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9300" *) and_dcpl_417;
  assign _03715_ = _05348_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9302" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c;
  assign FpFloatToInt_16U_5U_10U_and_57_nl = _03715_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9302" *) and_dcpl_433;
  assign _03716_ = chn_idata_data_sva_2_463_447_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9304" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c;
  assign FpFloatToInt_16U_5U_10U_and_58_nl = _03716_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9304" *) and_dcpl_433;
  assign _03717_ = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9306" *) _05349_;
  assign FpFloatToInt_16U_5U_10U_and_27_nl = _03717_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9306" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_23_nl = IsNaN_5U_10U_land_14_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9308" *) and_dcpl_433;
  assign and_2153_nl = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9320" *) nor_45_cse;
  assign and_987_rgt = mux_1892_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9322" *) and_dcpl_408;
  assign _03718_ = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9324" *) cfg_proc_precision_1_sva_st_65[1];
  assign and_989_rgt = _03718_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9324" *) and_dcpl_417;
  assign _03719_ = _05153_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9329" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c;
  assign FpFloatToInt_16U_5U_10U_and_43_nl = _03719_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9329" *) and_dcpl_433;
  assign _03720_ = chn_idata_data_sva_2_239_223_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9331" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c;
  assign FpFloatToInt_16U_5U_10U_and_44_nl = _03720_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9331" *) and_dcpl_433;
  assign _03721_ = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9333" *) _05350_;
  assign FpFloatToInt_16U_5U_10U_and_13_nl = _03721_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9333" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_22_nl = IsNaN_5U_10U_land_7_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9335" *) and_dcpl_433;
  assign _03722_ = _05351_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9346" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c;
  assign FpFloatToInt_16U_5U_10U_and_55_nl = _03722_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9346" *) and_dcpl_433;
  assign _03723_ = chn_idata_data_sva_2_431_415_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9348" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c;
  assign FpFloatToInt_16U_5U_10U_and_56_nl = _03723_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9348" *) and_dcpl_433;
  assign _03724_ = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9350" *) _05352_;
  assign FpFloatToInt_16U_5U_10U_and_25_nl = _03724_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9350" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_21_nl = IsNaN_5U_10U_land_13_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9352" *) and_dcpl_433;
  assign and_999_nl = _09534_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9353" *) and_dcpl_420;
  assign _03725_ = and_dcpl_499 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9354" *) _04947_;
  assign _03726_ = _03725_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9355" *) _04691_;
  assign _03727_ = _03726_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9355" *) cvt_unequal_tmp_20;
  assign and_1004_nl = _03727_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9355" *) or_400_cse_1;
  assign _03728_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9367" *) mux_2236_nl;
  assign and_2422_cse = cvt_unequal_tmp_20 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9368" *) or_4788_cse;
  assign and_2151_nl = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9369" *) nor_45_cse;
  assign and_1009_rgt = mux_1916_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9371" *) and_dcpl_408;
  assign _03729_ = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9373" *) cfg_proc_precision_1_sva_st_65[1];
  assign and_1011_rgt = _03729_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9373" *) and_dcpl_417;
  assign _03730_ = _05173_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9377" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c;
  assign FpFloatToInt_16U_5U_10U_and_45_nl = _03730_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9377" *) and_dcpl_433;
  assign _03731_ = chn_idata_data_sva_2_271_255_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9379" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c;
  assign FpFloatToInt_16U_5U_10U_and_46_nl = _03731_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9379" *) and_dcpl_433;
  assign _03732_ = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9381" *) _05354_;
  assign FpFloatToInt_16U_5U_10U_and_15_nl = _03732_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9381" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_20_nl = IsNaN_5U_10U_land_8_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9383" *) and_dcpl_433;
  assign _03733_ = _05355_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9395" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c;
  assign FpFloatToInt_16U_5U_10U_and_53_nl = _03733_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9395" *) and_dcpl_433;
  assign _03734_ = chn_idata_data_sva_2_399_383_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9397" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c;
  assign FpFloatToInt_16U_5U_10U_and_54_nl = _03734_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9397" *) and_dcpl_433;
  assign _03735_ = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9399" *) _05356_;
  assign FpFloatToInt_16U_5U_10U_and_23_nl = _03735_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9399" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_19_nl = IsNaN_5U_10U_land_12_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9401" *) and_dcpl_433;
  assign and_1023_nl = _09536_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9402" *) and_dcpl_420;
  assign _03736_ = and_3372_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9404" *) _04691_;
  assign _03737_ = _03736_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9404" *) cvt_unequal_tmp_20;
  assign and_1027_nl = _03737_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9404" *) or_5189_cse;
  assign and_2149_nl = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9405" *) nor_1048_cse;
  assign _03738_ = _05357_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9424" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c;
  assign FpFloatToInt_16U_5U_10U_and_47_nl = _03738_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9424" *) and_dcpl_433;
  assign _03739_ = chn_idata_data_sva_2_303_287_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9426" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c;
  assign FpFloatToInt_16U_5U_10U_and_48_nl = _03739_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9426" *) and_dcpl_433;
  assign _03740_ = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9428" *) _05358_;
  assign FpFloatToInt_16U_5U_10U_and_17_nl = _03740_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9428" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_18_nl = IsNaN_5U_10U_land_9_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9430" *) and_dcpl_433;
  assign and_1039_cse = mux_1142_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9440" *) and_dcpl_481;
  assign _03741_ = _05359_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9444" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c;
  assign FpFloatToInt_16U_5U_10U_and_51_nl = _03741_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9444" *) and_dcpl_433;
  assign _03742_ = chn_idata_data_sva_2_367_351_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9446" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c;
  assign FpFloatToInt_16U_5U_10U_and_52_nl = _03742_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9446" *) and_dcpl_433;
  assign _03743_ = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9448" *) _05360_;
  assign FpFloatToInt_16U_5U_10U_and_21_nl = _03743_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9448" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_17_nl = IsNaN_5U_10U_land_11_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9450" *) and_dcpl_433;
  assign _03744_ = _05361_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9461" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c;
  assign FpFloatToInt_16U_5U_10U_and_49_nl = _03744_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9461" *) and_dcpl_433;
  assign _03745_ = chn_idata_data_sva_2_335_319_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9463" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c;
  assign FpFloatToInt_16U_5U_10U_and_50_nl = _03745_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9463" *) and_dcpl_433;
  assign _03746_ = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9465" *) _05362_;
  assign FpFloatToInt_16U_5U_10U_and_19_nl = _03746_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9465" *) and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_16_nl = IsNaN_5U_10U_land_10_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9467" *) and_dcpl_433;
  assign cfg_out_precision_and_32_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9476" *) mux_938_nl;
  assign cvt_else_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9479" *) _05363_;
  assign _03747_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9482" *) _05364_;
  assign cvt_else_and_24_cse = _03747_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9482" *) _05365_;
  assign cvt_else_and_10_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9485" *) reg_cvt_else_cvt_else_nor_4_cse;
  assign _03748_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *) _05366_;
  assign cvt_else_and_34_cse = _03748_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *) _05367_;
  assign cvt_else_and_19_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9495" *) _05368_;
  assign IntShiftRightSat_49U_6U_17U_o_and_103_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9505" *) mux_1003_nl;
  assign _03749_ = cvt_1_FpMantRNE_17U_11U_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9507" *) cvt_unequal_tmp_20;
  assign and_1069_m1c = _03749_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9507" *) or_5189_cse;
  assign _03750_ = _04898_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9512" *) and_1069_m1c;
  assign _03751_ = _05128_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9513" *) cvt_unequal_tmp_20;
  assign _03752_ = _03751_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9513" *) or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_31_nl = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9515" *) and_1069_m1c;
  assign and_1078_cse = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9524" *) and_tmp_50;
  assign _03753_ = _07889_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9525" *) or_1159_cse;
  assign _03754_ = _03753_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9526" *) or_3538_cse;
  assign and_1077_rgt = _03754_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9526" *) and_dcpl_103;
  assign and_1080_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9527" *) cvt_2_FpMantRNE_17U_11U_else_and_1_tmp;
  assign _03755_ = _05200_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9533" *) and_1080_m1c;
  assign _03756_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9533" *) _05369_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_29_nl = cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9535" *) and_1080_m1c;
  assign FpIntToFloat_17U_5U_10U_is_inf_and_14_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9547" *) mux_1027_nl;
  assign and_1084_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9548" *) cvt_3_FpMantRNE_17U_11U_else_and_1_tmp;
  assign _03757_ = _04907_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9554" *) and_1084_m1c;
  assign _03758_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9554" *) _05370_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_27_nl = cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9556" *) and_1084_m1c;
  assign and_2186_cse = or_4524_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9566" *) chn_in_rsci_bawt;
  assign _03759_ = _09561_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9569" *) or_1159_cse;
  assign _03760_ = _03759_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9569" *) or_3538_cse;
  assign _03761_ = _03760_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9569" *) or_3542_cse;
  assign and_1091_rgt = _03761_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9569" *) and_dcpl_103;
  assign _03762_ = cvt_4_FpMantRNE_17U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9575" *) cvt_unequal_tmp_20;
  assign and_1093_m1c = _03762_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9575" *) or_5189_cse;
  assign _03763_ = _04287_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9581" *) and_1093_m1c;
  assign _03764_ = _05371_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9582" *) cvt_unequal_tmp_20;
  assign _03765_ = _03764_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9582" *) or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_25_nl = cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9584" *) and_1093_m1c;
  assign and_1097_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9589" *) cvt_5_FpMantRNE_17U_11U_else_and_1_tmp;
  assign _03766_ = _04910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9595" *) and_1097_m1c;
  assign _03767_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9595" *) _05372_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_23_nl = cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9597" *) and_1097_m1c;
  assign _03768_ = _07928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9603" *) or_1159_cse;
  assign _03769_ = _03768_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9603" *) or_3538_cse;
  assign _03770_ = _03769_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9603" *) or_3542_cse;
  assign and_1104_rgt = _03770_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9603" *) and_dcpl_103;
  assign _03771_ = and_tmp_225 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9605" *) and_dcpl_401;
  assign and_1106_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9608" *) cvt_6_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _03772_ = _04289_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9614" *) and_1106_m1c;
  assign _03773_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9614" *) _05160_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_21_nl = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9616" *) and_1106_m1c;
  assign and_1115_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9621" *) cvt_7_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _03774_ = _04291_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9627" *) and_1115_m1c;
  assign _03775_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9627" *) _05374_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_19_nl = cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9629" *) and_1115_m1c;
  assign and_1119_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9634" *) cvt_8_FpMantRNE_17U_11U_else_and_3_tmp;
  assign _03776_ = _04293_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9640" *) and_1119_m1c;
  assign _03777_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9640" *) _05375_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_17_nl = cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9642" *) and_1119_m1c;
  assign _03778_ = cvt_9_FpMantRNE_17U_11U_else_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9650" *) cvt_unequal_tmp_20;
  assign and_1123_m1c = _03778_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9650" *) or_5189_cse;
  assign _03779_ = _04928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9656" *) and_1123_m1c;
  assign _03780_ = _05376_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9657" *) cvt_unequal_tmp_20;
  assign _03781_ = _03780_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9657" *) or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_15_nl = cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9659" *) and_1123_m1c;
  assign _03782_ = mux_1142_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9664" *) and_dcpl_401;
  assign and_1132_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9666" *) cvt_10_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _03783_ = _04295_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9672" *) and_1132_m1c;
  assign _03784_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9672" *) _05377_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_13_nl = cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9674" *) and_1132_m1c;
  assign _03785_ = cvt_11_FpMantRNE_17U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9682" *) cvt_unequal_tmp_20;
  assign and_1141_m1c = _03785_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9682" *) or_5189_cse;
  assign _03786_ = _04297_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9688" *) and_1141_m1c;
  assign _03787_ = _05378_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9689" *) cvt_unequal_tmp_20;
  assign _03788_ = _03787_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9689" *) or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_11_nl = cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9691" *) and_1141_m1c;
  assign _03789_ = cvt_12_FpMantRNE_17U_11U_else_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9698" *) cvt_unequal_tmp_20;
  assign and_1145_m1c = _03789_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9698" *) or_5189_cse;
  assign _03790_ = _04299_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9704" *) and_1145_m1c;
  assign _03791_ = _05379_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9705" *) cvt_unequal_tmp_20;
  assign _03792_ = _03791_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9705" *) or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_9_nl = cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9707" *) and_1145_m1c;
  assign and_283_cse = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9712" *) mux_tmp_987;
  assign _03793_ = and_dcpl_499 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9713" *) and_dcpl_626;
  assign FpIntToFloat_17U_5U_10U_is_inf_and_8_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9714" *) _09565_;
  assign _03794_ = cvt_13_FpMantRNE_17U_11U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9716" *) cvt_unequal_tmp_20;
  assign and_1155_m1c = _03794_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9716" *) or_5189_cse;
  assign _03795_ = _04301_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9721" *) and_1155_m1c;
  assign _03796_ = _05380_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9722" *) cvt_unequal_tmp_20;
  assign _03797_ = _03796_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9722" *) or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_7_nl = cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9724" *) and_1155_m1c;
  assign and_1159_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9730" *) cvt_14_FpMantRNE_17U_11U_else_and_3_tmp;
  assign _03798_ = _04303_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9735" *) and_1159_m1c;
  assign _03799_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9735" *) _05381_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_5_nl = cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9737" *) and_1159_m1c;
  assign _03800_ = and_dcpl_473 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9749" *) and_dcpl_626;
  assign FpIntToFloat_17U_5U_10U_is_inf_and_10_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9749" *) _09566_;
  assign and_1172_m1c = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9750" *) cvt_15_FpMantRNE_17U_11U_else_and_3_tmp;
  assign _03801_ = _04305_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9755" *) and_1172_m1c;
  assign _03802_ = and_dcpl_420 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9755" *) _05169_;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_3_nl = cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9757" *) and_1172_m1c;
  assign _03803_ = cvt_16_FpMantRNE_17U_11U_else_and_4_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9764" *) cvt_unequal_tmp_20;
  assign and_1176_m1c = _03803_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9764" *) or_5189_cse;
  assign _03804_ = _04307_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9769" *) and_1176_m1c;
  assign _03805_ = _05382_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9770" *) cvt_unequal_tmp_20;
  assign _03806_ = _03805_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9770" *) or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_and_1_nl = cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl[4] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9772" *) and_1176_m1c;
  assign and_271_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9778" *) mux_tmp_986;
  assign cfg_proc_precision_and_40_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9780" *) mux_1267_nl;
  assign and_295_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9781" *) or_1159_cse;
  assign cfg_proc_precision_and_43_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9783" *) mux_1268_nl;
  assign _03807_ = _05121_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9785" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c;
  assign FpFloatToInt_16U_5U_10U_and_nl = _03807_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9785" *) and_dcpl_408;
  assign _03808_ = chn_idata_data_sva_2_47_31_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9787" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c;
  assign FpFloatToInt_16U_5U_10U_and_32_nl = _03808_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9787" *) and_dcpl_408;
  assign _03809_ = cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl[11] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9789" *) _05383_;
  assign FpFloatToInt_16U_5U_10U_and_1_nl = _03809_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9789" *) and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_o_int_and_15_nl = IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9791" *) and_dcpl_408;
  assign _03810_ = or_4862_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9792" *) _04691_;
  assign and_908_nl = _03810_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9792" *) and_dcpl_420;
  assign _03811_ = or_3696_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *) or_4862_cse;
  assign _03812_ = _03811_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *) or_4714_cse;
  assign _03813_ = _03812_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *) or_400_cse_1;
  assign _03814_ = _03813_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9831" *) or_5189_cse;
  assign _03815_ = _03814_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9832" *) main_stage_v_2;
  assign _03816_ = _03815_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9832" *) _03980_;
  assign FpIntToFloat_17U_5U_10U_is_inf_and_23_cse = _01459_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9838" *) _05384_;
  assign _03817_ = and_tmp_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9839" *) and_dcpl_363;
  assign and_1213_rgt = _03817_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9839" *) or_5189_cse;
  assign _03818_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9840" *) main_stage_v_2;
  assign FpIntToFloat_17U_5U_10U_is_inf_and_26_cse = _01459_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9850" *) _05385_;
  assign FpIntToFloat_17U_5U_10U_if_and_16_cse = IntShiftRightSat_49U_6U_17U_o_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9856" *) mux_1458_nl;
  assign _03819_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9861" *) mux_1463_cse;
  assign and_1247_rgt = or_3696_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9863" *) or_5189_cse;
  assign _03820_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9869" *) mux_1460_cse;
  assign _02350_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9873" *) FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse;
  assign FpIntToFloat_17U_5U_10U_if_and_18_cse = _02350_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9873" *) mux_1465_nl;
  assign and_1250_rgt = or_tmp_2960 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9874" *) or_5189_cse;
  assign _02349_ = and_tmp_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9877" *) and_dcpl_228;
  assign and_1249_cse = _02349_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9877" *) or_5189_cse;
  assign _03821_ = cfg_out_precision_1_sva_st_149[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9879" *) mux_786_cse_1;
  assign _03822_ = cfg_out_precision_1_sva_st_154[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9884" *) mux_1489_cse;
  assign FpIntToFloat_17U_5U_10U_if_and_22_cse = _02350_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9888" *) mux_1495_nl;
  assign FpIntToFloat_17U_5U_10U_if_and_27_cse = _02350_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9895" *) mux_1521_cse;
  assign _02600_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9899" *) _05022_;
  assign IntShiftRightSat_49U_6U_17U_o_and_107_cse = _02600_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9899" *) _05391_;
  assign _03823_ = cvt_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9902" *) _05392_;
  assign IntShiftRightSat_49U_6U_17U_o_and_108_cse = _03823_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9902" *) _05393_;
  assign IntShiftRightSat_49U_6U_17U_o_and_109_cse = _02600_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9905" *) _05394_;
  assign IntShiftRightSat_49U_6U_17U_o_and_111_cse = _03823_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9907" *) _05394_;
  assign IntShiftRightSat_49U_6U_17U_o_and_112_cse = _02600_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9910" *) _05395_;
  assign IntShiftRightSat_49U_6U_17U_o_and_114_cse = _03823_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9913" *) _05396_;
  assign IntShiftRightSat_49U_6U_17U_o_and_115_cse = _03823_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9916" *) _05397_;
  assign _03824_ = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9918" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2;
  assign _03825_ = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9920" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2;
  assign _03826_ = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9922" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2;
  assign _03827_ = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9924" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2;
  assign _03828_ = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9926" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2;
  assign _03829_ = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9928" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2;
  assign _03830_ = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9930" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2;
  assign _03831_ = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9932" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2;
  assign _03832_ = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9934" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2;
  assign _03833_ = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9936" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2;
  assign _03834_ = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9938" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2;
  assign _03835_ = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9940" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2;
  assign _03836_ = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9942" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2;
  assign _03837_ = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9944" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2;
  assign _03838_ = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9946" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2;
  assign _03839_ = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9948" *) FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2;
  assign and_1321_rgt = or_dcpl_320 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9949" *) or_5189_cse;
  assign and_1325_rgt = or_dcpl_322 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9950" *) or_5189_cse;
  assign and_1329_rgt = or_dcpl_324 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9951" *) or_5189_cse;
  assign and_1333_rgt = or_dcpl_326 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9952" *) or_5189_cse;
  assign and_1337_rgt = or_dcpl_328 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9953" *) or_5189_cse;
  assign and_1341_rgt = or_dcpl_330 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9954" *) or_5189_cse;
  assign and_1345_rgt = or_dcpl_332 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9955" *) or_5189_cse;
  assign and_1349_rgt = or_dcpl_334 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9956" *) or_5189_cse;
  assign and_1353_rgt = or_dcpl_336 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9957" *) or_5189_cse;
  assign and_1357_rgt = or_dcpl_338 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9958" *) or_5189_cse;
  assign and_1361_rgt = or_dcpl_340 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9959" *) or_5189_cse;
  assign and_1365_rgt = or_dcpl_342 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9960" *) or_5189_cse;
  assign and_1369_rgt = or_dcpl_344 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9961" *) or_5189_cse;
  assign and_1373_rgt = or_dcpl_346 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9962" *) or_5189_cse;
  assign and_1377_rgt = or_dcpl_348 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9963" *) or_5189_cse;
  assign and_1381_rgt = or_dcpl_350 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9964" *) or_5189_cse;
  assign _03840_ = cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9968" *) _05398_;
  assign IntSaturation_17U_16U_and_31_rgt = _03840_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9968" *) _04174_;
  assign IntSaturation_17U_16U_o_and_31_rgt = cvt_16_IntSaturation_17U_16U_if_acc_4_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9970" *) _04174_;
  assign _03841_ = cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9974" *) _05399_;
  assign IntSaturation_17U_16U_and_29_rgt = _03841_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9974" *) _04174_;
  assign IntSaturation_17U_16U_o_and_29_rgt = cvt_15_IntSaturation_17U_16U_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9976" *) _04174_;
  assign _03842_ = cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9980" *) _05400_;
  assign IntSaturation_17U_16U_and_27_rgt = _03842_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9980" *) _04174_;
  assign IntSaturation_17U_16U_o_and_27_rgt = cvt_14_IntSaturation_17U_16U_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9982" *) _04174_;
  assign _03843_ = cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9986" *) _05401_;
  assign IntSaturation_17U_16U_and_25_rgt = _03843_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9986" *) _04174_;
  assign IntSaturation_17U_16U_o_and_25_rgt = cvt_13_IntSaturation_17U_16U_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9988" *) _04174_;
  assign _03844_ = cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9992" *) _05402_;
  assign IntSaturation_17U_16U_and_23_rgt = _03844_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9992" *) _04174_;
  assign IntSaturation_17U_16U_o_and_23_rgt = cvt_12_IntSaturation_17U_16U_if_acc_3_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9994" *) _04174_;
  assign _03845_ = cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9998" *) _05403_;
  assign IntSaturation_17U_16U_and_21_rgt = _03845_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9998" *) _04174_;
  assign and_1021_cse = cfg_proc_precision_1_sva_st_101 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10098" *) 2'b10;
  assign _03865_ = cfg_proc_precision_rsci_d == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10120" *) 2'b10;
  assign _03866_ = chn_in_rsci_d_mxwt[502:493] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11529" *) 10'b1111111111;
  assign _03867_ = chn_in_rsci_d_mxwt[470:461] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11536" *) 10'b1111111111;
  assign _03868_ = chn_in_rsci_d_mxwt[438:429] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11543" *) 10'b1111111111;
  assign _03869_ = chn_in_rsci_d_mxwt[406:397] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11550" *) 10'b1111111111;
  assign _03870_ = chn_in_rsci_d_mxwt[374:365] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11557" *) 10'b1111111111;
  assign _03871_ = chn_in_rsci_d_mxwt[342:333] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11564" *) 10'b1111111111;
  assign _03872_ = chn_in_rsci_d_mxwt[310:301] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11571" *) 10'b1111111111;
  assign _03873_ = chn_in_rsci_d_mxwt[278:269] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11578" *) 10'b1111111111;
  assign _03874_ = chn_in_rsci_d_mxwt[246:237] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11585" *) 10'b1111111111;
  assign _03875_ = chn_in_rsci_d_mxwt[214:205] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11592" *) 10'b1111111111;
  assign _03876_ = chn_in_rsci_d_mxwt[182:173] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11599" *) 10'b1111111111;
  assign _03877_ = chn_in_rsci_d_mxwt[150:141] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11604" *) 10'b1111111111;
  assign _03878_ = chn_in_rsci_d_mxwt[158:151] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11606" *) 8'b11111111;
  assign _03879_ = chn_in_rsci_d_mxwt[118:109] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11613" *) 10'b1111111111;
  assign _03880_ = chn_in_rsci_d_mxwt[86:77] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11620" *) 10'b1111111111;
  assign _03881_ = chn_in_rsci_d_mxwt[54:45] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11627" *) 10'b1111111111;
  assign _03882_ = chn_in_rsci_d_mxwt[22:13] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11634" *) 10'b1111111111;
  assign _03883_ = FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11857" *) 11'b11111111111;
  assign _03884_ = FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11859" *) 11'b11111111111;
  assign _03885_ = cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11861" *) 11'b11111111111;
  assign _03886_ = cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11863" *) 11'b11111111111;
  assign _03887_ = cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11865" *) 11'b11111111111;
  assign _03888_ = cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11867" *) 11'b11111111111;
  assign _03889_ = cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11869" *) 11'b11111111111;
  assign _03890_ = cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11871" *) 11'b11111111111;
  assign _03891_ = FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11873" *) 11'b11111111111;
  assign _03892_ = cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11875" *) 11'b11111111111;
  assign _03893_ = cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11877" *) 11'b11111111111;
  assign _03894_ = cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11879" *) 11'b11111111111;
  assign _03895_ = cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11881" *) 11'b11111111111;
  assign _03896_ = cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11883" *) 11'b11111111111;
  assign _03897_ = cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11885" *) 11'b11111111111;
  assign _03898_ = cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[16:6] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11887" *) 11'b11111111111;
  assign _03899_ = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11933" *) 33'b111111111111111111111111111111111;
  assign _03900_ = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11981" *) 33'b111111111111111111111111111111111;
  assign _03901_ = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12021" *) 33'b111111111111111111111111111111111;
  assign _03902_ = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12069" *) 33'b111111111111111111111111111111111;
  assign _03903_ = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12117" *) 33'b111111111111111111111111111111111;
  assign _03904_ = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12157" *) 33'b111111111111111111111111111111111;
  assign _03905_ = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12197" *) 33'b111111111111111111111111111111111;
  assign _03906_ = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12245" *) 33'b111111111111111111111111111111111;
  assign _03907_ = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12293" *) 33'b111111111111111111111111111111111;
  assign _03908_ = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12333" *) 33'b111111111111111111111111111111111;
  assign _03909_ = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12381" *) 33'b111111111111111111111111111111111;
  assign _03910_ = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12429" *) 33'b111111111111111111111111111111111;
  assign _03911_ = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12469" *) 33'b111111111111111111111111111111111;
  assign _03912_ = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12509" *) 33'b111111111111111111111111111111111;
  assign _03913_ = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12549" *) 33'b111111111111111111111111111111111;
  assign _03914_ = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[48:16] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12589" *) 33'b111111111111111111111111111111111;
  assign _03915_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12613" *) 19'b1111111111111111111;
  assign _03916_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12641" *) 19'b1111111111111111111;
  assign _03917_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12669" *) 19'b1111111111111111111;
  assign _03918_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12697" *) 19'b1111111111111111111;
  assign _03919_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12725" *) 19'b1111111111111111111;
  assign _03920_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12753" *) 19'b1111111111111111111;
  assign _03921_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12781" *) 19'b1111111111111111111;
  assign _03922_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12809" *) 19'b1111111111111111111;
  assign _03923_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12837" *) 19'b1111111111111111111;
  assign _03924_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12865" *) 19'b1111111111111111111;
  assign _03925_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12893" *) 19'b1111111111111111111;
  assign _03926_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12921" *) 19'b1111111111111111111;
  assign _03927_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12949" *) 19'b1111111111111111111;
  assign _03928_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12977" *) 19'b1111111111111111111;
  assign _03929_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13005" *) 19'b1111111111111111111;
  assign _03930_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[43:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13033" *) 19'b1111111111111111111;
  assign cvt_else_equal_tmp = cfg_out_precision_1_sva_6 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13184" *) 1'b1;
  assign and_2136_cse = cfg_out_precision_1_sva_6 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13213" *) 2'b11;
  assign and_dcpl_3 = cfg_proc_precision_1_sva_st_64 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14098" *) 2'b10;
  assign _03931_ = cfg_out_precision_1_sva_st_113 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14473" *) 2'b10;
  assign _03932_ = reg_cfg_proc_precision_1_sva_st_40_cse == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14682" *) 2'b10;
  assign and_dcpl_228 = cfg_out_precision_1_sva_st_154 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14695" *) 2'b10;
  assign _03933_ = cfg_out_precision_1_sva_st_113 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14748" *) 1'b1;
  assign and_dcpl_479 = cfg_proc_precision_1_sva_st_89 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14750" *) 2'b10;
  assign _03934_ = cfg_proc_precision_1_sva_st_90 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14767" *) 2'b10;
  assign and_dcpl_535 = cfg_proc_precision_1_sva_st_102 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14768" *) 2'b10;
  assign and_1059_cse = cfg_proc_precision_1_sva_st_108 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14771" *) 2'b10;
  assign and_dcpl_942 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14823" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16;
  assign and_dcpl_946 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14825" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17;
  assign and_dcpl_950 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14826" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18;
  assign and_dcpl_954 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14829" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19;
  assign and_dcpl_958 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14830" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20;
  assign and_dcpl_962 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14833" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21;
  assign and_dcpl_966 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14836" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22;
  assign and_dcpl_970 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14837" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23;
  assign and_dcpl_974 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14838" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24;
  assign and_dcpl_978 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14840" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25;
  assign and_dcpl_982 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14842" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26;
  assign and_dcpl_987 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14843" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27;
  assign and_dcpl_991 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14845" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28;
  assign and_dcpl_995 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14846" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29;
  assign and_dcpl_999 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14847" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30;
  assign and_dcpl_1003 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14848" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31;
  assign _03935_ = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16303" *) 5'b11111;
  assign _03936_ = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16311" *) 5'b11111;
  assign _03937_ = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16319" *) 5'b11111;
  assign _03938_ = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16327" *) 5'b11111;
  assign _03939_ = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16335" *) 5'b11111;
  assign _03940_ = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16343" *) 5'b11111;
  assign _03941_ = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16351" *) 5'b11111;
  assign _03942_ = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16359" *) 5'b11111;
  assign _03943_ = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16367" *) 5'b11111;
  assign _03944_ = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16375" *) 5'b11111;
  assign _03945_ = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16383" *) 5'b11111;
  assign _03946_ = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16392" *) 5'b11111;
  assign _03947_ = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16400" *) 5'b11111;
  assign _03948_ = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16408" *) 5'b11111;
  assign _03949_ = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16416" *) 5'b11111;
  assign _03950_ = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16424" *) 5'b11111;
  assign _03951_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *) 4'b1111;
  assign _03952_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *) 4'b1111;
  assign _03953_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *) 4'b1111;
  assign _03954_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *) 4'b1111;
  assign _03955_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *) 4'b1111;
  assign _03956_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *) 4'b1111;
  assign _03957_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *) 4'b1111;
  assign _03958_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *) 4'b1111;
  assign _03959_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *) 4'b1111;
  assign _03960_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *) 4'b1111;
  assign _03961_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *) 4'b1111;
  assign _03962_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *) 4'b1111;
  assign _03963_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *) 4'b1111;
  assign and_2360_cse = cfg_proc_precision_1_sva_st_65 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18485" *) 2'b10;
  assign _03964_ = IntShiftRightSat_49U_6U_17U_i_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18754" *) { cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl };
  assign _03965_ = IntShiftRightSat_49U_6U_17U_i_15_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18759" *) { cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl };
  assign _03966_ = IntShiftRightSat_49U_6U_17U_i_14_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18762" *) { cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl };
  assign _03967_ = IntShiftRightSat_49U_6U_17U_i_13_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18765" *) { cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl };
  assign _03968_ = IntShiftRightSat_49U_6U_17U_i_12_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18768" *) { cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl };
  assign _03969_ = IntShiftRightSat_49U_6U_17U_i_11_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18771" *) { cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl };
  assign _03970_ = IntShiftRightSat_49U_6U_17U_i_10_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18774" *) { cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl };
  assign _03971_ = IntShiftRightSat_49U_6U_17U_i_9_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18777" *) { cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl };
  assign _03972_ = IntShiftRightSat_49U_6U_17U_i_8_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18780" *) { cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl };
  assign _03973_ = IntShiftRightSat_49U_6U_17U_i_7_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18783" *) { cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl };
  assign _03974_ = IntShiftRightSat_49U_6U_17U_i_6_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18786" *) { cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl };
  assign _03975_ = IntShiftRightSat_49U_6U_17U_i_5_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18789" *) { cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl };
  assign _03976_ = IntShiftRightSat_49U_6U_17U_i_4_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18792" *) { cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl };
  assign _03977_ = IntShiftRightSat_49U_6U_17U_i_3_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18795" *) { cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl };
  assign _03978_ = IntShiftRightSat_49U_6U_17U_i_2_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18798" *) { cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl };
  assign _03979_ = IntShiftRightSat_49U_6U_17U_i_1_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18801" *) { cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl };
  assign _03980_ = cfg_out_precision_1_sva_st_149 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19040" *) 2'b10;
  assign _03981_ = FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23360" *) 12'b111111111111;
  assign _03982_ = FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23387" *) 12'b111111111111;
  assign _03983_ = cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23406" *) 12'b111111111111;
  assign _03984_ = cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23420" *) 12'b111111111111;
  assign _03985_ = cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23429" *) 12'b111111111111;
  assign _03986_ = cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23447" *) 12'b111111111111;
  assign _03987_ = cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23459" *) 12'b111111111111;
  assign _03988_ = cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23475" *) 12'b111111111111;
  assign _03989_ = FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23493" *) 12'b111111111111;
  assign _03990_ = cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23504" *) 12'b111111111111;
  assign _03991_ = cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23516" *) 12'b111111111111;
  assign _03992_ = cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23537" *) 12'b111111111111;
  assign _03993_ = cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23546" *) 12'b111111111111;
  assign _03994_ = cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23567" *) 12'b111111111111;
  assign _03995_ = cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23576" *) 12'b111111111111;
  assign _03996_ = cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[16:5] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23585" *) 12'b111111111111;
  assign _03997_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24099" *) 4'b1111;
  assign _03998_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24110" *) 4'b1111;
  assign _03999_ = FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24119" *) 4'b1111;
  assign _04000_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9129" *) cfg_out_precision_1_sva_st_113;
  assign _04001_ = $signed(cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16437" *) $signed(cfg_scale_rsci_d);
  assign _04002_ = $signed(cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16439" *) $signed(cfg_scale_rsci_d);
  assign _04003_ = $signed(cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16441" *) $signed(cfg_scale_rsci_d);
  assign _04004_ = $signed(cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16496" *) $signed(cfg_scale_rsci_d);
  assign _04005_ = $signed(cvt_1_IntSubExt_32U_32U_33U_o_acc_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16515" *) $signed(cfg_scale_rsci_d);
  assign cvt_4_IntMulExt_33U_16U_49U_o_mul_2_nl = $signed(cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22421" *) $signed(cfg_scale_rsci_d);
  assign cvt_6_IntMulExt_33U_16U_49U_o_mul_2_nl = $signed(cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22426" *) $signed(cfg_scale_rsci_d);
  assign cvt_8_IntMulExt_33U_16U_49U_o_mul_3_nl = $signed(cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22431" *) $signed(cfg_scale_rsci_d);
  assign cvt_7_IntMulExt_33U_16U_49U_o_mul_2_nl = $signed(cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22436" *) $signed(cfg_scale_rsci_d);
  assign cvt_10_IntMulExt_33U_16U_49U_o_mul_2_nl = $signed(cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22441" *) $signed(cfg_scale_rsci_d);
  assign cvt_12_IntMulExt_33U_16U_49U_o_mul_3_nl = $signed(cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22446" *) $signed(cfg_scale_rsci_d);
  assign cvt_11_IntMulExt_33U_16U_49U_o_mul_2_nl = $signed(cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22451" *) $signed(cfg_scale_rsci_d);
  assign cvt_14_IntMulExt_33U_16U_49U_o_mul_3_nl = $signed(cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22456" *) $signed(cfg_scale_rsci_d);
  assign cvt_16_IntMulExt_33U_16U_49U_o_mul_4_nl = $signed(cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22461" *) $signed(cfg_scale_rsci_d);
  assign cvt_15_IntMulExt_33U_16U_49U_o_mul_3_nl = $signed(cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22466" *) $signed(cfg_scale_rsci_d);
  assign cvt_13_IntMulExt_33U_16U_49U_o_mul_2_nl = $signed(cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22471" *) $signed(cfg_scale_rsci_d);
  assign _04006_ = cfg_out_precision_1_sva_st_154 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10064" *) 1'b1;
  assign or_309_cse = cfg_out_precision_1_sva_st_149 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10065" *) 1'b1;
  assign or_183_cse_1 = reg_cfg_proc_precision_1_sva_st_40_cse != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10097" *) 2'b10;
  assign or_2251_nl = cfg_out_precision_1_sva_st_154 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10106" *) 2'b10;
  assign _04007_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10819" *) IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0;
  assign _04008_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10831" *) IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0;
  assign cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp = IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10834" *) { IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0 };
  assign _04009_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10846" *) IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0;
  assign cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp = IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10859" *) { IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0 };
  assign cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp = IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10862" *) { IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0 };
  assign _04010_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10874" *) IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0;
  assign cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp = IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10887" *) { IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0 };
  assign cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp = IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10910" *) { IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0 };
  assign cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp = IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10913" *) { IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0 };
  assign cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp = IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10916" *) { IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0 };
  assign _04011_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10928" *) IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0;
  assign cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp = IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11001" *) { IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0 };
  assign cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp = IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11004" *) { IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0 };
  assign _04012_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11410" *) IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0;
  assign _04013_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11412" *) IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0;
  assign _04014_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11415" *) IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0;
  assign _04015_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11418" *) IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0;
  assign _04016_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11421" *) IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0;
  assign _04017_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11423" *) IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0;
  assign _04018_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11425" *) IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0;
  assign _04019_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11427" *) IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0;
  assign _04020_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11429" *) IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0;
  assign _04021_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11432" *) IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0;
  assign _04022_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11435" *) IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0;
  assign _04023_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11523" *) chn_in_rsci_d_mxwt[502:480];
  assign _04024_ = chn_in_rsci_d_mxwt[510:503] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11524" *) 8'b11111111;
  assign _04025_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11530" *) chn_in_rsci_d_mxwt[470:448];
  assign _04026_ = chn_in_rsci_d_mxwt[478:471] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11531" *) 8'b11111111;
  assign _04027_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11537" *) chn_in_rsci_d_mxwt[438:416];
  assign _04028_ = chn_in_rsci_d_mxwt[446:439] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11538" *) 8'b11111111;
  assign _04029_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11544" *) chn_in_rsci_d_mxwt[406:384];
  assign _04030_ = chn_in_rsci_d_mxwt[414:407] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11545" *) 8'b11111111;
  assign _04031_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11551" *) chn_in_rsci_d_mxwt[374:352];
  assign _04032_ = chn_in_rsci_d_mxwt[382:375] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11552" *) 8'b11111111;
  assign _04033_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11558" *) chn_in_rsci_d_mxwt[342:320];
  assign _04034_ = chn_in_rsci_d_mxwt[350:343] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11559" *) 8'b11111111;
  assign _04035_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11565" *) chn_in_rsci_d_mxwt[310:288];
  assign _04036_ = chn_in_rsci_d_mxwt[318:311] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11566" *) 8'b11111111;
  assign _04037_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11572" *) chn_in_rsci_d_mxwt[278:256];
  assign _04038_ = chn_in_rsci_d_mxwt[286:279] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11573" *) 8'b11111111;
  assign _04039_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11579" *) chn_in_rsci_d_mxwt[246:224];
  assign _04040_ = chn_in_rsci_d_mxwt[254:247] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11580" *) 8'b11111111;
  assign _04041_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11586" *) chn_in_rsci_d_mxwt[214:192];
  assign _04042_ = chn_in_rsci_d_mxwt[222:215] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11587" *) 8'b11111111;
  assign _04043_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11593" *) chn_in_rsci_d_mxwt[182:160];
  assign _04044_ = chn_in_rsci_d_mxwt[190:183] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11594" *) 8'b11111111;
  assign _04045_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11605" *) chn_in_rsci_d_mxwt[150:128];
  assign _04046_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11607" *) chn_in_rsci_d_mxwt[118:96];
  assign _04047_ = chn_in_rsci_d_mxwt[126:119] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11608" *) 8'b11111111;
  assign _04048_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11614" *) chn_in_rsci_d_mxwt[86:64];
  assign _04049_ = chn_in_rsci_d_mxwt[94:87] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11615" *) 8'b11111111;
  assign _04050_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11621" *) chn_in_rsci_d_mxwt[54:32];
  assign _04051_ = chn_in_rsci_d_mxwt[62:55] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11622" *) 8'b11111111;
  assign _04052_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11628" *) chn_in_rsci_d_mxwt[22:0];
  assign _04053_ = chn_in_rsci_d_mxwt[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11629" *) 8'b11111111;
  assign cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp = IntShiftRightSat_49U_6U_17U_i_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11741" *) { IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0 };
  assign cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp = IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11744" *) { IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0 };
  assign cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp = IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11747" *) { IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0 };
  assign cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp = IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11750" *) { IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0 };
  assign cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp = IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11753" *) { IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0 };
  assign _04054_ = IntShiftRightSat_49U_6U_17U_i_2_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11759" *) { cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl };
  assign _04055_ = IntShiftRightSat_49U_6U_17U_i_4_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11765" *) { cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl };
  assign _04056_ = IntShiftRightSat_49U_6U_17U_i_3_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11771" *) { cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl };
  assign _04057_ = IntShiftRightSat_49U_6U_17U_i_6_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11777" *) { cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl };
  assign _04058_ = IntShiftRightSat_49U_6U_17U_i_8_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11783" *) { cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl };
  assign _04059_ = IntShiftRightSat_49U_6U_17U_i_7_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11789" *) { cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl };
  assign _04060_ = IntShiftRightSat_49U_6U_17U_i_5_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11795" *) { cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl };
  assign _04061_ = IntShiftRightSat_49U_6U_17U_i_10_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11801" *) { cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl };
  assign cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp = IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11804" *) { IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0 };
  assign _04062_ = IntShiftRightSat_49U_6U_17U_i_12_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11810" *) { cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl };
  assign _04063_ = IntShiftRightSat_49U_6U_17U_i_11_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11816" *) { cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl };
  assign cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp = IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11819" *) { IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0, IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0 };
  assign _04064_ = IntShiftRightSat_49U_6U_17U_i_14_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11825" *) { _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17], _03864_[17:9], cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl };
  assign _04065_ = IntShiftRightSat_49U_6U_17U_i_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11831" *) { cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17], cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl };
  assign _04066_ = IntShiftRightSat_49U_6U_17U_i_15_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11837" *) { cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17], cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl };
  assign _04067_ = IntShiftRightSat_49U_6U_17U_i_13_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11843" *) { cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17], cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl };
  assign _04068_ = IntShiftRightSat_49U_6U_17U_i_9_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11849" *) { cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17], cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl };
  assign _04069_ = IntShiftRightSat_49U_6U_17U_i_1_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11855" *) { cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17], cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl };
  assign _04070_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11935" *) cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16];
  assign _04071_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11983" *) cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16];
  assign _04072_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12023" *) cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16];
  assign _04073_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12071" *) cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16];
  assign _04074_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12119" *) cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16];
  assign _04075_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12159" *) cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16];
  assign _04076_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12199" *) cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16];
  assign _04077_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12247" *) cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16];
  assign _04078_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12295" *) cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16];
  assign _04079_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12335" *) cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16];
  assign _04080_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12383" *) cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16];
  assign _04081_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12431" *) cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[48:16];
  assign _04082_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12471" *) cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16];
  assign _04083_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12511" *) cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16];
  assign _04084_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12551" *) cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16];
  assign _04085_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12591" *) cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[48:16];
  assign _04086_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12615" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[43:25];
  assign _04087_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12643" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[43:25];
  assign _04088_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12671" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[43:25];
  assign _04089_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12699" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[43:25];
  assign _04090_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12727" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[43:25];
  assign _04091_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12755" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[43:25];
  assign _04092_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12783" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[43:25];
  assign _04093_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12811" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[43:25];
  assign _04094_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12839" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[43:25];
  assign _04095_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12867" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[43:25];
  assign _04096_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12895" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[43:25];
  assign _04097_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12923" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[43:25];
  assign _04098_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12951" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[43:25];
  assign _04099_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12979" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[43:25];
  assign _04100_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13007" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[43:25];
  assign _04101_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13035" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[43:25];
  assign or_1431_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13215" *) cfg_out_precision_1_sva_6;
  assign _04102_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13527" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva;
  assign _04103_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13528" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva;
  assign _04104_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13529" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva;
  assign _04105_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13543" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva;
  assign _04106_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13544" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva;
  assign _04107_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13545" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva;
  assign _04108_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13559" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva;
  assign _04109_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13560" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva;
  assign _04110_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13561" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva;
  assign _04111_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13575" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_4_sva;
  assign _04112_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13576" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_4_sva;
  assign _04113_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13577" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_4_sva;
  assign _04114_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13591" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_5_sva;
  assign _04115_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13592" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_5_sva;
  assign _04116_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13593" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_5_sva;
  assign _04117_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13607" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_6_sva;
  assign _04118_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13608" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_6_sva;
  assign _04119_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13609" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_6_sva;
  assign _04120_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13623" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_7_sva;
  assign _04121_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13624" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_7_sva;
  assign _04122_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13625" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_7_sva;
  assign _04123_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13639" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_8_sva;
  assign _04124_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13640" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_8_sva;
  assign _04125_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13641" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_8_sva;
  assign _04126_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13655" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_9_sva;
  assign _04127_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13656" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_9_sva;
  assign _04128_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13657" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_9_sva;
  assign _04129_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13671" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_10_sva;
  assign _04130_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13672" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_10_sva;
  assign _04131_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13673" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_10_sva;
  assign _04132_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13687" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_11_sva;
  assign _04133_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13688" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_11_sva;
  assign _04134_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13689" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_11_sva;
  assign _04135_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13703" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_12_sva;
  assign _04136_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13704" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_12_sva;
  assign _04137_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13705" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_12_sva;
  assign _04138_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13719" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_13_sva;
  assign _04139_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13720" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_13_sva;
  assign _04140_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13721" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_13_sva;
  assign _04141_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13735" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_14_sva;
  assign _04142_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13736" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_14_sva;
  assign _04143_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13737" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_14_sva;
  assign _04144_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13751" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_15_sva;
  assign _04145_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13752" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_15_sva;
  assign _04146_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13753" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_15_sva;
  assign _04147_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13767" *) FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva;
  assign _04148_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13768" *) FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva;
  assign _04149_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13769" *) FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva;
  assign or_4550_cse = cfg_proc_precision_1_sva_st_64 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14108" *) 2'b10;
  assign or_2242_nl = cfg_out_precision_rsci_d != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14124" *) 2'b10;
  assign or_4862_cse = cfg_proc_precision_1_sva_st_65 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14142" *) 2'b10;
  assign or_578_cse = cfg_out_precision_1_sva_st_149 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14190" *) 2'b10;
  assign or_425_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14214" *) cfg_out_precision_1_sva_st_113;
  assign or_461_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14317" *) cfg_out_precision_1_sva_st_149;
  assign _04150_ = cfg_out_precision_1_sva_6 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14501" *) 2'b10;
  assign or_1198_cse = cfg_out_precision_1_sva_st_113 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14509" *) 2'b10;
  assign _04151_ = cfg_out_precision_1_sva_st_156 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14525" *) 2'b10;
  assign or_1157_cse = cfg_out_precision_1_sva_6 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14563" *) 1'b1;
  assign or_300_cse = cfg_out_precision_1_sva_st_113 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14739" *) 1'b1;
  assign _04152_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16667" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_5_mx0;
  assign _04153_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16669" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_5_mx0;
  assign _04154_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16671" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_5_mx0;
  assign _04155_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16673" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_5_mx0;
  assign _04156_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16675" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_5_mx0;
  assign _04157_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16677" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_5_mx0;
  assign _04158_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16679" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_5_mx0;
  assign _04159_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16681" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_5_mx0;
  assign _04160_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16683" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_5_mx0;
  assign _04161_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16685" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_5_mx0;
  assign _04162_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16687" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_5_mx0;
  assign _04163_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16689" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_5_mx0;
  assign _04164_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16691" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_5_mx0;
  assign or_4524_cse = cfg_proc_precision_rsci_d != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *) 2'b10;
  assign or_961_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22543" *) cfg_out_precision_1_sva_st_154;
  assign _04165_ = cfg_out_precision_1_sva_st_136 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22924" *) 2'b10;
  assign or_1720_cse_1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21;
  assign or_5069_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23116" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30;
  assign _04166_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23307" *) cfg_out_precision_1_sva_st_136;
  assign _04167_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23326" *) cfg_out_precision_1_sva_st_144;
  assign or_1202_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16;
  assign _04168_ = cfg_out_precision_rsci_d != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23629" *) 1'b1;
  assign _04169_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24092" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_5_mx0;
  assign _04170_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24105" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_5_mx0;
  assign _04171_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24114" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_5_mx0;
  assign _04172_ = cfg_out_precision_1_sva_6 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8776" *) 2'b11;
  assign or_5254_cse = cfg_proc_precision_1_sva_st_108 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8803" *) 2'b10;
  assign or_400_cse_1 = cfg_proc_precision_1_sva_st_101 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8863" *) 2'b10;
  assign or_1159_cse = cfg_proc_precision_1_sva_st_66 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9083" *) 2'b10;
  assign or_3538_cse = cfg_proc_precision_1_sva_st_90 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9111" *) 2'b10;
  assign or_4714_cse = cfg_proc_precision_1_sva_st_89 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9144" *) 2'b10;
  assign or_3542_cse = cfg_proc_precision_1_sva_st_102 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9325" *) 2'b10;
  assign or_1596_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9528" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17;
  assign _04173_ = cfg_out_precision_1_sva_st_144 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *) 2'b10;
  assign or_1625_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9549" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18;
  assign or_1659_cse_1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9576" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19;
  assign or_1693_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9590" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20;
  assign or_1752_cse_1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9622" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22;
  assign or_1789_cse_1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9635" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23;
  assign or_1829_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9651" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24;
  assign or_1851_cse_1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9667" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25;
  assign or_1892_cse_1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9683" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26;
  assign or_1925_cse_1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9699" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27;
  assign or_5038_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9729" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28;
  assign or_5053_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9742" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29;
  assign or_5086_cse = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9777" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31;
  assign _04174_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10000" *) and_dcpl_93;
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10002" *) _05405_;
  assign _04175_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10004" *) cvt_10_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10008" *) _05407_;
  assign _04176_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10010" *) cvt_9_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10014" *) _05409_;
  assign _04177_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10016" *) cvt_8_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10020" *) _05411_;
  assign _04178_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10022" *) cvt_7_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10026" *) _05413_;
  assign _04179_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10028" *) cvt_6_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10032" *) _05415_;
  assign _04180_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10034" *) cvt_5_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10038" *) _05417_;
  assign _04181_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10040" *) cvt_4_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10044" *) _05419_;
  assign _04182_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10046" *) cvt_3_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10050" *) _05421_;
  assign _04183_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10052" *) cvt_2_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10056" *) _05423_;
  assign _04184_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10058" *) cvt_1_IntSaturation_17U_16U_if_acc_nl[2];
  assign _04185_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *) main_stage_v_1;
  assign _04186_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *) cvt_unequal_tmp_19;
  assign nor_1195_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *) _05425_;
  assign nor_1185_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10064" *) _05426_;
  assign _00058_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10065" *) main_stage_v_2;
  assign nor_1186_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10065" *) _05427_;
  assign _00064_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10072" *) and_1386_cse;
  assign _04187_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10076" *) and_tmp_16;
  assign _04188_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10081" *) and_tmp_19;
  assign _00065_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10095" *) and_2186_cse;
  assign _00018_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10099" *) mux_tmp_1276;
  assign _00019_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10101" *) mux_1284_nl;
  assign _04189_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10104" *) mux_1286_nl;
  assign FpIntToFloat_17U_5U_10U_if_nor_10_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10106" *) _05429_;
  assign FpIntToFloat_17U_5U_10U_if_nor_6_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10115" *) _05430_;
  assign cvt_cvt_nand_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10120" *) _03865_;
  assign _03847_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10137" *) chn_in_rsci_d_mxwt[26:24];
  assign _04190_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10140" *) chn_in_rsci_d_mxwt[30:23];
  assign _03848_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10149" *) chn_in_rsci_d_mxwt[58:56];
  assign _04191_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10153" *) chn_in_rsci_d_mxwt[62:55];
  assign _03849_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10161" *) chn_in_rsci_d_mxwt[90:88];
  assign _04192_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10165" *) chn_in_rsci_d_mxwt[94:87];
  assign _03850_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10173" *) chn_in_rsci_d_mxwt[122:120];
  assign _04193_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10177" *) chn_in_rsci_d_mxwt[126:119];
  assign _03851_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10185" *) chn_in_rsci_d_mxwt[154:152];
  assign _04194_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10189" *) chn_in_rsci_d_mxwt[158:151];
  assign _03852_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10197" *) chn_in_rsci_d_mxwt[186:184];
  assign _04195_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10201" *) chn_in_rsci_d_mxwt[190:183];
  assign _03853_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10209" *) chn_in_rsci_d_mxwt[218:216];
  assign _04196_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10213" *) chn_in_rsci_d_mxwt[222:215];
  assign _03854_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10221" *) chn_in_rsci_d_mxwt[250:248];
  assign _04197_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10225" *) chn_in_rsci_d_mxwt[254:247];
  assign _03855_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10233" *) chn_in_rsci_d_mxwt[282:280];
  assign _04198_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10237" *) chn_in_rsci_d_mxwt[286:279];
  assign _03856_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10245" *) chn_in_rsci_d_mxwt[314:312];
  assign _04199_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10249" *) chn_in_rsci_d_mxwt[318:311];
  assign _03857_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10257" *) chn_in_rsci_d_mxwt[346:344];
  assign _04200_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10261" *) chn_in_rsci_d_mxwt[350:343];
  assign _03858_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10269" *) chn_in_rsci_d_mxwt[378:376];
  assign _04201_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10273" *) chn_in_rsci_d_mxwt[382:375];
  assign _03859_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10281" *) chn_in_rsci_d_mxwt[410:408];
  assign _04202_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10285" *) chn_in_rsci_d_mxwt[414:407];
  assign _03860_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10293" *) chn_in_rsci_d_mxwt[442:440];
  assign _04203_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10297" *) chn_in_rsci_d_mxwt[446:439];
  assign _03861_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10305" *) chn_in_rsci_d_mxwt[474:472];
  assign _04204_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10309" *) chn_in_rsci_d_mxwt[478:471];
  assign _03862_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10317" *) chn_in_rsci_d_mxwt[506:504];
  assign _04205_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10321" *) chn_in_rsci_d_mxwt[510:503];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10398" *) _00075_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10401" *) _00076_;
  assign _04206_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10402" *) cvt_1_FpMantRNE_24U_11U_else_and_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10424" *) _00077_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10427" *) _00078_;
  assign _04207_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10428" *) cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10450" *) _00079_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10453" *) _00080_;
  assign _04208_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10454" *) cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10476" *) _00081_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10479" *) _00082_;
  assign _04209_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10480" *) cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10502" *) _00083_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10505" *) _00084_;
  assign _04210_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10506" *) cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10528" *) _00085_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10531" *) _00086_;
  assign _04211_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10532" *) cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10554" *) _00087_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10557" *) _00088_;
  assign _04212_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10558" *) cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10580" *) _00089_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10583" *) _00090_;
  assign _04213_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10584" *) cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10606" *) _00091_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10609" *) _00092_;
  assign _04214_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10610" *) cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10632" *) _00093_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10635" *) _00094_;
  assign _04215_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10636" *) cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10658" *) _00095_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10661" *) _00096_;
  assign _04216_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10662" *) cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10684" *) _00097_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10687" *) _00098_;
  assign _04217_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10688" *) cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10710" *) _00099_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10713" *) _00100_;
  assign _04218_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10714" *) cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10736" *) _00101_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10739" *) _00102_;
  assign _04219_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10740" *) cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10762" *) _00103_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10765" *) _00104_;
  assign _04220_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10766" *) cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10788" *) _00105_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10791" *) _00106_;
  assign _04221_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10792" *) cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2;
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_4_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10809" *) _05431_;
  assign IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10811" *) _00187_[2];
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10813" *) _00107_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10815" *) _00108_;
  assign _04222_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10817" *) _05432_;
  assign IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10817" *) _00203_[0];
  assign cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10819" *) _05434_;
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10821" *) _05435_;
  assign IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10823" *) _00188_[2];
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10825" *) _00109_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10827" *) _00110_;
  assign _04223_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10829" *) _05436_;
  assign IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10829" *) _00204_[0];
  assign cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10831" *) _05438_;
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10836" *) _05439_;
  assign IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10838" *) _00189_[2];
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10840" *) _00111_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10842" *) _00112_;
  assign _04224_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10844" *) _05440_;
  assign IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10844" *) _00205_[0];
  assign cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10846" *) _05442_;
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10848" *) or_dcpl_108;
  assign IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10850" *) or_dcpl_109;
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10852" *) _00113_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10854" *) _00114_;
  assign _04225_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10856" *) _05443_;
  assign IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10856" *) _00206_[0];
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10864" *) or_dcpl_110;
  assign IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10866" *) or_dcpl_111;
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10868" *) _00115_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10870" *) _00116_;
  assign _04226_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10872" *) _05444_;
  assign IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10872" *) _00207_[0];
  assign cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10874" *) _05446_;
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10876" *) or_dcpl_113;
  assign IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10878" *) or_dcpl_114;
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10880" *) _00117_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10882" *) _00118_;
  assign _04227_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10884" *) _05447_;
  assign IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10884" *) _00208_[0];
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10889" *) or_dcpl_115;
  assign IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10891" *) or_dcpl_116;
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10893" *) _00119_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10895" *) _00120_;
  assign _04228_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10897" *) _05448_;
  assign IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10897" *) _00209_[0];
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10899" *) or_dcpl_119;
  assign IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10901" *) or_dcpl_120;
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10903" *) _00121_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10905" *) _00122_;
  assign _04229_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10907" *) _05449_;
  assign IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10907" *) _00210_[0];
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10918" *) _05450_;
  assign IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10920" *) _00195_[2];
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10922" *) _00123_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10924" *) _00124_;
  assign _04230_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10926" *) _05451_;
  assign IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10926" *) _00211_[0];
  assign cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10928" *) _05453_;
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10930" *) or_dcpl_124;
  assign IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10932" *) or_dcpl_125;
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10934" *) _00125_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10936" *) _00126_;
  assign _04231_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10938" *) _05454_;
  assign IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10938" *) _00212_[0];
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10940" *) or_dcpl_126;
  assign IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10942" *) or_dcpl_127;
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10944" *) _00127_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10946" *) _00128_;
  assign _04232_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10948" *) _05455_;
  assign IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10948" *) _00213_[0];
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10950" *) or_dcpl_130;
  assign IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10952" *) or_dcpl_131;
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10954" *) _00129_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10956" *) _00130_;
  assign _04233_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10958" *) _05456_;
  assign IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10958" *) _00214_[0];
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10960" *) or_dcpl_132;
  assign IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10962" *) or_dcpl_133;
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10964" *) _00131_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10966" *) _00132_;
  assign _04234_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10968" *) _05457_;
  assign IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10968" *) _00215_[0];
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10970" *) or_dcpl_136;
  assign IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10972" *) or_dcpl_137;
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10974" *) _00133_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10976" *) _00134_;
  assign _04235_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10978" *) _05458_;
  assign IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10978" *) _00216_[0];
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10980" *) or_dcpl_139;
  assign IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10982" *) or_dcpl_140;
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10984" *) _00135_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10986" *) _00136_;
  assign _04236_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10988" *) _05459_;
  assign IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10988" *) _00217_[0];
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_24_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10990" *) or_dcpl_143;
  assign IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10992" *) or_dcpl_144;
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_22_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10994" *) _00137_;
  assign IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10996" *) _00138_;
  assign _04237_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10998" *) _05460_;
  assign IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10998" *) _00218_[0];
  assign _04238_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11006" *) _05461_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11006" *) _04519_;
  assign _04239_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11008" *) _05462_;
  assign _04240_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11011" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva[23:14];
  assign IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11014" *) _05383_;
  assign _04241_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11016" *) _05463_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11016" *) _04521_;
  assign _04242_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11018" *) _05464_;
  assign _04243_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11021" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva[23:14];
  assign IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11024" *) _05333_;
  assign _04244_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11026" *) _05465_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11026" *) _04523_;
  assign _00171_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11027" *) IntShiftRightSat_49U_6U_17U_o_16_3_sva_3;
  assign _00171_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11028" *) IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2[14:6];
  assign _04245_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11032" *) _05466_;
  assign _04246_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11035" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva[23:14];
  assign _04247_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11039" *) _05467_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11039" *) _04525_;
  assign _04248_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11041" *) _05468_;
  assign _04249_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11044" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva[23:14];
  assign _04250_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11048" *) _05469_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11048" *) _04527_;
  assign _00172_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11049" *) IntShiftRightSat_49U_6U_17U_o_16_5_sva_3;
  assign _00172_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11050" *) IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2[14:6];
  assign _04251_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11054" *) _05470_;
  assign _04252_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11057" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva[23:14];
  assign _04253_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11061" *) _05471_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11061" *) _04549_;
  assign _04254_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11063" *) _05472_;
  assign _04255_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11066" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_sva[23:14];
  assign _04256_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11070" *) _05473_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11070" *) _04529_;
  assign _04257_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11072" *) _05474_;
  assign _04258_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11075" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva[23:14];
  assign _04259_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11079" *) _05475_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11079" *) _04547_;
  assign _00173_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11080" *) IntShiftRightSat_49U_6U_17U_o_16_1_sva_3;
  assign _00173_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11081" *) IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2[14:6];
  assign _04260_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11085" *) _05476_;
  assign _04261_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11088" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva[23:14];
  assign IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11091" *) _05341_;
  assign _04262_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11093" *) _05477_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11093" *) _04531_;
  assign _04263_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11095" *) _05478_;
  assign _04264_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11098" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva[23:14];
  assign _04265_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11102" *) _05479_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11102" *) _04545_;
  assign _04266_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11104" *) _05480_;
  assign _04267_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11107" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva[23:14];
  assign _04268_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11111" *) _05481_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11111" *) _04533_;
  assign _04269_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11113" *) _05482_;
  assign _04270_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11116" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva[23:14];
  assign _04271_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11120" *) _05483_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11120" *) _04543_;
  assign _04272_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11122" *) _05484_;
  assign _04273_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11125" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva[23:14];
  assign _04274_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11129" *) _05485_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11129" *) _04535_;
  assign _00174_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11130" *) IntShiftRightSat_49U_6U_17U_o_16_9_sva_3;
  assign _00174_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11131" *) IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2[14:6];
  assign _04275_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11135" *) _05486_;
  assign _04276_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11138" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva[23:14];
  assign _04277_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11142" *) _05487_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11142" *) _04541_;
  assign _04278_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11144" *) _05488_;
  assign _04279_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11147" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva[23:14];
  assign _04280_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11151" *) _05489_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11151" *) _04537_;
  assign _04281_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11153" *) _05490_;
  assign _04282_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11156" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva[23:14];
  assign _04283_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11160" *) _05491_;
  assign FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11160" *) _04539_;
  assign _04284_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11162" *) _05492_;
  assign _04285_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11165" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva[23:14];
  assign _04286_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11235" *) cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign _04287_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11260" *) cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign _04288_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11261" *) _01463_;
  assign FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11262" *) _05493_;
  assign _04289_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11280" *) cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign _04290_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11281" *) _01465_;
  assign FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11282" *) _05494_;
  assign _04291_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11294" *) cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign _04292_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11295" *) _01467_;
  assign FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11296" *) _05495_;
  assign _04293_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11308" *) cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign _04294_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11309" *) _01469_;
  assign FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11310" *) _05496_;
  assign _04295_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11322" *) cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign _04296_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11323" *) _01471_;
  assign FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11324" *) _05497_;
  assign _04297_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11336" *) cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign _04298_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11337" *) _01473_;
  assign FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11338" *) _05498_;
  assign _04299_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11350" *) cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign _04300_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11351" *) _01475_;
  assign FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11352" *) _05499_;
  assign _04301_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11364" *) cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign _04302_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11365" *) _01477_;
  assign FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11366" *) _05500_;
  assign _04303_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11378" *) cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign _04304_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11379" *) _01479_;
  assign FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11380" *) _05501_;
  assign _04305_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11392" *) cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign _04306_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11393" *) _01481_;
  assign FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11394" *) _05502_;
  assign _04307_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11406" *) cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl[4];
  assign _04308_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11407" *) _01483_;
  assign FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11408" *) _05503_;
  assign cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11410" *) _05505_;
  assign cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11413" *) _05507_;
  assign cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11416" *) _05509_;
  assign cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11419" *) _05511_;
  assign cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11421" *) _05513_;
  assign cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11423" *) _05515_;
  assign cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11425" *) _05517_;
  assign cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11427" *) _05519_;
  assign cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11430" *) _05521_;
  assign cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11433" *) _05523_;
  assign cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11436" *) _05525_;
  assign _04309_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11523" *) _04023_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11524" *) _05718_;
  assign _04310_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11526" *) chn_in_rsci_d_mxwt[507];
  assign _04311_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11530" *) _04025_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11531" *) _05719_;
  assign _04312_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11533" *) chn_in_rsci_d_mxwt[475];
  assign _04313_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11537" *) _04027_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11538" *) _05720_;
  assign _04314_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11540" *) chn_in_rsci_d_mxwt[443];
  assign _04315_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11544" *) _04029_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11545" *) _05721_;
  assign _04316_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11547" *) chn_in_rsci_d_mxwt[411];
  assign _04317_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11551" *) _04031_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11552" *) _05722_;
  assign _04318_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11554" *) chn_in_rsci_d_mxwt[379];
  assign _04319_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11558" *) _04033_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11559" *) _05723_;
  assign _04320_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11561" *) chn_in_rsci_d_mxwt[347];
  assign _04321_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11565" *) _04035_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11566" *) _05724_;
  assign _04322_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11568" *) chn_in_rsci_d_mxwt[315];
  assign _04323_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11572" *) _04037_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11573" *) _05725_;
  assign _04324_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11575" *) chn_in_rsci_d_mxwt[283];
  assign _04325_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11579" *) _04039_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11580" *) _05726_;
  assign _04326_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11582" *) chn_in_rsci_d_mxwt[251];
  assign _04327_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11586" *) _04041_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11587" *) _05727_;
  assign _04328_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11589" *) chn_in_rsci_d_mxwt[219];
  assign _04329_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11593" *) _04043_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11594" *) _05728_;
  assign _04330_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11596" *) chn_in_rsci_d_mxwt[187];
  assign _04331_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11601" *) chn_in_rsci_d_mxwt[155];
  assign IsNaN_8U_23U_nor_4_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11605" *) _04045_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11606" *) _03878_;
  assign _04332_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11607" *) _04046_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11608" *) _05729_;
  assign _04333_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11610" *) chn_in_rsci_d_mxwt[123];
  assign _04334_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11614" *) _04048_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11615" *) _05730_;
  assign _04335_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11617" *) chn_in_rsci_d_mxwt[91];
  assign _04336_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11621" *) _04050_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11622" *) _05731_;
  assign _04337_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11624" *) chn_in_rsci_d_mxwt[59];
  assign _04338_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11628" *) _04052_;
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11629" *) _05732_;
  assign _04339_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11631" *) chn_in_rsci_d_mxwt[27];
  assign _00020_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11636" *) chn_idata_data_sva_1_27_0_1[27];
  assign _04341_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *) _05733_;
  assign _04342_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *) _05734_;
  assign _00021_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11642" *) chn_idata_data_sva_1_59_31_1[28];
  assign _04344_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *) _05735_;
  assign _04345_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *) _05736_;
  assign _00022_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11648" *) chn_idata_data_sva_1_91_63_1[28];
  assign _04347_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *) _05737_;
  assign _04348_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *) _05738_;
  assign _00023_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11654" *) chn_idata_data_sva_1_123_95_1[28];
  assign _04350_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *) _05739_;
  assign _04351_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *) _05740_;
  assign _00024_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11660" *) chn_idata_data_sva_1_155_127_1[28];
  assign _04353_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *) _05741_;
  assign _04354_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *) _05742_;
  assign _00025_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11666" *) chn_idata_data_sva_1_187_159_1[28];
  assign _04356_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *) _05743_;
  assign _04357_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *) _05744_;
  assign _00026_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11672" *) chn_idata_data_sva_1_219_191_1[28];
  assign _04359_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *) _05745_;
  assign _04360_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *) _05746_;
  assign _00027_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11678" *) chn_idata_data_sva_1_251_223_1[28];
  assign _04362_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *) _05747_;
  assign _04363_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *) _05748_;
  assign _00028_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11684" *) chn_idata_data_sva_1_283_255_1[28];
  assign _04365_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *) _05749_;
  assign _04366_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *) _05750_;
  assign _00029_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11690" *) chn_idata_data_sva_1_315_287_1[28];
  assign _04368_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *) _05751_;
  assign _04369_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *) _05752_;
  assign _00030_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11697" *) chn_idata_data_sva_1_347_319_1[28];
  assign _04371_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *) _05753_;
  assign _04372_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *) _05754_;
  assign _00031_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11704" *) chn_idata_data_sva_1_379_351_1[28];
  assign _04374_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *) _05755_;
  assign _04375_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *) _05756_;
  assign _00032_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11711" *) chn_idata_data_sva_1_411_383_1[28];
  assign _04377_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *) _05757_;
  assign _04378_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *) _05758_;
  assign _00033_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11718" *) chn_idata_data_sva_1_443_415_1[28];
  assign _04380_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *) _05759_;
  assign _04381_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *) _05760_;
  assign _00034_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11725" *) chn_idata_data_sva_1_475_447_1[28];
  assign _04383_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *) _05761_;
  assign _04384_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *) _05762_;
  assign _00035_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11732" *) chn_idata_data_sva_1_507_479_1[28];
  assign _04386_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *) _05763_;
  assign _04387_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *) _05764_;
  assign _04388_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11738" *) cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11759" *) _01502_;
  assign IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11765" *) _01503_;
  assign IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11771" *) _01504_;
  assign IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11777" *) _01505_;
  assign IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11783" *) _01506_;
  assign IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11789" *) _01507_;
  assign IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11795" *) _01508_;
  assign IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11801" *) _01509_;
  assign IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11810" *) _01510_;
  assign IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11816" *) _01511_;
  assign IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11825" *) _01512_;
  assign IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11831" *) _01513_;
  assign IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11837" *) _01514_;
  assign IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11843" *) _01515_;
  assign IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11849" *) _01516_;
  assign IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11855" *) _01517_;
  assign _00187_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11889" *) IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0[14];
  assign _00188_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11893" *) IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0[14];
  assign _04389_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11928" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[111];
  assign _04390_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11933" *) _03899_;
  assign _04391_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11935" *) _04070_;
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11935" *) _05319_;
  assign _00189_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11937" *) IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0[14];
  assign _00190_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11941" *) IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0[14];
  assign _04392_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11976" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[111];
  assign _04393_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11981" *) _03900_;
  assign _04394_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11983" *) _04071_;
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11983" *) _04857_;
  assign _04395_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12016" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[111];
  assign _04396_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12021" *) _03901_;
  assign _04397_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12023" *) _04072_;
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12023" *) _05320_;
  assign _00191_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12025" *) IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0[14];
  assign _00192_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12029" *) IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0[14];
  assign _04398_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12064" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[111];
  assign _04399_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12069" *) _03902_;
  assign _04400_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12071" *) _04073_;
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12071" *) _04860_;
  assign _00193_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12073" *) IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0[14];
  assign _00194_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12077" *) IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0[14];
  assign _04401_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12112" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[111];
  assign _04402_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12117" *) _03903_;
  assign _04403_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12119" *) _04074_;
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12119" *) _04863_;
  assign _04404_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12152" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[111];
  assign _04405_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12157" *) _03904_;
  assign _04406_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12159" *) _04075_;
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12159" *) _04861_;
  assign _04407_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12192" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[111];
  assign _04408_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12197" *) _03905_;
  assign _04409_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12199" *) _04076_;
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12199" *) _04859_;
  assign _00195_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12201" *) IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0[14];
  assign _00196_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12205" *) IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0[14];
  assign _04410_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12240" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[111];
  assign _04411_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12245" *) _03906_;
  assign _04412_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12247" *) _04077_;
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12247" *) _04864_;
  assign _00197_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12249" *) IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0[14];
  assign _00198_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12253" *) IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0[14];
  assign _04413_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12288" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[111];
  assign _04414_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12293" *) _03907_;
  assign _04415_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12295" *) _04078_;
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12295" *) _04866_;
  assign _04416_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12328" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[111];
  assign _04417_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12333" *) _03908_;
  assign _04418_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12335" *) _04079_;
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12335" *) _04865_;
  assign _00199_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12337" *) IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0[14];
  assign _00200_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12341" *) IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0[14];
  assign _04419_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12376" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[111];
  assign _04420_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12381" *) _03909_;
  assign _04421_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12383" *) _04080_;
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12383" *) _04869_;
  assign _00201_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12385" *) IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0[14];
  assign _00202_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12389" *) IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0[14];
  assign _04422_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12424" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[111];
  assign _04423_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12429" *) _03910_;
  assign _04424_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12431" *) _04081_;
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12431" *) _04873_;
  assign _04425_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12464" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[111];
  assign _04426_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12469" *) _03911_;
  assign _04427_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12471" *) _04082_;
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12471" *) _04871_;
  assign _04428_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12504" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[111];
  assign _04429_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12509" *) _03912_;
  assign _04430_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12511" *) _04083_;
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12511" *) _04868_;
  assign _04431_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12544" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[111];
  assign _04432_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12549" *) _03913_;
  assign _04433_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12551" *) _04084_;
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12551" *) _05324_;
  assign _04434_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12584" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[111];
  assign _04435_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12589" *) _03914_;
  assign _04436_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12591" *) _04085_;
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12591" *) _05318_;
  assign _04437_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12608" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[74];
  assign _04438_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12613" *) _03915_;
  assign _04439_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12615" *) _04086_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12615" *) _06787_;
  assign cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12617" *) _00139_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12619" *) _00140_;
  assign _04440_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12636" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[74];
  assign _04441_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12641" *) _03916_;
  assign _04442_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12643" *) _04087_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12643" *) _06818_;
  assign cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12645" *) _00141_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12647" *) _00142_;
  assign _04443_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12664" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[74];
  assign _04444_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12669" *) _03917_;
  assign _04445_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12671" *) _04088_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12671" *) _06849_;
  assign cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12673" *) _00143_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12675" *) _00144_;
  assign _04446_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12692" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[74];
  assign _04447_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12697" *) _03918_;
  assign _04448_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12699" *) _04089_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12699" *) _06880_;
  assign cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12701" *) _00145_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12703" *) _00146_;
  assign _04449_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12720" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[74];
  assign _04450_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12725" *) _03919_;
  assign _04451_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12727" *) _04090_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12727" *) _06911_;
  assign cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12729" *) _00147_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12731" *) _00148_;
  assign _04452_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12748" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[74];
  assign _04453_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12753" *) _03920_;
  assign _04454_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12755" *) _04091_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12755" *) _06942_;
  assign cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12757" *) _00149_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12759" *) _00150_;
  assign _04455_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12776" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[74];
  assign _04456_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12781" *) _03921_;
  assign _04457_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12783" *) _04092_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12783" *) _06973_;
  assign cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12785" *) _00151_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12787" *) _00152_;
  assign _04458_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12804" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[74];
  assign _04459_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12809" *) _03922_;
  assign _04460_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12811" *) _04093_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12811" *) _07004_;
  assign cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12813" *) _00153_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12815" *) _00154_;
  assign _04461_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12832" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[74];
  assign _04462_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12837" *) _03923_;
  assign _04463_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12839" *) _04094_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12839" *) _07035_;
  assign cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12841" *) _00155_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12843" *) _00156_;
  assign _04464_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12860" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[74];
  assign _04465_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12865" *) _03924_;
  assign _04466_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12867" *) _04095_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12867" *) _07066_;
  assign cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12869" *) _00157_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12871" *) _00158_;
  assign _04467_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12888" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[74];
  assign _04468_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12893" *) _03925_;
  assign _04469_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12895" *) _04096_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12895" *) _07097_;
  assign cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12897" *) _00159_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12899" *) _00160_;
  assign _04470_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12916" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[74];
  assign _04471_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12921" *) _03926_;
  assign _04472_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12923" *) _04097_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12923" *) _07128_;
  assign cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12925" *) _00161_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12927" *) _00162_;
  assign _04473_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12944" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[74];
  assign _04474_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12949" *) _03927_;
  assign _04475_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12951" *) _04098_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12951" *) _07159_;
  assign cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12953" *) _00163_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12955" *) _00164_;
  assign _04476_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12972" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[74];
  assign _04477_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12977" *) _03928_;
  assign _04478_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12979" *) _04099_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12979" *) _07190_;
  assign cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12981" *) _00165_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12983" *) _00166_;
  assign _04479_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13000" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[74];
  assign _04480_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13005" *) _03929_;
  assign _04481_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13007" *) _04100_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13007" *) _07221_;
  assign cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13009" *) _00167_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13011" *) _00168_;
  assign _04482_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13028" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[74];
  assign _04483_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13033" *) _03930_;
  assign _04484_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13035" *) _04101_;
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13035" *) _07252_;
  assign cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_22_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13037" *) _00169_;
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13039" *) _00170_;
  assign _04485_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13041" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16[4:1];
  assign _04486_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13050" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17[4:1];
  assign _04487_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13059" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18[4:1];
  assign _04488_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13068" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19[4:1];
  assign _04489_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13077" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20[4:1];
  assign _04490_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13086" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21[4:1];
  assign _04491_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13095" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22[4:1];
  assign _04492_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13104" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23[4:1];
  assign _04493_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13113" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24[4:1];
  assign _04494_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13122" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25[4:1];
  assign _04495_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13131" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26[4:1];
  assign _04496_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13140" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27[4:1];
  assign _04497_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13149" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28[4:1];
  assign _04498_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13158" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29[4:1];
  assign _04499_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13167" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30[4:1];
  assign _04500_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13176" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31[4:1];
  assign cvt_if_unequal_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13184" *) cvt_else_equal_tmp;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13193" *) _07333_;
  assign _04501_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13195" *) FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13207" *) _07334_;
  assign _04502_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13209" *) FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  assign cvt_else_nor_dfs = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13214" *) _07336_;
  assign cvt_else_equal_tmp_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13215" *) or_1431_nl;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13225" *) _07337_;
  assign _04503_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13227" *) FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13238" *) _07338_;
  assign _04504_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13240" *) FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13252" *) _07339_;
  assign _04505_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13254" *) FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13266" *) _07340_;
  assign _04506_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13268" *) FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13280" *) _07341_;
  assign _04507_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13282" *) FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13294" *) _07342_;
  assign _04508_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13296" *) FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13308" *) _07343_;
  assign _04509_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13310" *) FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13322" *) _07344_;
  assign _04510_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13324" *) FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13336" *) _07345_;
  assign _04511_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13338" *) FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13350" *) _07346_;
  assign _04512_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13352" *) FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13364" *) _07347_;
  assign _04513_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13366" *) FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13373" *) _07348_;
  assign _04514_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13375" *) cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13387" *) _07349_;
  assign _04515_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13389" *) FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13401" *) _07350_;
  assign _04516_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13403" *) FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  assign _04517_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13412" *) cfg_mode_eql_1_sva_6;
  assign _04518_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13416" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva[14:0];
  assign _04520_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13421" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva[14:0];
  assign _04522_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13426" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva[14:0];
  assign _04524_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13431" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva[14:0];
  assign _04526_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13436" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva[14:0];
  assign _04528_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13441" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva[14:0];
  assign _04530_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13446" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva[14:0];
  assign _04532_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13451" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva[14:0];
  assign _04534_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13456" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva[14:0];
  assign _04536_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13461" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva[14:0];
  assign _04538_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13466" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva[14:0];
  assign _04540_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13471" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva[14:0];
  assign _04542_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13476" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva[14:0];
  assign _04544_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13481" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva[14:0];
  assign _04546_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13486" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva[14:0];
  assign _04548_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13491" *) FpFloatToInt_16U_5U_10U_internal_int_24_1_sva[14:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13786" *) _04385_;
  assign _04550_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13790" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13794" *) _04382_;
  assign _04551_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13798" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13802" *) _04379_;
  assign _04552_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13806" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13810" *) _04376_;
  assign _04553_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13814" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13818" *) _04373_;
  assign _04554_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13822" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13826" *) _04370_;
  assign _04555_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13830" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13834" *) _04367_;
  assign _04556_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13838" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13842" *) _04364_;
  assign _04557_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13846" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13850" *) _04361_;
  assign _04558_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13854" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13858" *) _04358_;
  assign _04559_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13862" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13866" *) _04355_;
  assign _04560_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13870" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13874" *) _04352_;
  assign _04561_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13878" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13882" *) _04349_;
  assign _04562_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13886" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13890" *) _04346_;
  assign _04563_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13894" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13898" *) _04343_;
  assign _04564_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13902" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13906" *) _04340_;
  assign _04565_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13910" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2;
  assign _00203_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13912" *) IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0;
  assign _00204_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13916" *) IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0;
  assign _00205_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13920" *) IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0;
  assign _00206_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13924" *) IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0;
  assign _00207_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13928" *) IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0;
  assign _00208_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13932" *) IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0;
  assign _00209_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13936" *) IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0;
  assign _00210_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13940" *) IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0;
  assign _00211_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13944" *) IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0;
  assign _00212_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13948" *) IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0;
  assign _00213_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13952" *) IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0;
  assign _00214_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13956" *) IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0;
  assign _00215_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13960" *) IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0;
  assign _00216_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13964" *) IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0;
  assign _00217_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13968" *) IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0;
  assign _00218_[15:1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13972" *) IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13976" *) _07399_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13978" *) _07400_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13980" *) _07401_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13982" *) _07402_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13984" *) _07403_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13986" *) _07404_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13988" *) _07405_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13990" *) _07406_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13992" *) _07407_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13994" *) _07408_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13996" *) _07409_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13998" *) _07410_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14000" *) _07411_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14002" *) _07412_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14004" *) _07413_;
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14006" *) _07414_;
  assign cvt_asn_319 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14071" *) _07416_;
  assign _04566_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14072" *) cvt_unequal_tmp_21;
  assign _04567_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14107" *) and_dcpl_70;
  assign _04568_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14111" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign nor_8_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14115" *) or_4550_cse;
  assign _04569_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14121" *) and_tmp_12;
  assign nor_2056_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14121" *) _07420_;
  assign nor_2055_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14125" *) _07421_;
  assign not_tmp_119 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14127" *) _01542_;
  assign _04570_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14131" *) mux_tmp_120;
  assign nor_2054_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14131" *) _07422_;
  assign nor_2052_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14134" *) _07423_;
  assign _04571_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14136" *) mux_tmp_117;
  assign nor_2050_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14136" *) _07424_;
  assign _04572_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14139" *) and_tmp_33;
  assign nor_2049_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14139" *) _07425_;
  assign _04573_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14143" *) cfg_mode_eql_1_sva_4;
  assign nor_2029_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14143" *) _07426_;
  assign _04574_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14145" *) mux_188_nl;
  assign nand_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14145" *) _01543_;
  assign nor_2027_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14151" *) _07427_;
  assign _04575_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14153" *) mux_tmp_199;
  assign nor_2028_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14153" *) _07428_;
  assign _04576_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14156" *) _01544_;
  assign nor_2022_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14157" *) _07429_;
  assign nor_2021_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14159" *) _07430_;
  assign _00066_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14162" *) and_tmp_11;
  assign nor_50_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14164" *) or_4862_cse;
  assign _04577_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14174" *) _01546_;
  assign _00036_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14175" *) or_513_cse;
  assign _04578_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14184" *) mux_tmp_236;
  assign nor_2015_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14184" *) _07436_;
  assign _04579_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14186" *) mux_tmp_239;
  assign nor_2013_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14186" *) _07437_;
  assign _04580_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *) mux_344_cse;
  assign nor_2007_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *) or_2688_nl;
  assign nor_2009_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14192" *) or_2691_nl;
  assign nor_1995_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14195" *) or_2696_nl;
  assign nor_1997_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14198" *) or_2699_nl;
  assign not_tmp_270 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14200" *) _01548_;
  assign _04581_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14204" *) mux_tmp_259;
  assign nor_1988_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14204" *) _07446_;
  assign nor_1987_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14206" *) _07447_;
  assign nor_1983_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14212" *) _07448_;
  assign _04582_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14214" *) cvt_unequal_tmp_20;
  assign _00037_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14216" *) or_tmp_533;
  assign _00038_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14222" *) reg_cfg_proc_precision_1_sva_st_40_cse[1];
  assign _04583_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14225" *) mux_474_cse;
  assign nor_1975_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14225" *) or_2705_nl;
  assign nor_1977_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14227" *) or_2709_nl;
  assign _04584_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14229" *) and_tmp_50;
  assign nor_1974_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14229" *) _07454_;
  assign nor_1964_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14234" *) or_2714_nl;
  assign nor_1966_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14237" *) or_2717_nl;
  assign nor_151_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14239" *) or_400_cse_1;
  assign nor_1959_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14239" *) _07457_;
  assign nor_1955_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14242" *) _07459_;
  assign nor_1942_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14252" *) or_2723_nl;
  assign nor_1944_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14254" *) or_2727_nl;
  assign nor_1935_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14258" *) _07463_;
  assign nor_1922_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14267" *) or_2733_nl;
  assign nor_1924_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14269" *) or_2737_nl;
  assign _00039_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14271" *) cfg_proc_precision_1_sva_st_101[1];
  assign _04585_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14273" *) mux_tmp_415;
  assign nor_1919_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14273" *) _07466_;
  assign nor_1912_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14276" *) _07468_;
  assign _04586_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14278" *) mux_tmp_421;
  assign nor_1915_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14278" *) _07469_;
  assign _04587_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14284" *) mux_tmp_427;
  assign nor_1911_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14284" *) _07470_;
  assign _04588_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14286" *) mux_tmp_305;
  assign nor_1906_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14286" *) _07471_;
  assign _04589_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14288" *) mux_tmp_298;
  assign nor_1901_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14288" *) _07472_;
  assign _04590_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14290" *) mux_tmp_440;
  assign nor_1902_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14290" *) _07473_;
  assign nor_1892_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14293" *) or_2744_nl;
  assign nor_1894_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14295" *) or_2749_nl;
  assign nor_1891_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14299" *) _07476_;
  assign nor_1882_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14303" *) or_2754_nl;
  assign _04591_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14306" *) mux_1126_cse;
  assign nor_1884_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14306" *) or_2758_nl;
  assign nor_1872_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14309" *) _07481_;
  assign _04592_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14317" *) or_461_cse;
  assign nor_1858_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14321" *) or_2764_nl;
  assign nor_1860_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14323" *) or_2768_nl;
  assign nor_1851_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14326" *) _07487_;
  assign nor_1838_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14338" *) or_2774_nl;
  assign nor_1840_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14340" *) or_2778_nl;
  assign nor_1828_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14343" *) _07491_;
  assign _04593_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14347" *) _07492_;
  assign _04594_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14349" *) mux_tmp_565;
  assign nor_1827_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14349" *) _07493_;
  assign _04595_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14354" *) mux_tmp_577;
  assign nor_1815_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14354" *) _07494_;
  assign _04596_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14356" *) mux_tmp_578;
  assign nor_1816_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14356" *) _07495_;
  assign _04597_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14358" *) mux_tmp_579;
  assign nor_1817_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14358" *) _07496_;
  assign _04598_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14364" *) _01566_;
  assign _04599_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14368" *) mux_tmp_591;
  assign nor_1810_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14368" *) _07500_;
  assign _04600_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14370" *) mux_1460_cse;
  assign nor_1807_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14370" *) _07501_;
  assign _04601_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14374" *) _07502_;
  assign _04602_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14376" *) mux_tmp_600;
  assign nor_1803_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14376" *) _07503_;
  assign _04603_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14378" *) mux_tmp_601;
  assign nor_1804_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14378" *) _07504_;
  assign _04604_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14382" *) mux_tmp_612;
  assign nor_1795_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14382" *) _07505_;
  assign _04605_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14384" *) mux_tmp_613;
  assign nor_1796_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14384" *) _07506_;
  assign nor_1787_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14388" *) or_2784_nl;
  assign _04606_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14390" *) mux_382_cse;
  assign nor_1789_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14390" *) or_2789_nl;
  assign _04607_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14392" *) mux_1489_cse;
  assign nor_1780_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14392" *) _07509_;
  assign _04608_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14397" *) mux_tmp_638;
  assign nor_1774_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14397" *) _07510_;
  assign _04609_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14399" *) mux_tmp_639;
  assign nor_1775_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14399" *) _07511_;
  assign _04610_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14401" *) mux_tmp_640;
  assign nor_1776_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14401" *) _07512_;
  assign nor_1764_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14405" *) or_2796_nl;
  assign _04611_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14407" *) mux_417_cse;
  assign nor_1766_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14407" *) or_2802_nl;
  assign nor_1762_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14409" *) _07515_;
  assign _04612_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14413" *) _07516_;
  assign _04613_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14415" *) mux_tmp_678;
  assign nor_1748_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14415" *) _07517_;
  assign _04614_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14417" *) mux_tmp_679;
  assign nor_1749_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14417" *) _07518_;
  assign _04615_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14419" *) mux_tmp_680;
  assign nor_1750_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14419" *) _07519_;
  assign _04616_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14423" *) mux_tmp_692;
  assign nor_1738_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14423" *) _07520_;
  assign _04617_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14425" *) mux_tmp_693;
  assign nor_1739_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14425" *) _07521_;
  assign _04618_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14427" *) mux_tmp_694;
  assign nor_1740_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14427" *) _07522_;
  assign nor_1728_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14431" *) or_2809_nl;
  assign nor_1730_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14433" *) or_2815_nl;
  assign nor_1718_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14435" *) _07525_;
  assign _04619_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14437" *) mux_tmp_719;
  assign nor_1719_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14437" *) _07526_;
  assign _04620_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14441" *) _07527_;
  assign _04621_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14443" *) mux_tmp_723;
  assign nor_1711_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14443" *) _07528_;
  assign _04622_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14445" *) mux_tmp_724;
  assign nor_1712_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14445" *) _07529_;
  assign _04623_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14447" *) mux_tmp_725;
  assign nor_1713_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14447" *) _07530_;
  assign _04624_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14449" *) mux_tmp_726;
  assign nor_1714_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14449" *) _07531_;
  assign _04625_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14453" *) mux_tmp_739;
  assign nor_1699_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14453" *) _07532_;
  assign _04626_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14455" *) mux_tmp_740;
  assign nor_1700_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14455" *) _07533_;
  assign _04627_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14457" *) mux_tmp_741;
  assign nor_1701_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14457" *) _07534_;
  assign _04628_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14459" *) mux_tmp_742;
  assign nor_1702_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14459" *) _07535_;
  assign nor_1687_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14463" *) or_2823_nl;
  assign nor_1689_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14465" *) or_2830_nl;
  assign _04629_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14467" *) mux_tmp_658;
  assign nor_1685_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14467" *) _07538_;
  assign _04630_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14469" *) mux_tmp_765;
  assign nor_1686_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14469" *) _07539_;
  assign _04631_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14471" *) main_stage_v_3;
  assign or_tmp_1393 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14473" *) _01571_;
  assign nor_1672_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14485" *) or_1159_cse;
  assign nor_1545_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14485" *) _07541_;
  assign nor_1534_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14488" *) _07542_;
  assign _04632_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14490" *) mux_tmp_986;
  assign nor_1535_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14490" *) _07543_;
  assign _04633_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14494" *) _01572_;
  assign _04634_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14500" *) mux_tmp_987;
  assign nor_1486_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14500" *) _07545_;
  assign _04635_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14504" *) reg_chn_out_rsci_ld_core_psct_cse;
  assign _04636_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14507" *) mux_tmp_1038;
  assign nor_1487_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14507" *) _07549_;
  assign _04637_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14513" *) and_tmp_171;
  assign _00040_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14514" *) or_tmp_1650;
  assign _04638_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14522" *) and_tmp_168;
  assign nor_1464_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14522" *) _07552_;
  assign _04639_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14527" *) and_tmp_169;
  assign nor_1455_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14527" *) _07553_;
  assign _04640_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14540" *) mux_tmp_1100;
  assign nor_1446_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14540" *) _07558_;
  assign _04641_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14546" *) and_tmp_175;
  assign _00041_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14547" *) or_tmp_1780;
  assign nor_213_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14557" *) or_3538_cse;
  assign nor_1387_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14557" *) _07561_;
  assign _04642_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14559" *) mux_tmp_1196;
  assign nor_1388_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14559" *) _07562_;
  assign nand_202_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14561" *) _01575_;
  assign nor_1371_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14564" *) _07563_;
  assign _04643_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14566" *) mux_tmp_1225;
  assign nor_1372_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14566" *) _07564_;
  assign _04644_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14568" *) mux_tmp_1226;
  assign nor_1373_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14568" *) _07565_;
  assign _00042_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14573" *) or_tmp_2136;
  assign _00043_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14579" *) mux_1272_nl;
  assign nor_1320_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14581" *) or_tmp_2139;
  assign _00044_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14590" *) mux_1328_nl;
  assign _00045_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14595" *) mux_tmp_1332;
  assign _04645_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14607" *) _07478_;
  assign not_tmp_1709 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14615" *) _07569_;
  assign nand_tmp_48 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14616" *) _01576_;
  assign _04646_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14624" *) _07570_;
  assign _04647_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14625" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _00063_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14628" *) chn_in_rsci_bawt;
  assign nand_230_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14656" *) _01578_;
  assign _04648_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14675" *) chn_out_rsci_bawt;
  assign _04649_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14684" *) _03932_;
  assign or_dcpl_30 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14684" *) _01582_;
  assign nor_tmp_636 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14698" *) _07612_;
  assign not_tmp_2254 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14702" *) _01583_;
  assign _00070_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14733" *) and_tmp_225;
  assign nor_1063_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14733" *) _07614_;
  assign _04650_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14737" *) cfg_out_precision_1_sva_st_113[1];
  assign _04651_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14742" *) cfg_proc_precision_1_sva_st_65[0];
  assign _04652_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14750" *) and_dcpl_479;
  assign or_dcpl_151 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14750" *) _01589_;
  assign and_dcpl_444 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14751" *) or_425_cse;
  assign nor_1053_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14754" *) _07616_;
  assign _04653_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14764" *) and_tmp_165;
  assign nor_1025_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14764" *) _07617_;
  assign _04654_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14767" *) _03934_;
  assign or_dcpl_178 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14767" *) _01591_;
  assign _00069_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14777" *) mux_tmp_455;
  assign _04655_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14788" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl[8];
  assign _04656_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14789" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8];
  assign _04657_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14790" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _04658_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14791" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _04659_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14792" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _04660_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14793" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _04661_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14794" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _04662_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14795" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _04663_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14796" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _04664_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14797" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _04665_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14798" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _04666_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14799" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _04667_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14800" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _04668_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14801" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _04669_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14802" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _04670_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14803" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _04671_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14804" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign _04672_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14805" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign _04673_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14806" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _04674_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14807" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _04675_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14808" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _04676_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14809" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _04677_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14810" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _04678_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14811" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _04679_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14812" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign _04680_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14813" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign _04681_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14814" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _04682_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14815" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _04683_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14816" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign _04684_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14817" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _04685_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14818" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8];
  assign _04686_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14819" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8];
  assign _04687_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14849" *) cfg_proc_precision_rsci_d[1];
  assign _04688_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14854" *) _01603_;
  assign _04689_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14859" *) cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign _04690_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14862" *) _07644_;
  assign _04691_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14881" *) cfg_out_precision_1_sva_st_113[0];
  assign _04692_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14883" *) cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11];
  assign _04693_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14886" *) _07647_;
  assign nor_2040_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14973" *) or_5189_cse;
  assign _04694_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *) _07652_;
  assign _04695_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14983" *) _07654_;
  assign _04696_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *) _07657_;
  assign _00046_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14988" *) mux_tmp_2203;
  assign _04697_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14990" *) _01621_;
  assign _04698_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14992" *) and_dcpl_626;
  assign _00047_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15000" *) or_tmp;
  assign _00048_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15004" *) or_tmp_4080;
  assign _00049_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15010" *) or_tmp_4081;
  assign _00050_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15016" *) or_tmp_4082;
  assign _00051_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15021" *) or_tmp_4084;
  assign _00052_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15028" *) or_tmp_4086;
  assign _00053_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15033" *) or_tmp_4087;
  assign _00054_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15042" *) or_tmp_4092;
  assign _00055_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15046" *) or_tmp_4095;
  assign _00056_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15052" *) or_tmp_4097;
  assign _04699_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15056" *) FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6;
  assign _04700_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15057" *) IsNaN_5U_10U_land_2_lpi_1_dfm_4;
  assign _04701_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15058" *) FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  assign _04702_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15059" *) IsNaN_5U_10U_land_3_lpi_1_dfm_5;
  assign _04703_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15060" *) FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7;
  assign _04704_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15061" *) IsNaN_5U_10U_land_4_lpi_1_dfm_5;
  assign _04705_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15062" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7;
  assign _04706_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15063" *) IsNaN_5U_10U_land_5_lpi_1_dfm_5;
  assign _04707_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15064" *) FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7;
  assign _04708_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15065" *) IsNaN_5U_10U_land_6_lpi_1_dfm_5;
  assign _04709_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15066" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  assign _04710_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15067" *) IsNaN_5U_10U_land_7_lpi_1_dfm_6;
  assign _04711_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15068" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  assign _04712_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15069" *) IsNaN_5U_10U_land_8_lpi_1_dfm_5;
  assign _04713_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15070" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  assign _04714_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15071" *) IsNaN_5U_10U_land_9_lpi_1_dfm_5;
  assign _04715_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15072" *) FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7;
  assign _04716_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15073" *) IsNaN_5U_10U_land_lpi_1_dfm_5;
  assign _04717_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15074" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7;
  assign _04718_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15075" *) IsNaN_5U_10U_land_1_lpi_1_dfm_3;
  assign _04719_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15076" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  assign _04720_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15077" *) IsNaN_5U_10U_land_10_lpi_1_dfm_5;
  assign _04721_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15078" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  assign _04722_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15079" *) IsNaN_5U_10U_land_11_lpi_1_dfm_5;
  assign _04723_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15080" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7;
  assign _04724_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15081" *) IsNaN_5U_10U_land_12_lpi_1_dfm_5;
  assign _04725_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15082" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  assign _04726_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15083" *) IsNaN_5U_10U_land_13_lpi_1_dfm_5;
  assign _04727_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15084" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  assign _04728_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15085" *) IsNaN_5U_10U_land_14_lpi_1_dfm_6;
  assign _04729_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15086" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  assign _04730_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15087" *) IsNaN_5U_10U_land_15_lpi_1_dfm_3;
  assign _04731_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15094" *) main_stage_en_1;
  assign _04732_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15094" *) _01654_;
  assign _04733_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15369" *) mux_2302_nl;
  assign _04734_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15383" *) mux_2308_nl;
  assign _04735_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15396" *) mux_2314_nl;
  assign _04736_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15410" *) mux_2320_nl;
  assign _04737_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15424" *) mux_2327_nl;
  assign _04738_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15438" *) mux_2332_nl;
  assign _04739_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15452" *) mux_2338_nl;
  assign _04740_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15466" *) mux_2344_nl;
  assign _04741_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15480" *) mux_2349_nl;
  assign _04742_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15622" *) and_dcpl_105;
  assign _04743_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15630" *) main_stage_v_1_mx0c1;
  assign _04744_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15654" *) mux_8_nl;
  assign _04745_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15664" *) mux_10_nl;
  assign _04746_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15726" *) mux_14_nl;
  assign _04747_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15736" *) mux_16_nl;
  assign _04748_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15754" *) mux_19_nl;
  assign _04749_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15764" *) mux_21_nl;
  assign _04750_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15782" *) mux_24_nl;
  assign _04751_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15792" *) mux_26_nl;
  assign _04752_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15801" *) mux_28_nl;
  assign _04753_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15810" *) mux_30_nl;
  assign _04754_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15820" *) mux_32_nl;
  assign _04755_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15829" *) mux_34_nl;
  assign _04756_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15838" *) mux_36_nl;
  assign _04757_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15848" *) mux_38_nl;
  assign _04758_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15857" *) mux_41_nl;
  assign _04759_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15866" *) mux_42_nl;
  assign _04760_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15876" *) mux_44_nl;
  assign _04761_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15894" *) mux_47_nl;
  assign _04762_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15904" *) mux_49_nl;
  assign _04763_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15922" *) mux_52_nl;
  assign _04764_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15932" *) mux_54_nl;
  assign _04765_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15941" *) mux_56_nl;
  assign _04766_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15950" *) mux_58_nl;
  assign _04767_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15960" *) mux_60_nl;
  assign _04768_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15978" *) mux_63_nl;
  assign _04769_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15988" *) mux_65_nl;
  assign _04770_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16006" *) mux_68_nl;
  assign _04771_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16016" *) mux_70_nl;
  assign _04772_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16025" *) mux_72_nl;
  assign _04773_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16034" *) mux_74_nl;
  assign _04774_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16044" *) mux_76_nl;
  assign _04775_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16062" *) mux_79_nl;
  assign _04776_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16072" *) mux_81_nl;
  assign _04777_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16090" *) mux_84_nl;
  assign _04778_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16100" *) mux_86_nl;
  assign _04779_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16118" *) mux_89_nl;
  assign _04780_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16128" *) mux_91_nl;
  assign _04781_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7];
  assign _04782_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16305" *) _01745_;
  assign _04783_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _04784_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16313" *) _01748_;
  assign _04785_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _04786_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16321" *) _01751_;
  assign _04787_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _04788_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16329" *) _01754_;
  assign _04789_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _04790_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16337" *) _01757_;
  assign _04791_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _04792_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16345" *) _01760_;
  assign _04793_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _04794_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16353" *) _01763_;
  assign _04795_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _04796_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16361" *) _01766_;
  assign _04797_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _04798_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16369" *) _01769_;
  assign _04799_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _04800_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16377" *) _01772_;
  assign _04801_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _04802_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16385" *) _01775_;
  assign _04803_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _04804_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16394" *) _01778_;
  assign _04805_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _04806_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16402" *) _01781_;
  assign _04807_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _04808_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16410" *) _01784_;
  assign _04809_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _04810_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16418" *) _01787_;
  assign _04811_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7];
  assign _04812_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16426" *) _01790_;
  assign _04813_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16523" *) main_stage_v_2_mx0c1;
  assign _04814_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16667" *) _04152_;
  assign _04815_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *) _01796_;
  assign _04816_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *) _07696_;
  assign _04817_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16669" *) _04153_;
  assign _04818_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *) _01797_;
  assign _04819_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *) _07697_;
  assign _04820_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16671" *) _04154_;
  assign _04821_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *) _01798_;
  assign _04822_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *) _07698_;
  assign _04823_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16673" *) _04155_;
  assign _04824_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *) _01799_;
  assign _04825_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *) _07699_;
  assign _04826_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16675" *) _04156_;
  assign _04827_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *) _01800_;
  assign _04828_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *) _07700_;
  assign _04829_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16677" *) _04157_;
  assign _04830_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *) _01801_;
  assign _04831_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *) _07701_;
  assign _04832_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16679" *) _04158_;
  assign _04833_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *) _01802_;
  assign _04834_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *) _07702_;
  assign _04835_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16681" *) _04159_;
  assign _04836_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *) _01803_;
  assign _04837_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *) _07703_;
  assign _04838_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16683" *) _04160_;
  assign _04839_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *) _01804_;
  assign _04840_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *) _07704_;
  assign _04841_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16685" *) _04161_;
  assign _04842_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *) _01805_;
  assign _04843_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *) _07705_;
  assign _04844_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16687" *) _04162_;
  assign _04845_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *) _01806_;
  assign _04846_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *) _07706_;
  assign _04847_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16689" *) _04163_;
  assign _04848_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *) _01807_;
  assign _04849_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *) _07707_;
  assign _04850_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16691" *) _04164_;
  assign _04851_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *) _01808_;
  assign _04852_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *) _07708_;
  assign _04853_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16792" *) mux_167_nl;
  assign _04854_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16942" *) mux_191_nl;
  assign _04855_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16961" *) mux_192_nl;
  assign _04856_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17000" *) mux_tmp_245;
  assign _04858_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17257" *) _07726_;
  assign _04862_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17443" *) _07730_;
  assign _04867_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *) mux_tmp_585;
  assign _04870_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17838" *) _07738_;
  assign _04872_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17894" *) _07740_;
  assign _04874_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17955" *) main_stage_v_3_mx0c1;
  assign _04875_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18532" *) mux_899_nl;
  assign _04876_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18755" *) _07784_;
  assign _04877_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18760" *) _07785_;
  assign _04878_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18763" *) _07786_;
  assign _04879_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18766" *) _07787_;
  assign _04880_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18769" *) _07788_;
  assign _04881_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18772" *) _07789_;
  assign _04882_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18775" *) _07790_;
  assign _04883_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18778" *) _07791_;
  assign _04884_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18781" *) _07792_;
  assign _04885_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18784" *) _07793_;
  assign _04886_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18787" *) _07794_;
  assign _04887_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18790" *) _07795_;
  assign _04888_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18793" *) _07796_;
  assign _04889_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18796" *) _07797_;
  assign _04890_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18799" *) _07798_;
  assign _04891_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18802" *) _07799_;
  assign _04892_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18882" *) _07800_;
  assign _04893_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18883" *) mux_954_nl;
  assign _04894_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18899" *) _07801_;
  assign _04895_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18900" *) mux_964_nl;
  assign _04896_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18938" *) mux_995_nl;
  assign _04897_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18959" *) _07802_;
  assign _04898_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18988" *) cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl[4];
  assign _04899_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18989" *) _02055_;
  assign _04900_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18990" *) _07803_;
  assign _04901_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18997" *) cfg_mode_eql_1_sva_5;
  assign _04902_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18998" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  assign _04903_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18999" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign _04904_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19028" *) mux_1018_nl;
  assign _04905_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19038" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _04906_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19039" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _04907_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19060" *) cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign _04908_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19061" *) _02089_;
  assign _04909_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19062" *) _07805_;
  assign _04910_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19063" *) cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign _04911_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19064" *) _02091_;
  assign _04912_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19065" *) _07806_;
  assign _04913_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19073" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _04914_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19074" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _04915_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19104" *) mux_1054_nl;
  assign _04916_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19115" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _04917_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19116" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign _04918_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19135" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _04919_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19166" *) mux_1077_nl;
  assign _04920_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19177" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _04921_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19178" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign _04922_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19197" *) mux_1091_nl;
  assign _04923_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19208" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _04924_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19209" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign _04925_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19228" *) mux_1116_nl;
  assign _04926_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19239" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _04927_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19240" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign _04928_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19259" *) cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign _04929_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19260" *) _02196_;
  assign _04930_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19261" *) _07808_;
  assign _04931_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19269" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _04932_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19270" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _04933_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19310" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _04934_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19311" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign _04935_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19329" *) mux_1163_nl;
  assign _04936_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19341" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _04937_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19342" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign _04938_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19360" *) mux_1179_nl;
  assign _04939_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19372" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _04940_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19373" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign _04941_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19405" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _04942_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19406" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign _04943_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19424" *) mux_1204_nl;
  assign _04944_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19432" *) mux_1213_nl;
  assign _04945_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19442" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _04946_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19443" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign _04947_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19461" *) cfg_out_precision_1_sva_st_149[1];
  assign _04948_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19492" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _04949_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19493" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign _04950_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19513" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2;
  assign _04951_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19514" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign _04952_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19576" *) _07809_;
  assign _04953_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19577" *) _07810_;
  assign _04954_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19586" *) mux_2249_nl;
  assign _04955_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19805" *) mux_1533_nl;
  assign _04956_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20069" *) mux_1569_nl;
  assign _04957_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *) mux_tmp_6;
  assign _04958_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20088" *) mux_1573_nl;
  assign _04959_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20107" *) mux_1577_nl;
  assign _04960_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20126" *) mux_1581_nl;
  assign _04961_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20145" *) mux_1585_nl;
  assign _04962_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20164" *) mux_1589_nl;
  assign _04963_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20202" *) mux_1595_nl;
  assign _04964_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20221" *) mux_1599_nl;
  assign _04965_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20240" *) mux_1603_nl;
  assign _04966_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20278" *) mux_1609_nl;
  assign _04967_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20297" *) mux_1613_nl;
  assign _04968_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20316" *) mux_1617_nl;
  assign _04969_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20335" *) mux_1621_nl;
  assign _04970_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20354" *) mux_1625_nl;
  assign _04971_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20581" *) cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign _04972_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20583" *) cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign _04973_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20585" *) cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign _04974_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20587" *) cvt_1_IntSaturation_17U_16U_else_if_acc_nl[2];
  assign _04975_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20589" *) cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl[2];
  assign _04976_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20591" *) cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign _04977_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20593" *) cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign _04978_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20595" *) cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign _04979_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20597" *) cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign _04980_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20599" *) cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign _04981_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20601" *) cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign _04982_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20603" *) cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign _04983_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20605" *) cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign _04984_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20607" *) cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign _04985_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20609" *) cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign _04986_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *) _07882_;
  assign _04987_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *) _07884_;
  assign _04988_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *) _07888_;
  assign _04989_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *) _07891_;
  assign _04990_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *) _07895_;
  assign _04991_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *) _07898_;
  assign _04992_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *) _07902_;
  assign _04993_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *) _07903_;
  assign _04994_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20903" *) _07907_;
  assign _04995_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20913" *) _07910_;
  assign _04996_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *) _07914_;
  assign _04997_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *) _07915_;
  assign _04998_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *) _07919_;
  assign _04999_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *) _07920_;
  assign _05000_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *) _07927_;
  assign _05001_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *) _07930_;
  assign _05002_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20978" *) _07934_;
  assign _05003_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20988" *) _07937_;
  assign _05004_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *) _07942_;
  assign _05005_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *) _07944_;
  assign _05006_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *) _07948_;
  assign _05007_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *) _07949_;
  assign _05008_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *) _07956_;
  assign _05009_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *) _07959_;
  assign _05010_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *) _07964_;
  assign _05011_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *) _07968_;
  assign _05012_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *) _07974_;
  assign _00071_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21083" *) mux_1142_cse;
  assign _05013_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *) _07976_;
  assign _05014_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *) _07983_;
  assign _05015_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *) _07986_;
  assign _05016_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *) _07991_;
  assign _05017_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *) _07995_;
  assign _05018_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21152" *) mux_1415_nl;
  assign _05019_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *) or_dcpl_386;
  assign _05020_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *) mux_tmp_114;
  assign _05021_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21179" *) _07997_;
  assign _05022_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *) or_dcpl_16;
  assign _05023_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *) mux_tmp_122;
  assign nor_1992_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21234" *) or_tmp_3032;
  assign _05024_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *) _08002_;
  assign _05025_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *) _08006_;
  assign _05026_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *) _08010_;
  assign _05027_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *) _08014_;
  assign _05028_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *) _08018_;
  assign _05029_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *) _08022_;
  assign _05030_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *) _08026_;
  assign _05031_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *) _08030_;
  assign _05032_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *) _08034_;
  assign _05033_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *) _08038_;
  assign _05034_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *) _08042_;
  assign _05035_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *) _08046_;
  assign _05036_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *) _08050_;
  assign _05037_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *) _08054_;
  assign _05038_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *) _08058_;
  assign _05039_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *) _08062_;
  assign _05040_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21417" *) or_tmp_4102;
  assign _05041_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21420" *) or_5175_tmp;
  assign _05042_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21423" *) or_5177_tmp;
  assign _05043_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21426" *) or_5181_tmp;
  assign _05044_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21462" *) or_5174_tmp;
  assign _05045_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21467" *) or_5176_tmp;
  assign _05046_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21474" *) or_5178_tmp;
  assign _05047_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21480" *) or_5179_tmp;
  assign _05048_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21485" *) or_5180_tmp;
  assign _05049_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21493" *) or_5182_tmp;
  assign _05050_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21499" *) or_5183_tmp;
  assign _05051_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21504" *) or_5184_tmp;
  assign _05052_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21512" *) or_5185_tmp;
  assign _05053_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21517" *) or_5186_tmp;
  assign _05054_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21522" *) or_5188_tmp;
  assign _05055_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21528" *) or_5187_tmp;
  assign _00057_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21533" *) mux_2361_nl;
  assign _05056_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21547" *) cvt_1_IntSaturation_17U_8U_else_if_acc_nl[10];
  assign _05057_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21574" *) cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign _05058_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21600" *) cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign _05059_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21627" *) cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign _05060_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21654" *) cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign _05061_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21681" *) cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign _05062_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21708" *) cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign _05063_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21735" *) cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign _05064_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21762" *) cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign _05065_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21789" *) cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign _05066_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21816" *) cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign _05067_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21843" *) cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign _05068_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21870" *) cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign _05069_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21920" *) cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign _05070_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21935" *) cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl[10];
  assign nor_2081_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *) _08066_;
  assign _05071_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21963" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2;
  assign nor_2082_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21965" *) _08069_;
  assign _05072_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21967" *) or_4524_cse;
  assign _05073_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21970" *) _08070_;
  assign _05074_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21971" *) _08071_;
  assign _05075_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21981" *) _02659_;
  assign _05076_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21982" *) _08072_;
  assign nor_2075_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22006" *) _08085_;
  assign _05077_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22008" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign nor_2076_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22010" *) _08088_;
  assign nor_2073_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22029" *) _08099_;
  assign _05078_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22031" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign nor_2074_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22033" *) _08102_;
  assign nor_2071_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22052" *) _08113_;
  assign _05079_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22054" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign nor_2072_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22056" *) _08116_;
  assign _05080_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22075" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign nand_235_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22096" *) _02662_;
  assign _05081_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22104" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign nand_234_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22125" *) _02664_;
  assign nand_233_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22147" *) _02666_;
  assign nor_2069_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22155" *) _08170_;
  assign _05082_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22157" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign nor_2070_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22159" *) _08173_;
  assign nor_2067_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22178" *) _08184_;
  assign _05083_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22180" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign nor_2068_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22182" *) _08187_;
  assign _05084_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22201" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign nand_232_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22224" *) _02668_;
  assign nor_2065_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22232" *) _08214_;
  assign _05085_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22234" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign nor_2066_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22236" *) _08217_;
  assign nor_2063_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22255" *) _08228_;
  assign _05086_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22257" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign nor_2064_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22259" *) _08231_;
  assign _05087_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22278" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign nand_231_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22301" *) _02670_;
  assign nor_2061_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22309" *) _08258_;
  assign _05088_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22311" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign nor_2062_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22313" *) _08261_;
  assign nor_2059_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22332" *) _08272_;
  assign _05089_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22334" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign nor_2060_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22336" *) _08275_;
  assign nor_2057_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22355" *) _08286_;
  assign _05090_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22357" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2;
  assign nor_2058_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22359" *) _08289_;
  assign _00219_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22482" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0;
  assign _00219_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22483" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign nor_2048_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22486" *) _08299_;
  assign _00220_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22488" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0;
  assign _00220_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22489" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00221_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22491" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0;
  assign _00221_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22492" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00222_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22494" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0;
  assign _00222_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22495" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00223_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22497" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0;
  assign _00223_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22498" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00224_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22501" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0;
  assign _00224_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22502" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00225_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22504" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0;
  assign _00225_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22505" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00226_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22507" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0;
  assign _00226_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22508" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00227_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22511" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00227_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22511" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0;
  assign _00228_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22514" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00228_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22514" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0;
  assign _00229_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22517" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00229_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22517" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0;
  assign _00230_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22520" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00230_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22520" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0;
  assign _00231_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22522" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0;
  assign _00231_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22523" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00232_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22526" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00232_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22526" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0;
  assign _00233_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22529" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00233_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22529" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0;
  assign _00234_[2:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22534" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0[3:1];
  assign _00234_[3] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22534" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0;
  assign nor_2020_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22543" *) _08300_;
  assign nor_2016_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22550" *) _08301_;
  assign nor_2017_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22553" *) _08303_;
  assign nor_1993_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22586" *) _08306_;
  assign _05091_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22590" *) and_tmp_67;
  assign nor_1991_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22590" *) _08307_;
  assign _05092_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22594" *) mux_tmp_294;
  assign nor_1984_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22594" *) _08308_;
  assign _05093_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22597" *) mux_tmp_299;
  assign nor_1985_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22597" *) _08309_;
  assign nor_1962_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22625" *) _08312_;
  assign _00059_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22626" *) or_tmp_218;
  assign _05094_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22634" *) mux_tmp_351;
  assign nor_1951_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22634" *) _08313_;
  assign _05095_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22637" *) mux_tmp_356;
  assign nor_1952_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22637" *) _08314_;
  assign _05096_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22650" *) mux_tmp_386;
  assign nor_1931_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22650" *) _08315_;
  assign _05097_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22653" *) mux_tmp_391;
  assign nor_1932_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22653" *) _08316_;
  assign _05098_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22666" *) mux_tmp_422;
  assign nor_1907_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22666" *) _08317_;
  assign _05099_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22669" *) mux_tmp_428;
  assign nor_1908_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22669" *) _08318_;
  assign _05100_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22702" *) mux_tmp_481;
  assign nor_1868_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22702" *) _08319_;
  assign _05101_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22705" *) mux_tmp_487;
  assign nor_1869_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22705" *) _08320_;
  assign _05102_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22720" *) mux_tmp_519;
  assign nor_1847_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22720" *) _08321_;
  assign _05103_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22723" *) mux_tmp_525;
  assign nor_1848_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22723" *) _08322_;
  assign _05104_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22738" *) mux_tmp_560;
  assign nor_1822_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22738" *) _08323_;
  assign _05105_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22741" *) mux_tmp_566;
  assign nor_1823_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22741" *) _08324_;
  assign _05106_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22747" *) mux_tmp_580;
  assign nor_1814_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22747" *) _08325_;
  assign _05107_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22753" *) mux_tmp_592;
  assign nor_1809_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22753" *) _08326_;
  assign _05108_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22758" *) mux_tmp_597;
  assign nor_1800_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22758" *) _08328_;
  assign _05109_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22761" *) mux_tmp_602;
  assign nor_1801_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22761" *) _08329_;
  assign nor_1793_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22765" *) _08330_;
  assign _05110_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22768" *) mux_tmp_614;
  assign nor_1794_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22768" *) _08331_;
  assign _05111_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22781" *) mux_tmp_641;
  assign nor_1773_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22781" *) _08332_;
  assign _05112_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22798" *) mux_tmp_634;
  assign nor_1745_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22798" *) _08334_;
  assign _05113_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22801" *) mux_tmp_681;
  assign nor_1746_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22801" *) _08335_;
  assign _05114_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22807" *) mux_tmp_695;
  assign nor_1737_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22807" *) _08336_;
  assign _05115_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22811" *) or_tmp_3840;
  assign nor_2290_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22811" *) _08337_;
  assign _05116_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22823" *) mux_tmp_720;
  assign nor_1708_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22823" *) _08339_;
  assign _05117_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22826" *) mux_tmp_727;
  assign nor_1709_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22826" *) _08340_;
  assign nor_1697_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22830" *) _08341_;
  assign _05118_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22833" *) mux_tmp_743;
  assign nor_1698_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22833" *) _08342_;
  assign _05119_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22837" *) or_tmp_3849;
  assign nor_2287_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22837" *) _08343_;
  assign _00060_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22842" *) or_tmp_306;
  assign _00175_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22846" *) IntShiftRightSat_49U_6U_17U_o_16_10_sva_2;
  assign _00175_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22847" *) IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2[14:6];
  assign _00176_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22849" *) IntShiftRightSat_49U_6U_17U_o_16_2_sva_2;
  assign _00176_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22850" *) IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2[14:6];
  assign _00177_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22852" *) IntShiftRightSat_49U_6U_17U_o_16_4_sva_2;
  assign _00177_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22853" *) IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2[14:6];
  assign _00178_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22855" *) IntShiftRightSat_49U_6U_17U_o_16_6_sva_2;
  assign _00178_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22856" *) IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2[14:6];
  assign _00179_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22858" *) IntShiftRightSat_49U_6U_17U_o_16_7_sva_2;
  assign _00179_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22859" *) IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2[14:6];
  assign _00180_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22861" *) IntShiftRightSat_49U_6U_17U_o_16_sva_2;
  assign _00180_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22862" *) IntShiftRightSat_49U_6U_17U_o_15_1_sva_2[14:6];
  assign _00181_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22864" *) IntShiftRightSat_49U_6U_17U_o_16_8_sva_2;
  assign _00181_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22865" *) IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2[14:6];
  assign _00182_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22867" *) IntShiftRightSat_49U_6U_17U_o_16_15_sva_2;
  assign _00182_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22868" *) IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2[14:6];
  assign _00183_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22870" *) IntShiftRightSat_49U_6U_17U_o_16_13_sva_2;
  assign _00183_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22871" *) IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2[14:6];
  assign _00184_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22873" *) IntShiftRightSat_49U_6U_17U_o_16_11_sva_2;
  assign _00184_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22874" *) IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2[14:6];
  assign _00185_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22876" *) IntShiftRightSat_49U_6U_17U_o_16_12_sva_2;
  assign _00185_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22877" *) IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2[14:6];
  assign _05120_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22879" *) _08344_;
  assign nor_1667_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22880" *) _08347_;
  assign _05121_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22882" *) chn_idata_data_sva_2_47_31_1[0];
  assign nor_1670_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22883" *) _08349_;
  assign nand_208_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22887" *) _02696_;
  assign _05122_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22890" *) _08350_;
  assign nor_1671_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22893" *) _08351_;
  assign _05123_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22895" *) cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl[11];
  assign nor_1665_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22896" *) _08353_;
  assign _05124_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22899" *) _08354_;
  assign _05125_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22901" *) mux_813_cse;
  assign nand_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22901" *) _02697_;
  assign nor_1658_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22906" *) _08357_;
  assign _05126_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22909" *) _08358_;
  assign nand_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22911" *) _02698_;
  assign _05127_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22916" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp;
  assign _05128_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *) cvt_1_FpMantRNE_17U_11U_else_and_tmp;
  assign _05129_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *) _08361_;
  assign _05130_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *) _08362_;
  assign nand_4_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *) _02699_;
  assign nor_1653_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22923" *) _08364_;
  assign nor_1655_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22927" *) _08367_;
  assign _05131_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22931" *) cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign nor_1652_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22932" *) _08370_;
  assign _05132_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22935" *) _08371_;
  assign nand_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22937" *) _02700_;
  assign _05133_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22947" *) cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign nor_1649_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22948" *) _08374_;
  assign _05134_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22951" *) _08375_;
  assign nand_6_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22953" *) _02701_;
  assign _05135_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22957" *) chn_idata_data_sva_2_143_127_1[0];
  assign _05136_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22962" *) IsNaN_5U_10U_land_4_lpi_1_dfm_4;
  assign _05137_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22965" *) cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign nor_1646_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22966" *) _08378_;
  assign _05138_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22969" *) _08379_;
  assign nand_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22971" *) _02705_;
  assign _05139_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22975" *) chn_idata_data_sva_2_175_159_1[0];
  assign nor_1636_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22976" *) _08383_;
  assign _05140_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22977" *) _08384_;
  assign nor_1637_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22978" *) _08387_;
  assign nor_1640_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22982" *) _08389_;
  assign nand_206_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22986" *) _02706_;
  assign _05141_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22989" *) _08390_;
  assign nor_1641_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22992" *) _08391_;
  assign _05142_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22994" *) cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign nor_1634_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22995" *) _08393_;
  assign _05143_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22998" *) _08394_;
  assign nand_9_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23000" *) _02707_;
  assign nor_1625_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *) _08399_;
  assign nor_1628_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23010" *) _08402_;
  assign _05144_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23016" *) cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign nor_1623_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23017" *) _08404_;
  assign _05145_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23020" *) _08405_;
  assign nand_10_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23022" *) _02708_;
  assign _05146_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23026" *) cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign nor_1620_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23027" *) _08408_;
  assign _05147_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23030" *) _08409_;
  assign nand_11_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23032" *) _02709_;
  assign _05148_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23036" *) chn_idata_data_sva_2_495_479_1[0];
  assign nor_1610_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23037" *) _08413_;
  assign _05149_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23038" *) _08414_;
  assign nor_1611_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23039" *) _08417_;
  assign nor_1614_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23043" *) _08419_;
  assign nand_205_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23047" *) _02710_;
  assign _05150_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23050" *) _08420_;
  assign nor_1615_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23053" *) _08421_;
  assign _05151_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23055" *) cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign nor_1608_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23056" *) _08423_;
  assign _05152_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23059" *) _08424_;
  assign nand_13_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23061" *) _02711_;
  assign _05153_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23065" *) chn_idata_data_sva_2_239_223_1[0];
  assign nor_1598_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23066" *) _08428_;
  assign _05154_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23067" *) _08429_;
  assign nor_1599_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23068" *) _08432_;
  assign nor_1602_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23072" *) _08434_;
  assign nand_204_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23076" *) _02712_;
  assign _05155_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23079" *) _08435_;
  assign nor_1603_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23082" *) _08436_;
  assign _05156_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23084" *) cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign nor_1596_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23085" *) _08438_;
  assign _05157_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23088" *) _08439_;
  assign nand_15_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23090" *) _02713_;
  assign nand_16_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23094" *) _02714_;
  assign _05158_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23095" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_5;
  assign _05159_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *) _08442_;
  assign nand_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *) _02715_;
  assign _05160_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *) cvt_6_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _05161_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *) _08443_;
  assign _05162_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *) or_1720_cse_1;
  assign _05163_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *) _08444_;
  assign _05164_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *) _02716_;
  assign nor_1584_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23112" *) or_1196_cse;
  assign _05165_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23113" *) cvt_15_FpMantRNE_17U_11U_else_and_3_svs;
  assign _05166_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23113" *) _08449_;
  assign _05167_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23114" *) mux_tmp_416;
  assign _05168_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23117" *) _08451_;
  assign _05169_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23119" *) cvt_15_FpMantRNE_17U_11U_else_and_3_tmp;
  assign nor_1585_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23122" *) _08453_;
  assign nor_1588_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23129" *) _08458_;
  assign _05170_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23132" *) or_4788_cse;
  assign _05171_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23134" *) cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign nor_1583_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23135" *) _08460_;
  assign _05172_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23138" *) _08461_;
  assign nand_21_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23140" *) _02717_;
  assign _05173_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23144" *) chn_idata_data_sva_2_271_255_1[0];
  assign nor_1574_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23145" *) _08465_;
  assign _05174_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23146" *) _08466_;
  assign nor_1575_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23147" *) _08469_;
  assign nor_1577_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23151" *) _08471_;
  assign nor_1578_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23153" *) _08473_;
  assign nand_22_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23160" *) _02718_;
  assign nor_1579_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23162" *) _08475_;
  assign _05175_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23164" *) cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign nor_1572_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23165" *) _08477_;
  assign _05176_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23168" *) _08478_;
  assign nand_23_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23170" *) _02719_;
  assign _05177_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23174" *) cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign nor_1569_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23175" *) _08481_;
  assign _05178_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23178" *) _08482_;
  assign nand_24_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23180" *) _02720_;
  assign _05179_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23184" *) cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign nor_1566_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23185" *) _08485_;
  assign _05180_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23188" *) _08486_;
  assign nand_25_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23190" *) _02721_;
  assign _05181_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23194" *) cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign nor_1563_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23195" *) _08489_;
  assign _05182_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23198" *) _08490_;
  assign nand_26_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23200" *) _02722_;
  assign nor_1557_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23304" *) _08495_;
  assign _05183_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23308" *) _08499_;
  assign _05184_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23309" *) _08500_;
  assign nor_1558_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23309" *) _08501_;
  assign _00186_[10] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23311" *) IntShiftRightSat_49U_6U_17U_o_16_14_sva_2;
  assign _00186_[8:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23312" *) IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2[14:6];
  assign _05185_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23316" *) and_tmp_166;
  assign nor_1555_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23316" *) _08502_;
  assign _05186_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *) _08505_;
  assign _05187_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *) _08506_;
  assign nor_1547_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *) _08507_;
  assign _05188_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *) _08509_;
  assign _05189_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *) _08510_;
  assign nor_1548_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *) _08511_;
  assign _05190_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *) _08513_;
  assign _05191_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *) _08514_;
  assign nor_1537_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *) _08515_;
  assign _05192_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *) _08517_;
  assign _05193_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *) _08518_;
  assign nor_1538_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *) _08519_;
  assign _05194_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *) _08521_;
  assign _05195_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *) _08522_;
  assign nor_1526_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *) _08523_;
  assign _05196_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *) _08525_;
  assign _05197_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *) _08526_;
  assign nor_1527_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *) _08527_;
  assign nor_1519_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23356" *) _08530_;
  assign nor_1521_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *) _08534_;
  assign _05198_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23360" *) _03981_;
  assign _05199_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *) or_1202_cse;
  assign nor_2461_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *) _08538_;
  assign nor_1510_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23369" *) _08540_;
  assign nor_1511_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23371" *) _08542_;
  assign _05200_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23380" *) cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign _05201_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23380" *) _02724_;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23381" *) _08543_;
  assign _05202_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23382" *) mux_tmp_944;
  assign nor_1508_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23382" *) _08544_;
  assign _05203_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23387" *) _03982_;
  assign _05204_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *) _08548_;
  assign _05205_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *) _02727_;
  assign nor_2457_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *) _08549_;
  assign _05206_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23406" *) _03983_;
  assign _05207_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *) _08553_;
  assign _05208_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *) _02729_;
  assign nor_2453_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *) _08554_;
  assign _05209_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23420" *) _03984_;
  assign _05210_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *) _08559_;
  assign _05211_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *) _02731_;
  assign nor_2449_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *) _08560_;
  assign _05212_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23429" *) _03985_;
  assign _05213_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *) _08564_;
  assign _05214_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *) _02733_;
  assign nor_2445_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *) _08565_;
  assign nor_1465_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23439" *) _08567_;
  assign nor_1466_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23441" *) _08569_;
  assign _05215_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23447" *) _03986_;
  assign _05216_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *) _08574_;
  assign _05217_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *) _02735_;
  assign nor_2441_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *) _08575_;
  assign _05218_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23459" *) _03987_;
  assign _05219_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *) _08580_;
  assign _05220_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *) _02737_;
  assign nor_2437_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *) _08581_;
  assign _05221_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23475" *) _03988_;
  assign _05222_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *) _08586_;
  assign _05223_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *) _02739_;
  assign nor_2433_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *) _08587_;
  assign nor_1433_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23491" *) _08591_;
  assign _05224_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23493" *) _03989_;
  assign _05225_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *) _08595_;
  assign _05226_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *) _02741_;
  assign nor_2429_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *) _08596_;
  assign _05227_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23504" *) _03990_;
  assign _05228_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *) _08599_;
  assign _05229_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *) _02744_;
  assign nor_2425_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *) _08600_;
  assign _05230_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23516" *) _03991_;
  assign _05231_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *) _08603_;
  assign _05232_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *) _02746_;
  assign _05233_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *) _08604_;
  assign _05234_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23530" *) _02747_;
  assign nor_1403_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23530" *) _08605_;
  assign _05235_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23537" *) _03992_;
  assign _05236_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *) _08608_;
  assign _05237_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *) _02749_;
  assign _05238_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *) _08609_;
  assign _05239_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23546" *) _03993_;
  assign _05240_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *) _08612_;
  assign _05241_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *) _02752_;
  assign nor_2411_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *) _08613_;
  assign _05242_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23556" *) _08614_;
  assign nand_45_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23556" *) _02753_;
  assign nand_201_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23557" *) _02755_;
  assign _05243_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23562" *) _08615_;
  assign nand_46_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23562" *) _02756_;
  assign nand_199_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23563" *) _02758_;
  assign _05244_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23567" *) _03994_;
  assign _05245_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *) _08618_;
  assign _05246_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *) _02761_;
  assign nor_2406_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *) _08619_;
  assign _05247_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23576" *) _03995_;
  assign _05248_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *) _08622_;
  assign _05249_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *) _02764_;
  assign nor_2401_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *) _08623_;
  assign _05250_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23585" *) _03996_;
  assign _05251_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *) _08627_;
  assign _05252_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *) _02766_;
  assign nor_2396_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *) _08628_;
  assign _05253_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23595" *) mux_tmp_1227;
  assign nor_1351_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23595" *) _08629_;
  assign _05254_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23599" *) and_283_cse;
  assign nor_1338_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23599" *) _08630_;
  assign nor_2251_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23602" *) _08631_;
  assign nor_2252_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23606" *) _08632_;
  assign _00061_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23608" *) mux_tmp_1419;
  assign _00062_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23615" *) mux_1426_nl;
  assign _05255_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23620" *) _02767_;
  assign nor_2113_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23620" *) _08633_;
  assign _05256_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23622" *) mux_tmp_1469;
  assign nor_1303_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23622" *) _08634_;
  assign _05257_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23625" *) _02768_;
  assign nor_1302_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23625" *) _08635_;
  assign _00235_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23633" *) chn_in_rsci_d_mxwt[23];
  assign nor_1263_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23636" *) _08636_;
  assign nor_1264_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23642" *) _08642_;
  assign nor_1261_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23647" *) _08648_;
  assign _05258_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23650" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2;
  assign _05259_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23651" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2;
  assign nor_1262_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23653" *) _08653_;
  assign _00236_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23656" *) chn_in_rsci_d_mxwt[55];
  assign nor_1259_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23659" *) _08654_;
  assign nor_1260_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23665" *) _08660_;
  assign nor_1257_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23670" *) _08666_;
  assign _05260_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23673" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _05261_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23674" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign nor_1258_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23676" *) _08671_;
  assign _00237_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23679" *) chn_in_rsci_d_mxwt[87];
  assign nor_1255_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23682" *) _08672_;
  assign nor_1256_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23688" *) _08678_;
  assign nor_1253_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23693" *) _08684_;
  assign _05262_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23696" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _05263_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23697" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign nor_1254_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23699" *) _08689_;
  assign _00238_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23702" *) chn_in_rsci_d_mxwt[119];
  assign nor_1251_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23705" *) _08690_;
  assign nor_1252_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23711" *) _08696_;
  assign nor_1249_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23716" *) _08702_;
  assign _05264_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23719" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _05265_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23720" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign nor_1250_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23722" *) _08707_;
  assign _00239_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23725" *) chn_in_rsci_d_mxwt[151];
  assign _05266_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23726" *) or_tmp_2466;
  assign nor_1247_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23728" *) _08712_;
  assign nor_1099_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23729" *) or_tmp_2469;
  assign nor_1248_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23734" *) _08719_;
  assign _05267_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *) _02778_;
  assign nor_1245_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *) _08720_;
  assign _05268_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23742" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _05269_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23743" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign nor_1246_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23745" *) _08724_;
  assign _00240_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23748" *) chn_in_rsci_d_mxwt[183];
  assign nor_1243_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23751" *) _08727_;
  assign nor_1244_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23757" *) _08733_;
  assign nor_1241_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23762" *) _08739_;
  assign _05270_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23765" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _05271_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23766" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign nor_1242_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23768" *) _08744_;
  assign _00241_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23771" *) chn_in_rsci_d_mxwt[215];
  assign nor_1239_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23774" *) _08747_;
  assign nor_1240_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23780" *) _08753_;
  assign nor_1237_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23785" *) _08759_;
  assign _05272_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23788" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _05273_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23789" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign nor_1238_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23791" *) _08764_;
  assign _00242_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23794" *) chn_in_rsci_d_mxwt[247];
  assign nor_1235_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23797" *) _08765_;
  assign nor_1236_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23803" *) _08771_;
  assign nor_1233_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23808" *) _08777_;
  assign _05274_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23811" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _05275_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23812" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign nor_1234_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23814" *) _08782_;
  assign _00243_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23817" *) chn_in_rsci_d_mxwt[279];
  assign nor_1231_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23820" *) _08783_;
  assign nor_1232_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23826" *) _08789_;
  assign nor_1229_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23831" *) _08795_;
  assign _05276_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23834" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _05277_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23835" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign nor_1230_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23837" *) _08800_;
  assign _00244_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23840" *) chn_in_rsci_d_mxwt[311];
  assign nor_1227_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23843" *) _08803_;
  assign nor_1228_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23849" *) _08809_;
  assign nor_1225_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23854" *) _08815_;
  assign _05278_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23857" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _05279_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23858" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign nor_1226_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23860" *) _08820_;
  assign _00245_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23863" *) chn_in_rsci_d_mxwt[343];
  assign nor_1223_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23866" *) _08821_;
  assign nor_1224_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23872" *) _08827_;
  assign nor_1221_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23877" *) _08833_;
  assign _05280_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23880" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _05281_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23881" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign nor_1222_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23883" *) _08838_;
  assign _00246_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23886" *) chn_in_rsci_d_mxwt[375];
  assign nor_1219_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23889" *) _08839_;
  assign nor_1220_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23895" *) _08845_;
  assign nor_1217_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23900" *) _08851_;
  assign _05282_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23903" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _05283_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23904" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign nor_1218_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23906" *) _08856_;
  assign _00247_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23909" *) chn_in_rsci_d_mxwt[407];
  assign nor_1215_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23912" *) _08859_;
  assign nor_1216_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23918" *) _08865_;
  assign nor_1213_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23923" *) _08871_;
  assign _05284_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23926" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _05285_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23927" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign nor_1214_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23929" *) _08876_;
  assign _00248_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23932" *) chn_in_rsci_d_mxwt[439];
  assign nor_1211_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23935" *) _08877_;
  assign nor_1212_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23941" *) _08883_;
  assign nor_1209_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23946" *) _08889_;
  assign _05286_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23949" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _05287_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23950" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign nor_1210_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23952" *) _08894_;
  assign _00249_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23955" *) chn_in_rsci_d_mxwt[471];
  assign nor_1207_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23958" *) _08895_;
  assign nor_1208_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23964" *) _08901_;
  assign nor_1205_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23969" *) _08907_;
  assign _05288_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23972" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _05289_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23973" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign nor_1206_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23975" *) _08912_;
  assign _00250_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23978" *) chn_in_rsci_d_mxwt[503];
  assign nor_1203_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23981" *) _08913_;
  assign nor_1204_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23987" *) _08919_;
  assign nor_1201_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23992" *) _08925_;
  assign _05290_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23995" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2;
  assign _05291_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23996" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2;
  assign nor_1202_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23998" *) _08930_;
  assign _05292_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *) _02792_;
  assign nor_1200_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *) _08946_;
  assign _05293_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24063" *) _02795_;
  assign nor_1198_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24063" *) _08955_;
  assign IsNaN_5U_10U_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24092" *) _04169_;
  assign IsNaN_5U_10U_IsNaN_5U_10U_nand_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24099" *) _02796_;
  assign IsNaN_5U_10U_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24105" *) _04170_;
  assign IsNaN_5U_10U_IsNaN_5U_10U_nand_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24110" *) _02797_;
  assign IsNaN_5U_10U_nor_14_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24114" *) _04171_;
  assign IsNaN_5U_10U_IsNaN_5U_10U_nand_14_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24119" *) _02798_;
  assign _05294_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24123" *) mux_tmp_129;
  assign _05295_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24125" *) and_tmp_18;
  assign _05296_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24127" *) mux_tmp_151;
  assign _05297_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24132" *) _02799_;
  assign _00067_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24221" *) mux_1437_cse;
  assign _05298_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24229" *) _02800_;
  assign nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6907" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6913" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6919" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6925" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6931" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6937" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6943" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6949" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6955" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6961" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6967" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6973" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6979" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6985" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6991" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:6997" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1[0];
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7122" *) chn_idata_data_sva_1_27_0_1[23];
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7131" *) chn_idata_data_sva_1_59_31_1[24];
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7140" *) chn_idata_data_sva_1_91_63_1[24];
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7149" *) chn_idata_data_sva_1_123_95_1[24];
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7158" *) chn_idata_data_sva_1_155_127_1[24];
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7167" *) chn_idata_data_sva_1_187_159_1[24];
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7176" *) chn_idata_data_sva_1_219_191_1[24];
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7185" *) chn_idata_data_sva_1_251_223_1[24];
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7194" *) chn_idata_data_sva_1_283_255_1[24];
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7203" *) chn_idata_data_sva_1_315_287_1[24];
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7212" *) chn_idata_data_sva_1_347_319_1[24];
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7221" *) chn_idata_data_sva_1_379_351_1[24];
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7230" *) chn_idata_data_sva_1_411_383_1[24];
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7239" *) chn_idata_data_sva_1_443_415_1[24];
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7248" *) chn_idata_data_sva_1_475_447_1[24];
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7257" *) chn_idata_data_sva_1_507_479_1[24];
  assign _05299_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8774" *) or_dcpl_4;
  assign _05300_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8799" *) mux_2355_nl;
  assign _05301_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8821" *) IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  assign nand_219_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8822" *) _03632_;
  assign nor_2047_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8824" *) or_306_cse;
  assign _05302_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8825" *) IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  assign nor_2046_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8827" *) or_tmp_378;
  assign _05303_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8830" *) IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  assign _05304_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8831" *) IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  assign _05305_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8841" *) IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  assign _05306_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8845" *) mux_169_nl;
  assign _05307_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8846" *) IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  assign _05308_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8847" *) IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  assign _05309_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8848" *) IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  assign nor_45_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8849" *) or_309_cse;
  assign _05310_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8853" *) IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  assign _05311_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8854" *) IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  assign _05312_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8855" *) IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  assign _05313_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8856" *) IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  assign _05314_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8857" *) IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  assign _05315_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8858" *) IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  assign _05316_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8859" *) IsNaN_8U_23U_land_lpi_1_dfm_3;
  assign _05317_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8861" *) mux_tmp_200;
  assign nor_2026_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8861" *) _09460_;
  assign nor_57_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8874" *) or_1198_cse;
  assign nor_2011_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8879" *) _09462_;
  assign nor_63_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8885" *) or_578_cse;
  assign nor_2004_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8886" *) or_243_nl;
  assign nor_2005_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8888" *) _09464_;
  assign nor_1980_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8897" *) _09466_;
  assign _00068_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8902" *) mux_tmp_321;
  assign nor_2150_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8911" *) or_183_cse_1;
  assign nor_1314_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8913" *) or_tmp_3763;
  assign nor_2326_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8913" *) _09468_;
  assign nor_1958_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8932" *) _09470_;
  assign _05321_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8947" *) _09471_;
  assign _05322_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8954" *) mux_tmp_345;
  assign nor_1939_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8954" *) _09472_;
  assign nor_1917_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8964" *) _09473_;
  assign _05323_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8966" *) mux_tmp_435;
  assign nor_1898_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8966" *) _09474_;
  assign _05325_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8979" *) mux_tmp_317;
  assign nor_1875_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8979" *) _09476_;
  assign _05326_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9007" *) or_tmp_3379;
  assign nor_2300_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9007" *) _09477_;
  assign _05327_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9011" *) _09478_;
  assign _05328_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9016" *) or_tmp_3025;
  assign nand_51_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9016" *) _03664_;
  assign nor_1772_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9025" *) _09479_;
  assign nand_225_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9032" *) _03666_;
  assign _05329_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9045" *) mux_1463_cse;
  assign nor_1761_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9045" *) _09481_;
  assign _05330_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9051" *) _03671_;
  assign _00072_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9063" *) mux_tmp_1813;
  assign _05331_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9071" *) mux_tmp_766;
  assign nor_1683_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9071" *) _09483_;
  assign nor_1674_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9073" *) _09484_;
  assign nor_1056_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9082" *) _09487_;
  assign nor_1666_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9085" *) _08363_;
  assign nor_1669_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9087" *) _09489_;
  assign nor_1664_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9092" *) or_dcpl_147;
  assign nor_1659_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9096" *) _09494_;
  assign nor_1661_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9099" *) _09497_;
  assign nand_207_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9107" *) _03676_;
  assign nor_2099_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9110" *) or_4709_cse;
  assign _05332_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9120" *) chn_idata_data_sva_2_79_63_1[0];
  assign nor_2100_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9131" *) _08368_;
  assign nor_2101_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9133" *) _09500_;
  assign nor_2285_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9142" *) or_300_cse;
  assign nor_2219_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9144" *) or_4714_cse;
  assign _05334_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9151" *) chn_idata_data_sva_2_111_95_1[0];
  assign _05335_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9156" *) IsNaN_5U_10U_land_3_lpi_1_dfm_4;
  assign _05336_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9167" *) _03685_;
  assign nor_2284_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9167" *) _09501_;
  assign _05337_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9169" *) _09502_;
  assign nor_1049_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9176" *) _09508_;
  assign nor_1048_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9178" *) _09509_;
  assign _05338_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9183" *) chn_idata_data_sva_2_511_1;
  assign _05339_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9188" *) IsNaN_5U_10U_land_lpi_1_dfm_4;
  assign _05340_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9217" *) IsNaN_5U_10U_land_5_lpi_1_dfm_4;
  assign nor_1624_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9228" *) _09515_;
  assign nor_1630_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9229" *) _09517_;
  assign nor_1629_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9230" *) or_1157_cse;
  assign nor_1626_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9231" *) _09519_;
  assign nor_1040_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9234" *) _09521_;
  assign _05342_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9264" *) or_4749_cse;
  assign nor_1033_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9271" *) _09527_;
  assign _05343_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9276" *) chn_idata_data_sva_2_207_191_1[0];
  assign _05344_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9281" *) IsNaN_5U_10U_land_6_lpi_1_dfm_4;
  assign _05345_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *) _09528_;
  assign _05346_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *) _03709_;
  assign _05347_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *) _09529_;
  assign _05348_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9301" *) chn_idata_data_sva_2_463_447_1[0];
  assign _05349_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9306" *) IsNaN_5U_10U_land_14_lpi_1_dfm_5;
  assign nor_2142_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9310" *) _09532_;
  assign nor_2143_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9312" *) _09533_;
  assign nor_183_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9325" *) or_3542_cse;
  assign _05350_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9333" *) IsNaN_5U_10U_land_7_lpi_1_dfm_5;
  assign nor_1589_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9342" *) or_5254_cse;
  assign _05351_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9345" *) chn_idata_data_sva_2_431_415_1[0];
  assign _05352_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9350" *) IsNaN_5U_10U_land_13_lpi_1_dfm_4;
  assign nor_2269_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9364" *) _09535_;
  assign _05353_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9367" *) _03728_;
  assign _05354_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9381" *) IsNaN_5U_10U_land_8_lpi_1_dfm_4;
  assign _05355_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9394" *) chn_idata_data_sva_2_399_383_1[0];
  assign _05356_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9399" *) IsNaN_5U_10U_land_12_lpi_1_dfm_4;
  assign _05357_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9423" *) chn_idata_data_sva_2_303_287_1[0];
  assign _05358_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9428" *) IsNaN_5U_10U_land_9_lpi_1_dfm_4;
  assign _05359_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9443" *) chn_idata_data_sva_2_367_351_1[0];
  assign _05360_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9448" *) IsNaN_5U_10U_land_11_lpi_1_dfm_4;
  assign _05361_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9460" *) chn_idata_data_sva_2_335_319_1[0];
  assign _05362_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9465" *) IsNaN_5U_10U_land_10_lpi_1_dfm_4;
  assign nor_1556_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9477" *) or_1483_nl;
  assign _05363_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9479" *) fsm_output[0];
  assign _05364_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9481" *) _09537_;
  assign _05365_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9482" *) mux_948_nl;
  assign reg_cvt_else_cvt_else_nor_4_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9484" *) _09538_;
  assign _00073_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9487" *) or_5379_cse;
  assign nor_1536_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9489" *) _09539_;
  assign _05366_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *) _09541_;
  assign _05367_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *) mux_991_nl;
  assign _05368_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9495" *) _09542_;
  assign nor_1523_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9497" *) _09544_;
  assign nor_1524_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9499" *) _08497_;
  assign nor_1525_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9501" *) _09547_;
  assign _00001_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9508" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16;
  assign _00002_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9519" *) mux_1966_itm;
  assign _00003_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9529" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17;
  assign _05369_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9533" *) cvt_2_FpMantRNE_17U_11U_else_and_1_tmp;
  assign nor_1500_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *) _09554_;
  assign nor_1498_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9544" *) _09558_;
  assign _00004_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9550" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18;
  assign _05370_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9554" *) cvt_3_FpMantRNE_17U_11U_else_and_1_tmp;
  assign nor_1488_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9562" *) _09559_;
  assign nor_1489_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9564" *) _09560_;
  assign _00005_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9577" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19;
  assign _05371_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9581" *) cvt_4_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _00006_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9591" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20;
  assign _05372_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9595" *) cvt_5_FpMantRNE_17U_11U_else_and_1_tmp;
  assign _05373_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9606" *) mux_tmp_960;
  assign nor_1463_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9606" *) _09562_;
  assign _00007_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9610" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21;
  assign _00008_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9623" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22;
  assign _05374_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9627" *) cvt_7_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _00009_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9636" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23;
  assign _05375_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9640" *) cvt_8_FpMantRNE_17U_11U_else_and_3_tmp;
  assign nor_1434_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9647" *) _09563_;
  assign _00010_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9652" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24;
  assign _05376_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9656" *) cvt_9_FpMantRNE_17U_11U_else_and_1_tmp;
  assign _00011_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9668" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25;
  assign _05377_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9672" *) cvt_10_FpMantRNE_17U_11U_else_and_2_tmp;
  assign nor_1415_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9679" *) _09564_;
  assign _00012_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9684" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26;
  assign _05378_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9688" *) cvt_11_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _00013_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9700" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27;
  assign _05379_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9704" *) cvt_12_FpMantRNE_17U_11U_else_and_3_tmp;
  assign _00014_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9717" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28;
  assign _05380_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9721" *) cvt_13_FpMantRNE_17U_11U_else_and_2_tmp;
  assign _00015_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9731" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29;
  assign _05381_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9735" *) cvt_14_FpMantRNE_17U_11U_else_and_3_tmp;
  assign _00016_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9751" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30;
  assign _00017_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9765" *) libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31;
  assign _05382_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9769" *) cvt_16_FpMantRNE_17U_11U_else_and_4_tmp;
  assign _00000_[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9826" *) mux_2020_nl;
  assign _00000_[1] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9826" *) mux_2015_nl;
  assign _00074_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9835" *) mux_1343_nl;
  assign _05384_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9838" *) mux_1345_nl;
  assign nand_190_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9840" *) _03818_;
  assign _05385_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9850" *) mux_1442_nl;
  assign nor_1309_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9852" *) _09568_;
  assign nor_1310_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9854" *) _09569_;
  assign nor_1306_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9858" *) _09570_;
  assign _05386_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9861" *) _03819_;
  assign nor_2130_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9861" *) _09571_;
  assign _05387_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9864" *) mux_1466_cse;
  assign nor_1305_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9864" *) _09572_;
  assign _05388_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9869" *) _03820_;
  assign nor_2114_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9869" *) _09573_;
  assign nor_1301_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9875" *) _09574_;
  assign _05389_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9879" *) _03821_;
  assign nor_2127_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9879" *) _09575_;
  assign nor_1287_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9881" *) _09576_;
  assign _05390_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9884" *) _03822_;
  assign nor_2110_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9884" *) _09577_;
  assign nand_171_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9889" *) and_2487_nl;
  assign nor_1271_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9891" *) _09579_;
  assign _05391_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9899" *) mux_124_nl;
  assign _05392_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9901" *) or_dcpl_32;
  assign _05393_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9902" *) mux_130_nl;
  assign _05394_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9905" *) mux_133_cse;
  assign _05395_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9910" *) mux_118_nl;
  assign _05396_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9913" *) mux_149_nl;
  assign _05397_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9916" *) mux_152_nl;
  assign nand_164_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9918" *) _03824_;
  assign nand_162_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9920" *) _03825_;
  assign nand_160_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9922" *) _03826_;
  assign nand_158_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9924" *) _03827_;
  assign nand_156_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9926" *) _03828_;
  assign nand_153_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9928" *) _03829_;
  assign nand_151_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9930" *) _03830_;
  assign nand_149_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9932" *) _03831_;
  assign nand_147_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9934" *) _03832_;
  assign nand_145_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9936" *) _03833_;
  assign nand_143_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9938" *) _03834_;
  assign nand_141_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9940" *) _03835_;
  assign nand_139_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9942" *) _03836_;
  assign nand_137_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9944" *) _03837_;
  assign nand_135_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9946" *) _03838_;
  assign nand_133_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9948" *) _03839_;
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9966" *) _09581_;
  assign _05398_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9968" *) cvt_16_IntSaturation_17U_16U_if_acc_4_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9972" *) _09583_;
  assign _05399_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9974" *) cvt_15_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9978" *) _09585_;
  assign _05400_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9980" *) cvt_14_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9984" *) _09587_;
  assign _05401_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9986" *) cvt_13_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9990" *) _09589_;
  assign _05402_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9992" *) cvt_12_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9996" *) _09591_;
  assign _05403_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9998" *) cvt_11_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _05404_ = cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10002" *) cvt_10_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _05405_ = _05404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10002" *) and_dcpl_93;
  assign _05406_ = cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10008" *) cvt_9_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _05407_ = _05406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10008" *) and_dcpl_93;
  assign _05408_ = cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10014" *) cvt_8_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _05409_ = _05408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10014" *) and_dcpl_93;
  assign _05410_ = cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10020" *) cvt_7_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _05411_ = _05410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10020" *) and_dcpl_93;
  assign _05412_ = cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10026" *) cvt_6_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _05413_ = _05412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10026" *) and_dcpl_93;
  assign _05414_ = cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10032" *) cvt_5_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _05415_ = _05414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10032" *) and_dcpl_93;
  assign _05416_ = cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10038" *) cvt_4_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _05417_ = _05416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10038" *) and_dcpl_93;
  assign _05418_ = cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10044" *) cvt_3_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _05419_ = _05418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10044" *) and_dcpl_93;
  assign _05420_ = cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10050" *) cvt_2_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _05421_ = _05420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10050" *) and_dcpl_93;
  assign _05422_ = cvt_1_IntSaturation_17U_16U_else_if_acc_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10056" *) cvt_1_IntSaturation_17U_16U_if_acc_nl[2];
  assign _05423_ = _05422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10056" *) and_dcpl_93;
  assign _05424_ = _04185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *) _04186_;
  assign _05425_ = _05424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10061" *) cfg_mode_eql_1_sva_4;
  assign _05426_ = _04006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10064" *) _04185_;
  assign _05427_ = or_309_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10065" *) _00058_;
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse = _01445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10071" *) and_1385_rgt;
  assign or_479_nl = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10072" *) _00064_;
  assign or_547_nl = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10076" *) _04187_;
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse = _01448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10080" *) and_1385_rgt;
  assign or_626_nl = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10081" *) _04188_;
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_15_cse = _01453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10087" *) and_1385_rgt;
  assign _05428_ = _01455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10091" *) and_1385_rgt;
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_8_cse = _01458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10094" *) and_1385_rgt;
  assign or_5379_cse = _00065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10095" *) main_stage_v_1;
  assign or_186_cse = or_183_cse_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10097" *) and_dcpl_3;
  assign or_dcpl_16 = or_dcpl_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10106" *) _04185_;
  assign _05429_ = or_dcpl_16 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10106" *) or_2251_nl;
  assign or_217_nl = or_2251_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10107" *) _04187_;
  assign or_226_nl = or_2251_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10111" *) _04188_;
  assign or_dcpl_32 = or_dcpl_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10115" *) or_dcpl_30;
  assign _05430_ = or_dcpl_32 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10115" *) or_2251_nl;
  assign or_243_nl = or_2251_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10116" *) _00064_;
  assign _05431_ = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10809" *) cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp;
  assign _00187_[2] = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_4_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10811" *) cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp;
  assign _05432_ = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10817" *) cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp;
  assign _00203_[0] = _04222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10817" *) cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp;
  assign _05433_ = IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10819" *) _04007_;
  assign _05434_ = _05433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10819" *) IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0;
  assign _05435_ = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10821" *) cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign _00188_[2] = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10823" *) cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _05436_ = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10829" *) cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _00204_[0] = _04223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10829" *) cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign _05437_ = IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10831" *) _04008_;
  assign _05438_ = _05437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10831" *) IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0;
  assign _05439_ = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10836" *) cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign _00189_[2] = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10838" *) cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _05440_ = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10844" *) cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _00205_[0] = _04224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10844" *) cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign _05441_ = IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10846" *) _04009_;
  assign _05442_ = _05441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10846" *) IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0;
  assign or_dcpl_108 = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10848" *) cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_109 = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10850" *) cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _05443_ = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10856" *) cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _00206_[0] = _04225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10856" *) cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_110 = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10864" *) cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign or_dcpl_111 = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10866" *) cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _05444_ = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10872" *) cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _00207_[0] = _04226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10872" *) cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign _05445_ = IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10874" *) _04010_;
  assign _05446_ = _05445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10874" *) IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0;
  assign or_dcpl_113 = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10876" *) cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_114 = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10878" *) cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _05447_ = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10884" *) cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _00208_[0] = _04227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10884" *) cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_115 = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10889" *) cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_116 = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10891" *) cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _05448_ = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10897" *) cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _00209_[0] = _04228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10897" *) cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_119 = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10899" *) cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign or_dcpl_120 = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10901" *) cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _05449_ = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10907" *) cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _00210_[0] = _04229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10907" *) cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign _05450_ = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10918" *) cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign _00195_[2] = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10920" *) cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _05451_ = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10926" *) cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign _00211_[0] = _04230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10926" *) cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign _05452_ = IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10928" *) _04011_;
  assign _05453_ = _05452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10928" *) IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0;
  assign or_dcpl_124 = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10930" *) cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_125 = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10932" *) cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _05454_ = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10938" *) cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _00212_[0] = _04231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10938" *) cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_126 = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10940" *) cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_127 = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10942" *) cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _05455_ = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10948" *) cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _00213_[0] = _04232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10948" *) cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_130 = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10950" *) cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign or_dcpl_131 = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10952" *) cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _05456_ = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10958" *) cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _00214_[0] = _04233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10958" *) cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign or_dcpl_132 = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10960" *) cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_133 = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10962" *) cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _05457_ = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10968" *) cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign _00215_[0] = _04234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10968" *) cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_136 = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10970" *) cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign or_dcpl_137 = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10972" *) cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _05458_ = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10978" *) cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _00216_[0] = _04235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10978" *) cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign or_dcpl_139 = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10980" *) cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign or_dcpl_140 = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10982" *) cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _05459_ = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10988" *) cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign _00217_[0] = _04236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10988" *) cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  assign or_dcpl_143 = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10990" *) cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp;
  assign or_dcpl_144 = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_24_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10992" *) cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp;
  assign _05460_ = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10998" *) cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp;
  assign _00218_[0] = _04237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:10998" *) cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp;
  assign _05461_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11006" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva;
  assign _04519_ = _04238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11006" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva;
  assign _05462_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11008" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva;
  assign cvt_1_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_nl = _04239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11009" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva;
  assign _05383_ = IsNaN_5U_10U_nor_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11014" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2;
  assign _05463_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11016" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva;
  assign _04521_ = _04241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11016" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva;
  assign _05464_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11018" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva;
  assign cvt_2_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl = _04242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11019" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva;
  assign _05333_ = IsNaN_5U_10U_nor_1_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11024" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  assign _05465_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11026" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva;
  assign _04523_ = _04244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11026" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva;
  assign _05466_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11032" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva;
  assign cvt_3_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl = _04245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11033" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva;
  assign _05467_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11039" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva;
  assign _04525_ = _04247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11039" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva;
  assign _05468_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11041" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva;
  assign cvt_4_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl = _04248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11042" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva;
  assign _05469_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11048" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva;
  assign _04527_ = _04250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11048" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva;
  assign _05470_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11054" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva;
  assign cvt_5_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl = _04251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11055" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva;
  assign _05471_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11061" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva;
  assign _04549_ = _04253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11061" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva;
  assign _05472_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11063" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva;
  assign cvt_16_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_4_nl = _04254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11064" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva;
  assign _05473_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11070" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva;
  assign _04529_ = _04256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11070" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva;
  assign _05474_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11072" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva;
  assign cvt_6_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl = _04257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11073" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva;
  assign _05475_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11079" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva;
  assign _04547_ = _04259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11079" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva;
  assign _05476_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11085" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva;
  assign cvt_15_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl = _04260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11086" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva;
  assign _05341_ = IsNaN_5U_10U_nor_14_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11091" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2;
  assign _05477_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11093" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva;
  assign _04531_ = _04262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11093" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva;
  assign _05478_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11095" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva;
  assign cvt_7_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl = _04263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11096" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva;
  assign _05479_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11102" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva;
  assign _04545_ = _04265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11102" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva;
  assign _05480_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11104" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva;
  assign cvt_14_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl = _04266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11105" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva;
  assign _05481_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11111" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva;
  assign _04533_ = _04268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11111" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva;
  assign _05482_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11113" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva;
  assign cvt_8_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl = _04269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11114" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva;
  assign _05483_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11120" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva;
  assign _04543_ = _04271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11120" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva;
  assign _05484_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11122" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva;
  assign cvt_13_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl = _04272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11123" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva;
  assign _05485_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11129" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva;
  assign _04535_ = _04274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11129" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva;
  assign _05486_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11135" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva;
  assign cvt_9_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl = _04275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11136" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva;
  assign _05487_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11142" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva;
  assign _04541_ = _04277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11142" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva;
  assign _05488_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11144" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva;
  assign cvt_12_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl = _04278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11145" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva;
  assign _05489_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11151" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva;
  assign _04537_ = _04280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11151" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva;
  assign _05490_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11153" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva;
  assign cvt_10_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl = _04281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11154" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva;
  assign _05491_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11160" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva;
  assign _04539_ = _04283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11160" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva;
  assign _05492_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[25] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11162" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva;
  assign cvt_11_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl = _04284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11163" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_13_nl = _01462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11235" *) cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1;
  assign or_3872_nl = and_dcpl_954 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11255" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign _05493_ = _01464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11262" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign or_3891_nl = and_dcpl_962 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11275" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign _05494_ = _01466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11282" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign or_3900_nl = and_dcpl_966 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11289" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign _05495_ = _01468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11296" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign or_3911_nl = and_dcpl_970 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11303" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign _05496_ = _01470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11310" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign or_3932_nl = and_dcpl_978 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11317" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign _05497_ = _01472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11324" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign or_3942_nl = and_dcpl_982 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11331" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign _05498_ = _01474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11338" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign or_3953_nl = and_dcpl_987 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11345" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign _05499_ = _01476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11352" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign or_3965_nl = and_dcpl_991 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11359" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign _05500_ = _01478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11366" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign or_3977_nl = and_dcpl_995 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11373" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign _05501_ = _01480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11380" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign or_3989_nl = and_dcpl_999 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11387" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign _05502_ = _01482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11394" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign or_3999_nl = and_dcpl_1003 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11401" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign _05503_ = _01484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11408" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2;
  assign _05504_ = IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11410" *) _04012_;
  assign _05505_ = _05504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11410" *) IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0;
  assign _05506_ = IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11412" *) _04013_;
  assign _05507_ = _05506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11413" *) IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0;
  assign _05508_ = IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11415" *) _04014_;
  assign _05509_ = _05508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11416" *) IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0;
  assign _05510_ = IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11418" *) _04015_;
  assign _05511_ = _05510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11419" *) IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0;
  assign _05512_ = IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11421" *) _04016_;
  assign _05513_ = _05512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11421" *) IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0;
  assign _05514_ = IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11423" *) _04017_;
  assign _05515_ = _05514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11423" *) IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0;
  assign _05516_ = IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11425" *) _04018_;
  assign _05517_ = _05516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11425" *) IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0;
  assign _05518_ = IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11427" *) _04019_;
  assign _05519_ = _05518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11427" *) IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0;
  assign _05520_ = IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11429" *) _04020_;
  assign _05521_ = _05520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11430" *) IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0;
  assign _05522_ = IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11432" *) _04021_;
  assign _05523_ = _05522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11433" *) IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0;
  assign _05524_ = IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11435" *) _04022_;
  assign _05525_ = _05524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11436" *) IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0;
  assign _05526_ = chn_in_rsci_d_mxwt[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11438" *) chn_in_rsci_d_mxwt[1];
  assign _05527_ = _05526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11438" *) chn_in_rsci_d_mxwt[2];
  assign _05528_ = _05527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11439" *) chn_in_rsci_d_mxwt[3];
  assign _05529_ = _05528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11439" *) chn_in_rsci_d_mxwt[4];
  assign _05530_ = _05529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11439" *) chn_in_rsci_d_mxwt[5];
  assign _05531_ = _05530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11440" *) chn_in_rsci_d_mxwt[6];
  assign _05532_ = _05531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11440" *) chn_in_rsci_d_mxwt[7];
  assign _05533_ = _05532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11440" *) chn_in_rsci_d_mxwt[8];
  assign _05534_ = _05533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *) chn_in_rsci_d_mxwt[9];
  assign _05535_ = _05534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *) chn_in_rsci_d_mxwt[10];
  assign _05536_ = _05535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *) chn_in_rsci_d_mxwt[11];
  assign _05537_ = _05536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11441" *) chn_in_rsci_d_mxwt[13];
  assign _05538_ = chn_in_rsci_d_mxwt[32] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11443" *) chn_in_rsci_d_mxwt[33];
  assign _05539_ = _05538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11443" *) chn_in_rsci_d_mxwt[34];
  assign _05540_ = _05539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11444" *) chn_in_rsci_d_mxwt[35];
  assign _05541_ = _05540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11444" *) chn_in_rsci_d_mxwt[36];
  assign _05542_ = _05541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11444" *) chn_in_rsci_d_mxwt[37];
  assign _05543_ = _05542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11445" *) chn_in_rsci_d_mxwt[38];
  assign _05544_ = _05543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11445" *) chn_in_rsci_d_mxwt[39];
  assign _05545_ = _05544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11445" *) chn_in_rsci_d_mxwt[40];
  assign _05546_ = _05545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *) chn_in_rsci_d_mxwt[41];
  assign _05547_ = _05546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *) chn_in_rsci_d_mxwt[42];
  assign _05548_ = _05547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *) chn_in_rsci_d_mxwt[43];
  assign _05549_ = _05548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11446" *) chn_in_rsci_d_mxwt[45];
  assign _05550_ = chn_in_rsci_d_mxwt[64] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11448" *) chn_in_rsci_d_mxwt[65];
  assign _05551_ = _05550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11448" *) chn_in_rsci_d_mxwt[66];
  assign _05552_ = _05551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11449" *) chn_in_rsci_d_mxwt[67];
  assign _05553_ = _05552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11449" *) chn_in_rsci_d_mxwt[68];
  assign _05554_ = _05553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11449" *) chn_in_rsci_d_mxwt[69];
  assign _05555_ = _05554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11450" *) chn_in_rsci_d_mxwt[70];
  assign _05556_ = _05555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11450" *) chn_in_rsci_d_mxwt[71];
  assign _05557_ = _05556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11450" *) chn_in_rsci_d_mxwt[72];
  assign _05558_ = _05557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *) chn_in_rsci_d_mxwt[73];
  assign _05559_ = _05558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *) chn_in_rsci_d_mxwt[74];
  assign _05560_ = _05559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *) chn_in_rsci_d_mxwt[75];
  assign _05561_ = _05560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11451" *) chn_in_rsci_d_mxwt[77];
  assign _05562_ = chn_in_rsci_d_mxwt[96] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11453" *) chn_in_rsci_d_mxwt[97];
  assign _05563_ = _05562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11453" *) chn_in_rsci_d_mxwt[98];
  assign _05564_ = _05563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11454" *) chn_in_rsci_d_mxwt[99];
  assign _05565_ = _05564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11454" *) chn_in_rsci_d_mxwt[100];
  assign _05566_ = _05565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11454" *) chn_in_rsci_d_mxwt[101];
  assign _05567_ = _05566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11455" *) chn_in_rsci_d_mxwt[102];
  assign _05568_ = _05567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11455" *) chn_in_rsci_d_mxwt[103];
  assign _05569_ = _05568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11455" *) chn_in_rsci_d_mxwt[104];
  assign _05570_ = _05569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *) chn_in_rsci_d_mxwt[105];
  assign _05571_ = _05570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *) chn_in_rsci_d_mxwt[106];
  assign _05572_ = _05571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *) chn_in_rsci_d_mxwt[107];
  assign _05573_ = _05572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11456" *) chn_in_rsci_d_mxwt[109];
  assign _05574_ = chn_in_rsci_d_mxwt[128] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11458" *) chn_in_rsci_d_mxwt[129];
  assign _05575_ = _05574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11458" *) chn_in_rsci_d_mxwt[130];
  assign _05576_ = _05575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11459" *) chn_in_rsci_d_mxwt[131];
  assign _05577_ = _05576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11459" *) chn_in_rsci_d_mxwt[132];
  assign _05578_ = _05577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11459" *) chn_in_rsci_d_mxwt[133];
  assign _05579_ = _05578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11460" *) chn_in_rsci_d_mxwt[134];
  assign _05580_ = _05579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11460" *) chn_in_rsci_d_mxwt[135];
  assign _05581_ = _05580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11460" *) chn_in_rsci_d_mxwt[136];
  assign _05582_ = _05581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *) chn_in_rsci_d_mxwt[137];
  assign _05583_ = _05582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *) chn_in_rsci_d_mxwt[138];
  assign _05584_ = _05583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *) chn_in_rsci_d_mxwt[139];
  assign _05585_ = _05584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11461" *) chn_in_rsci_d_mxwt[141];
  assign _05586_ = chn_in_rsci_d_mxwt[160] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11463" *) chn_in_rsci_d_mxwt[161];
  assign _05587_ = _05586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11463" *) chn_in_rsci_d_mxwt[162];
  assign _05588_ = _05587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11464" *) chn_in_rsci_d_mxwt[163];
  assign _05589_ = _05588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11464" *) chn_in_rsci_d_mxwt[164];
  assign _05590_ = _05589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11464" *) chn_in_rsci_d_mxwt[165];
  assign _05591_ = _05590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11465" *) chn_in_rsci_d_mxwt[166];
  assign _05592_ = _05591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11465" *) chn_in_rsci_d_mxwt[167];
  assign _05593_ = _05592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11465" *) chn_in_rsci_d_mxwt[168];
  assign _05594_ = _05593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *) chn_in_rsci_d_mxwt[169];
  assign _05595_ = _05594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *) chn_in_rsci_d_mxwt[170];
  assign _05596_ = _05595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *) chn_in_rsci_d_mxwt[171];
  assign _05597_ = _05596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11466" *) chn_in_rsci_d_mxwt[173];
  assign _05598_ = chn_in_rsci_d_mxwt[192] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11468" *) chn_in_rsci_d_mxwt[193];
  assign _05599_ = _05598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11468" *) chn_in_rsci_d_mxwt[194];
  assign _05600_ = _05599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11469" *) chn_in_rsci_d_mxwt[195];
  assign _05601_ = _05600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11469" *) chn_in_rsci_d_mxwt[196];
  assign _05602_ = _05601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11469" *) chn_in_rsci_d_mxwt[197];
  assign _05603_ = _05602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11470" *) chn_in_rsci_d_mxwt[198];
  assign _05604_ = _05603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11470" *) chn_in_rsci_d_mxwt[199];
  assign _05605_ = _05604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11470" *) chn_in_rsci_d_mxwt[200];
  assign _05606_ = _05605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *) chn_in_rsci_d_mxwt[201];
  assign _05607_ = _05606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *) chn_in_rsci_d_mxwt[202];
  assign _05608_ = _05607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *) chn_in_rsci_d_mxwt[203];
  assign _05609_ = _05608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11471" *) chn_in_rsci_d_mxwt[205];
  assign _05610_ = chn_in_rsci_d_mxwt[224] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11473" *) chn_in_rsci_d_mxwt[225];
  assign _05611_ = _05610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11473" *) chn_in_rsci_d_mxwt[226];
  assign _05612_ = _05611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11474" *) chn_in_rsci_d_mxwt[227];
  assign _05613_ = _05612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11474" *) chn_in_rsci_d_mxwt[228];
  assign _05614_ = _05613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11474" *) chn_in_rsci_d_mxwt[229];
  assign _05615_ = _05614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11475" *) chn_in_rsci_d_mxwt[230];
  assign _05616_ = _05615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11475" *) chn_in_rsci_d_mxwt[231];
  assign _05617_ = _05616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11475" *) chn_in_rsci_d_mxwt[232];
  assign _05618_ = _05617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *) chn_in_rsci_d_mxwt[233];
  assign _05619_ = _05618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *) chn_in_rsci_d_mxwt[234];
  assign _05620_ = _05619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *) chn_in_rsci_d_mxwt[235];
  assign _05621_ = _05620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11476" *) chn_in_rsci_d_mxwt[237];
  assign _05622_ = chn_in_rsci_d_mxwt[256] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11478" *) chn_in_rsci_d_mxwt[257];
  assign _05623_ = _05622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11478" *) chn_in_rsci_d_mxwt[258];
  assign _05624_ = _05623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11479" *) chn_in_rsci_d_mxwt[259];
  assign _05625_ = _05624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11479" *) chn_in_rsci_d_mxwt[260];
  assign _05626_ = _05625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11479" *) chn_in_rsci_d_mxwt[261];
  assign _05627_ = _05626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11480" *) chn_in_rsci_d_mxwt[262];
  assign _05628_ = _05627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11480" *) chn_in_rsci_d_mxwt[263];
  assign _05629_ = _05628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11480" *) chn_in_rsci_d_mxwt[264];
  assign _05630_ = _05629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *) chn_in_rsci_d_mxwt[265];
  assign _05631_ = _05630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *) chn_in_rsci_d_mxwt[266];
  assign _05632_ = _05631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *) chn_in_rsci_d_mxwt[267];
  assign _05633_ = _05632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11481" *) chn_in_rsci_d_mxwt[269];
  assign _05634_ = chn_in_rsci_d_mxwt[288] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11483" *) chn_in_rsci_d_mxwt[289];
  assign _05635_ = _05634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11484" *) chn_in_rsci_d_mxwt[290];
  assign _05636_ = _05635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11484" *) chn_in_rsci_d_mxwt[291];
  assign _05637_ = _05636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11484" *) chn_in_rsci_d_mxwt[292];
  assign _05638_ = _05637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11485" *) chn_in_rsci_d_mxwt[293];
  assign _05639_ = _05638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11485" *) chn_in_rsci_d_mxwt[294];
  assign _05640_ = _05639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11485" *) chn_in_rsci_d_mxwt[295];
  assign _05641_ = _05640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11486" *) chn_in_rsci_d_mxwt[296];
  assign _05642_ = _05641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11486" *) chn_in_rsci_d_mxwt[297];
  assign _05643_ = _05642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11486" *) chn_in_rsci_d_mxwt[298];
  assign _05644_ = _05643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11487" *) chn_in_rsci_d_mxwt[299];
  assign _05645_ = _05644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11487" *) chn_in_rsci_d_mxwt[301];
  assign _05646_ = chn_in_rsci_d_mxwt[320] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11489" *) chn_in_rsci_d_mxwt[321];
  assign _05647_ = _05646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11490" *) chn_in_rsci_d_mxwt[322];
  assign _05648_ = _05647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11490" *) chn_in_rsci_d_mxwt[323];
  assign _05649_ = _05648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11490" *) chn_in_rsci_d_mxwt[324];
  assign _05650_ = _05649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11491" *) chn_in_rsci_d_mxwt[325];
  assign _05651_ = _05650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11491" *) chn_in_rsci_d_mxwt[326];
  assign _05652_ = _05651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11491" *) chn_in_rsci_d_mxwt[327];
  assign _05653_ = _05652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11492" *) chn_in_rsci_d_mxwt[328];
  assign _05654_ = _05653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11492" *) chn_in_rsci_d_mxwt[329];
  assign _05655_ = _05654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11492" *) chn_in_rsci_d_mxwt[330];
  assign _05656_ = _05655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11493" *) chn_in_rsci_d_mxwt[331];
  assign _05657_ = _05656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11493" *) chn_in_rsci_d_mxwt[333];
  assign _05658_ = chn_in_rsci_d_mxwt[352] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11495" *) chn_in_rsci_d_mxwt[353];
  assign _05659_ = _05658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11496" *) chn_in_rsci_d_mxwt[354];
  assign _05660_ = _05659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11496" *) chn_in_rsci_d_mxwt[355];
  assign _05661_ = _05660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11496" *) chn_in_rsci_d_mxwt[356];
  assign _05662_ = _05661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11497" *) chn_in_rsci_d_mxwt[357];
  assign _05663_ = _05662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11497" *) chn_in_rsci_d_mxwt[358];
  assign _05664_ = _05663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11497" *) chn_in_rsci_d_mxwt[359];
  assign _05665_ = _05664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11498" *) chn_in_rsci_d_mxwt[360];
  assign _05666_ = _05665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11498" *) chn_in_rsci_d_mxwt[361];
  assign _05667_ = _05666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11498" *) chn_in_rsci_d_mxwt[362];
  assign _05668_ = _05667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11499" *) chn_in_rsci_d_mxwt[363];
  assign _05669_ = _05668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11499" *) chn_in_rsci_d_mxwt[365];
  assign _05670_ = chn_in_rsci_d_mxwt[384] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11501" *) chn_in_rsci_d_mxwt[385];
  assign _05671_ = _05670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11502" *) chn_in_rsci_d_mxwt[386];
  assign _05672_ = _05671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11502" *) chn_in_rsci_d_mxwt[387];
  assign _05673_ = _05672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11502" *) chn_in_rsci_d_mxwt[388];
  assign _05674_ = _05673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11503" *) chn_in_rsci_d_mxwt[389];
  assign _05675_ = _05674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11503" *) chn_in_rsci_d_mxwt[390];
  assign _05676_ = _05675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11503" *) chn_in_rsci_d_mxwt[391];
  assign _05677_ = _05676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11504" *) chn_in_rsci_d_mxwt[392];
  assign _05678_ = _05677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11504" *) chn_in_rsci_d_mxwt[393];
  assign _05679_ = _05678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11504" *) chn_in_rsci_d_mxwt[394];
  assign _05680_ = _05679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11505" *) chn_in_rsci_d_mxwt[395];
  assign _05681_ = _05680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11505" *) chn_in_rsci_d_mxwt[397];
  assign _05682_ = chn_in_rsci_d_mxwt[416] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11507" *) chn_in_rsci_d_mxwt[417];
  assign _05683_ = _05682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11508" *) chn_in_rsci_d_mxwt[418];
  assign _05684_ = _05683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11508" *) chn_in_rsci_d_mxwt[419];
  assign _05685_ = _05684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11508" *) chn_in_rsci_d_mxwt[420];
  assign _05686_ = _05685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11509" *) chn_in_rsci_d_mxwt[421];
  assign _05687_ = _05686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11509" *) chn_in_rsci_d_mxwt[422];
  assign _05688_ = _05687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11509" *) chn_in_rsci_d_mxwt[423];
  assign _05689_ = _05688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11510" *) chn_in_rsci_d_mxwt[424];
  assign _05690_ = _05689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11510" *) chn_in_rsci_d_mxwt[425];
  assign _05691_ = _05690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11510" *) chn_in_rsci_d_mxwt[426];
  assign _05692_ = _05691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11511" *) chn_in_rsci_d_mxwt[427];
  assign _05693_ = _05692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11511" *) chn_in_rsci_d_mxwt[429];
  assign _05694_ = chn_in_rsci_d_mxwt[448] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11513" *) chn_in_rsci_d_mxwt[449];
  assign _05695_ = _05694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11514" *) chn_in_rsci_d_mxwt[450];
  assign _05696_ = _05695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11514" *) chn_in_rsci_d_mxwt[451];
  assign _05697_ = _05696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11514" *) chn_in_rsci_d_mxwt[452];
  assign _05698_ = _05697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11515" *) chn_in_rsci_d_mxwt[453];
  assign _05699_ = _05698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11515" *) chn_in_rsci_d_mxwt[454];
  assign _05700_ = _05699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11515" *) chn_in_rsci_d_mxwt[455];
  assign _05701_ = _05700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11516" *) chn_in_rsci_d_mxwt[456];
  assign _05702_ = _05701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11516" *) chn_in_rsci_d_mxwt[457];
  assign _05703_ = _05702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11516" *) chn_in_rsci_d_mxwt[458];
  assign _05704_ = _05703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11517" *) chn_in_rsci_d_mxwt[459];
  assign _05705_ = _05704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11517" *) chn_in_rsci_d_mxwt[461];
  assign _05706_ = chn_in_rsci_d_mxwt[480] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11519" *) chn_in_rsci_d_mxwt[481];
  assign _05707_ = _05706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11519" *) chn_in_rsci_d_mxwt[482];
  assign _05708_ = _05707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11520" *) chn_in_rsci_d_mxwt[483];
  assign _05709_ = _05708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11520" *) chn_in_rsci_d_mxwt[484];
  assign _05710_ = _05709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11520" *) chn_in_rsci_d_mxwt[485];
  assign _05711_ = _05710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11521" *) chn_in_rsci_d_mxwt[486];
  assign _05712_ = _05711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11521" *) chn_in_rsci_d_mxwt[487];
  assign _05713_ = _05712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11521" *) chn_in_rsci_d_mxwt[488];
  assign _05714_ = _05713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *) chn_in_rsci_d_mxwt[489];
  assign _05715_ = _05714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *) chn_in_rsci_d_mxwt[490];
  assign _05716_ = _05715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *) chn_in_rsci_d_mxwt[491];
  assign _05717_ = _05716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11522" *) chn_in_rsci_d_mxwt[493];
  assign _05718_ = _04309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11524" *) _04024_;
  assign _05719_ = _04311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11531" *) _04026_;
  assign _05720_ = _04313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11538" *) _04028_;
  assign _05721_ = _04315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11545" *) _04030_;
  assign _05722_ = _04317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11552" *) _04032_;
  assign _05723_ = _04319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11559" *) _04034_;
  assign _05724_ = _04321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11566" *) _04036_;
  assign _05725_ = _04323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11573" *) _04038_;
  assign _05726_ = _04325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11580" *) _04040_;
  assign _05727_ = _04327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11587" *) _04042_;
  assign _05728_ = _04329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11594" *) _04044_;
  assign _05729_ = _04332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11608" *) _04047_;
  assign _05730_ = _04334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11615" *) _04049_;
  assign _05731_ = _04336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11622" *) _04051_;
  assign _05732_ = _04338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11629" *) _04053_;
  assign _05733_ = _01485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *) nand_164_cse;
  assign _05734_ = _04341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0 = _04342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11640" *) IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  assign _05735_ = _01486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *) nand_162_cse;
  assign _05736_ = _04344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0 = _04345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11646" *) IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  assign _05737_ = _01487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *) nand_160_cse;
  assign _05738_ = _04347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0 = _04348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11652" *) IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  assign _05739_ = _01488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *) nand_158_cse;
  assign _05740_ = _04350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0 = _04351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11658" *) IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  assign _05741_ = _01489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *) nand_156_cse;
  assign _05742_ = _04353_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0 = _04354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11664" *) nor_1099_cse;
  assign _05743_ = _01490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *) nand_153_cse;
  assign _05744_ = _04356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0 = _04357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11670" *) IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  assign _05745_ = _01491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *) nand_151_cse;
  assign _05746_ = _04359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0 = _04360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11676" *) IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  assign _05747_ = _01492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *) nand_149_cse;
  assign _05748_ = _04362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0 = _04363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11682" *) IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  assign _05749_ = _01493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *) nand_147_cse;
  assign _05750_ = _04365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0 = _04366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11688" *) IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  assign _05751_ = _01494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *) nand_145_cse;
  assign _05752_ = _04368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11694" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0 = _04369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11695" *) IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  assign _05753_ = _01495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *) nand_143_cse;
  assign _05754_ = _04371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11701" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0 = _04372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11702" *) IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  assign _05755_ = _01496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *) nand_141_cse;
  assign _05756_ = _04374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11708" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0 = _04375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11709" *) IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  assign _05757_ = _01497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *) nand_139_cse;
  assign _05758_ = _04377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11715" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0 = _04378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11716" *) IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  assign _05759_ = _01498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *) nand_137_cse;
  assign _05760_ = _04380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11722" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0 = _04381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11723" *) IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  assign _05761_ = _01499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *) nand_135_cse;
  assign _05762_ = _04383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11729" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0 = _04384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11730" *) IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  assign _05763_ = _01500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *) nand_133_cse;
  assign _05764_ = _04386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *) FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0 = _04387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11736" *) IsNaN_8U_23U_land_lpi_1_dfm_3;
  assign IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0 = _01501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11738" *) cvt_14_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _05765_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11898" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[1];
  assign _05766_ = _05765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11898" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[2];
  assign _05767_ = _05766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11899" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[3];
  assign _05768_ = _05767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11899" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[4];
  assign _05769_ = _05768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11900" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[5];
  assign _05770_ = _05769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11900" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[6];
  assign _05771_ = _05770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11901" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[7];
  assign _05772_ = _05771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11901" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[8];
  assign _05773_ = _05772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11902" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[9];
  assign _05774_ = _05773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11902" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[10];
  assign _05775_ = _05774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11903" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[11];
  assign _05776_ = _05775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11903" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[12];
  assign _05777_ = _05776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11904" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[13];
  assign _05778_ = _05777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11904" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[14];
  assign _05779_ = _05778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11905" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[15];
  assign _05780_ = _05779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11905" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[16];
  assign _05781_ = _05780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11906" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[17];
  assign _05782_ = _05781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11906" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[18];
  assign _05783_ = _05782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11907" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[19];
  assign _05784_ = _05783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11907" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[20];
  assign _05785_ = _05784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11908" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[21];
  assign _05786_ = _05785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11908" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[22];
  assign _05787_ = _05786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11909" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[23];
  assign _05788_ = _05787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11909" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[24];
  assign _05789_ = _05788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11910" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[25];
  assign _05790_ = _05789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11910" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[26];
  assign _05791_ = _05790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11911" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[27];
  assign _05792_ = _05791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11911" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[28];
  assign _05793_ = _05792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11912" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[29];
  assign _05794_ = _05793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11912" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[30];
  assign _05795_ = _05794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11913" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[31];
  assign _05796_ = _05795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11913" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[32];
  assign _05797_ = _05796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11914" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[33];
  assign _05798_ = _05797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11914" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[34];
  assign _05799_ = _05798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11915" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[35];
  assign _05800_ = _05799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11915" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[36];
  assign _05801_ = _05800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11916" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[37];
  assign _05802_ = _05801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11916" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[38];
  assign _05803_ = _05802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11917" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[39];
  assign _05804_ = _05803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11917" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[40];
  assign _05805_ = _05804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11918" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[41];
  assign _05806_ = _05805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11918" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[42];
  assign _05807_ = _05806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11919" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[43];
  assign _05808_ = _05807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11919" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[44];
  assign _05809_ = _05808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11920" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[45];
  assign _05810_ = _05809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11920" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[46];
  assign _05811_ = _05810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11921" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[47];
  assign _05812_ = _05811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11921" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[48];
  assign _05813_ = _05812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11922" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[49];
  assign _05814_ = _05813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11922" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[50];
  assign _05815_ = _05814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11923" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[51];
  assign _05816_ = _05815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11923" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[52];
  assign _05817_ = _05816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11924" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[53];
  assign _05818_ = _05817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11924" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[54];
  assign _05819_ = _05818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11925" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[55];
  assign _05820_ = _05819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11925" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[56];
  assign _05821_ = _05820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11926" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[57];
  assign _05822_ = _05821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11926" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[58];
  assign _05823_ = _05822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11927" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[59];
  assign _05824_ = _05823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11927" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[60];
  assign _05825_ = _05824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11928" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[61];
  assign _05826_ = _05825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11928" *) _04389_;
  assign _05319_ = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11935" *) _04391_;
  assign _05827_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11946" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[1];
  assign _05828_ = _05827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11946" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[2];
  assign _05829_ = _05828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11947" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[3];
  assign _05830_ = _05829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11947" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[4];
  assign _05831_ = _05830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11948" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[5];
  assign _05832_ = _05831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11948" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[6];
  assign _05833_ = _05832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11949" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[7];
  assign _05834_ = _05833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11949" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[8];
  assign _05835_ = _05834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11950" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[9];
  assign _05836_ = _05835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11950" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[10];
  assign _05837_ = _05836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11951" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[11];
  assign _05838_ = _05837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11951" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[12];
  assign _05839_ = _05838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11952" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[13];
  assign _05840_ = _05839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11952" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[14];
  assign _05841_ = _05840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11953" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[15];
  assign _05842_ = _05841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11953" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[16];
  assign _05843_ = _05842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11954" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[17];
  assign _05844_ = _05843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11954" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[18];
  assign _05845_ = _05844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11955" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[19];
  assign _05846_ = _05845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11955" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[20];
  assign _05847_ = _05846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11956" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[21];
  assign _05848_ = _05847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11956" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[22];
  assign _05849_ = _05848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11957" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[23];
  assign _05850_ = _05849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11957" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[24];
  assign _05851_ = _05850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11958" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[25];
  assign _05852_ = _05851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11958" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[26];
  assign _05853_ = _05852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11959" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[27];
  assign _05854_ = _05853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11959" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[28];
  assign _05855_ = _05854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11960" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[29];
  assign _05856_ = _05855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11960" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[30];
  assign _05857_ = _05856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11961" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[31];
  assign _05858_ = _05857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11961" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[32];
  assign _05859_ = _05858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11962" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[33];
  assign _05860_ = _05859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11962" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[34];
  assign _05861_ = _05860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11963" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[35];
  assign _05862_ = _05861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11963" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[36];
  assign _05863_ = _05862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11964" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[37];
  assign _05864_ = _05863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11964" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[38];
  assign _05865_ = _05864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11965" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[39];
  assign _05866_ = _05865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11965" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[40];
  assign _05867_ = _05866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11966" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[41];
  assign _05868_ = _05867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11966" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[42];
  assign _05869_ = _05868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11967" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[43];
  assign _05870_ = _05869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11967" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[44];
  assign _05871_ = _05870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11968" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[45];
  assign _05872_ = _05871_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11968" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[46];
  assign _05873_ = _05872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11969" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[47];
  assign _05874_ = _05873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11969" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[48];
  assign _05875_ = _05874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11970" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[49];
  assign _05876_ = _05875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11970" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[50];
  assign _05877_ = _05876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11971" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[51];
  assign _05878_ = _05877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11971" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[52];
  assign _05879_ = _05878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11972" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[53];
  assign _05880_ = _05879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11972" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[54];
  assign _05881_ = _05880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11973" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[55];
  assign _05882_ = _05881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11973" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[56];
  assign _05883_ = _05882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11974" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[57];
  assign _05884_ = _05883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11974" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[58];
  assign _05885_ = _05884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11975" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[59];
  assign _05886_ = _05885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11975" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[60];
  assign _05887_ = _05886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11976" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[61];
  assign _05888_ = _05887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11976" *) _04392_;
  assign _04857_ = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11983" *) _04394_;
  assign _05889_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11986" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[1];
  assign _05890_ = _05889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11986" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[2];
  assign _05891_ = _05890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11987" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[3];
  assign _05892_ = _05891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11987" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[4];
  assign _05893_ = _05892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11988" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[5];
  assign _05894_ = _05893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11988" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[6];
  assign _05895_ = _05894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11989" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[7];
  assign _05896_ = _05895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11989" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[8];
  assign _05897_ = _05896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11990" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[9];
  assign _05898_ = _05897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11990" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[10];
  assign _05899_ = _05898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11991" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[11];
  assign _05900_ = _05899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11991" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[12];
  assign _05901_ = _05900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11992" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[13];
  assign _05902_ = _05901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11992" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[14];
  assign _05903_ = _05902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11993" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[15];
  assign _05904_ = _05903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11993" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[16];
  assign _05905_ = _05904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11994" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[17];
  assign _05906_ = _05905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11994" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[18];
  assign _05907_ = _05906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11995" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[19];
  assign _05908_ = _05907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11995" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[20];
  assign _05909_ = _05908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11996" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[21];
  assign _05910_ = _05909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11996" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[22];
  assign _05911_ = _05910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11997" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[23];
  assign _05912_ = _05911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11997" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[24];
  assign _05913_ = _05912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11998" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[25];
  assign _05914_ = _05913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11998" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[26];
  assign _05915_ = _05914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11999" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[27];
  assign _05916_ = _05915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:11999" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[28];
  assign _05917_ = _05916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12000" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[29];
  assign _05918_ = _05917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12000" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[30];
  assign _05919_ = _05918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12001" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[31];
  assign _05920_ = _05919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12001" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[32];
  assign _05921_ = _05920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12002" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[33];
  assign _05922_ = _05921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12002" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[34];
  assign _05923_ = _05922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12003" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[35];
  assign _05924_ = _05923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12003" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[36];
  assign _05925_ = _05924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12004" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[37];
  assign _05926_ = _05925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12004" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[38];
  assign _05927_ = _05926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12005" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[39];
  assign _05928_ = _05927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12005" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[40];
  assign _05929_ = _05928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12006" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[41];
  assign _05930_ = _05929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12006" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[42];
  assign _05931_ = _05930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12007" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[43];
  assign _05932_ = _05931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12007" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[44];
  assign _05933_ = _05932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12008" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[45];
  assign _05934_ = _05933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12008" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[46];
  assign _05935_ = _05934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12009" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[47];
  assign _05936_ = _05935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12009" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[48];
  assign _05937_ = _05936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12010" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[49];
  assign _05938_ = _05937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12010" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[50];
  assign _05939_ = _05938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12011" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[51];
  assign _05940_ = _05939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12011" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[52];
  assign _05941_ = _05940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12012" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[53];
  assign _05942_ = _05941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12012" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[54];
  assign _05943_ = _05942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12013" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[55];
  assign _05944_ = _05943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12013" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[56];
  assign _05945_ = _05944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12014" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[57];
  assign _05946_ = _05945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12014" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[58];
  assign _05947_ = _05946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12015" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[59];
  assign _05948_ = _05947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12015" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[60];
  assign _05949_ = _05948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12016" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[61];
  assign _05950_ = _05949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12016" *) _04395_;
  assign _05320_ = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12023" *) _04397_;
  assign _05951_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12034" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[1];
  assign _05952_ = _05951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12034" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[2];
  assign _05953_ = _05952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12035" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[3];
  assign _05954_ = _05953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12035" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[4];
  assign _05955_ = _05954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12036" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[5];
  assign _05956_ = _05955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12036" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[6];
  assign _05957_ = _05956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12037" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[7];
  assign _05958_ = _05957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12037" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[8];
  assign _05959_ = _05958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12038" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[9];
  assign _05960_ = _05959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12038" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[10];
  assign _05961_ = _05960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12039" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[11];
  assign _05962_ = _05961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12039" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[12];
  assign _05963_ = _05962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12040" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[13];
  assign _05964_ = _05963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12040" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[14];
  assign _05965_ = _05964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12041" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[15];
  assign _05966_ = _05965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12041" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[16];
  assign _05967_ = _05966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12042" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[17];
  assign _05968_ = _05967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12042" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[18];
  assign _05969_ = _05968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12043" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[19];
  assign _05970_ = _05969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12043" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[20];
  assign _05971_ = _05970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12044" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[21];
  assign _05972_ = _05971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12044" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[22];
  assign _05973_ = _05972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12045" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[23];
  assign _05974_ = _05973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12045" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[24];
  assign _05975_ = _05974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12046" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[25];
  assign _05976_ = _05975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12046" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[26];
  assign _05977_ = _05976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12047" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[27];
  assign _05978_ = _05977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12047" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[28];
  assign _05979_ = _05978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12048" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[29];
  assign _05980_ = _05979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12048" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[30];
  assign _05981_ = _05980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12049" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[31];
  assign _05982_ = _05981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12049" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[32];
  assign _05983_ = _05982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12050" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[33];
  assign _05984_ = _05983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12050" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[34];
  assign _05985_ = _05984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12051" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[35];
  assign _05986_ = _05985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12051" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[36];
  assign _05987_ = _05986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12052" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[37];
  assign _05988_ = _05987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12052" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[38];
  assign _05989_ = _05988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12053" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[39];
  assign _05990_ = _05989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12053" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[40];
  assign _05991_ = _05990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12054" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[41];
  assign _05992_ = _05991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12054" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[42];
  assign _05993_ = _05992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12055" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[43];
  assign _05994_ = _05993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12055" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[44];
  assign _05995_ = _05994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12056" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[45];
  assign _05996_ = _05995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12056" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[46];
  assign _05997_ = _05996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12057" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[47];
  assign _05998_ = _05997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12057" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[48];
  assign _05999_ = _05998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12058" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[49];
  assign _06000_ = _05999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12058" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[50];
  assign _06001_ = _06000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12059" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[51];
  assign _06002_ = _06001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12059" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[52];
  assign _06003_ = _06002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12060" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[53];
  assign _06004_ = _06003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12060" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[54];
  assign _06005_ = _06004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12061" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[55];
  assign _06006_ = _06005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12061" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[56];
  assign _06007_ = _06006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12062" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[57];
  assign _06008_ = _06007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12062" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[58];
  assign _06009_ = _06008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12063" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[59];
  assign _06010_ = _06009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12063" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[60];
  assign _06011_ = _06010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12064" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[61];
  assign _06012_ = _06011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12064" *) _04398_;
  assign _04860_ = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12071" *) _04400_;
  assign _06013_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12082" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[1];
  assign _06014_ = _06013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12082" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[2];
  assign _06015_ = _06014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12083" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[3];
  assign _06016_ = _06015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12083" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[4];
  assign _06017_ = _06016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12084" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[5];
  assign _06018_ = _06017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12084" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[6];
  assign _06019_ = _06018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12085" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[7];
  assign _06020_ = _06019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12085" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[8];
  assign _06021_ = _06020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12086" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[9];
  assign _06022_ = _06021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12086" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[10];
  assign _06023_ = _06022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12087" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[11];
  assign _06024_ = _06023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12087" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[12];
  assign _06025_ = _06024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12088" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[13];
  assign _06026_ = _06025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12088" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[14];
  assign _06027_ = _06026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12089" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[15];
  assign _06028_ = _06027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12089" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[16];
  assign _06029_ = _06028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12090" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[17];
  assign _06030_ = _06029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12090" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[18];
  assign _06031_ = _06030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12091" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[19];
  assign _06032_ = _06031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12091" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[20];
  assign _06033_ = _06032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12092" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[21];
  assign _06034_ = _06033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12092" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[22];
  assign _06035_ = _06034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12093" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[23];
  assign _06036_ = _06035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12093" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[24];
  assign _06037_ = _06036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12094" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[25];
  assign _06038_ = _06037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12094" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[26];
  assign _06039_ = _06038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12095" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[27];
  assign _06040_ = _06039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12095" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[28];
  assign _06041_ = _06040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12096" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[29];
  assign _06042_ = _06041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12096" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[30];
  assign _06043_ = _06042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12097" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[31];
  assign _06044_ = _06043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12097" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[32];
  assign _06045_ = _06044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12098" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[33];
  assign _06046_ = _06045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12098" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[34];
  assign _06047_ = _06046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12099" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[35];
  assign _06048_ = _06047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12099" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[36];
  assign _06049_ = _06048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12100" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[37];
  assign _06050_ = _06049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12100" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[38];
  assign _06051_ = _06050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12101" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[39];
  assign _06052_ = _06051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12101" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[40];
  assign _06053_ = _06052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12102" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[41];
  assign _06054_ = _06053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12102" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[42];
  assign _06055_ = _06054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12103" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[43];
  assign _06056_ = _06055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12103" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[44];
  assign _06057_ = _06056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12104" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[45];
  assign _06058_ = _06057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12104" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[46];
  assign _06059_ = _06058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12105" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[47];
  assign _06060_ = _06059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12105" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[48];
  assign _06061_ = _06060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12106" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[49];
  assign _06062_ = _06061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12106" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[50];
  assign _06063_ = _06062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12107" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[51];
  assign _06064_ = _06063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12107" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[52];
  assign _06065_ = _06064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12108" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[53];
  assign _06066_ = _06065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12108" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[54];
  assign _06067_ = _06066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12109" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[55];
  assign _06068_ = _06067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12109" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[56];
  assign _06069_ = _06068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12110" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[57];
  assign _06070_ = _06069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12110" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[58];
  assign _06071_ = _06070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12111" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[59];
  assign _06072_ = _06071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12111" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[60];
  assign _06073_ = _06072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12112" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[61];
  assign _06074_ = _06073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12112" *) _04401_;
  assign _04863_ = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12119" *) _04403_;
  assign _06075_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12122" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[1];
  assign _06076_ = _06075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12122" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[2];
  assign _06077_ = _06076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12123" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[3];
  assign _06078_ = _06077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12123" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[4];
  assign _06079_ = _06078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12124" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[5];
  assign _06080_ = _06079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12124" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[6];
  assign _06081_ = _06080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12125" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[7];
  assign _06082_ = _06081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12125" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[8];
  assign _06083_ = _06082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12126" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[9];
  assign _06084_ = _06083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12126" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[10];
  assign _06085_ = _06084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12127" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[11];
  assign _06086_ = _06085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12127" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[12];
  assign _06087_ = _06086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12128" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[13];
  assign _06088_ = _06087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12128" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[14];
  assign _06089_ = _06088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12129" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[15];
  assign _06090_ = _06089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12129" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[16];
  assign _06091_ = _06090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12130" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[17];
  assign _06092_ = _06091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12130" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[18];
  assign _06093_ = _06092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12131" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[19];
  assign _06094_ = _06093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12131" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[20];
  assign _06095_ = _06094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12132" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[21];
  assign _06096_ = _06095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12132" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[22];
  assign _06097_ = _06096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12133" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[23];
  assign _06098_ = _06097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12133" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[24];
  assign _06099_ = _06098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12134" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[25];
  assign _06100_ = _06099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12134" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[26];
  assign _06101_ = _06100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12135" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[27];
  assign _06102_ = _06101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12135" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[28];
  assign _06103_ = _06102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12136" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[29];
  assign _06104_ = _06103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12136" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[30];
  assign _06105_ = _06104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12137" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[31];
  assign _06106_ = _06105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12137" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[32];
  assign _06107_ = _06106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12138" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[33];
  assign _06108_ = _06107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12138" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[34];
  assign _06109_ = _06108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12139" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[35];
  assign _06110_ = _06109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12139" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[36];
  assign _06111_ = _06110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12140" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[37];
  assign _06112_ = _06111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12140" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[38];
  assign _06113_ = _06112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12141" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[39];
  assign _06114_ = _06113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12141" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[40];
  assign _06115_ = _06114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12142" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[41];
  assign _06116_ = _06115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12142" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[42];
  assign _06117_ = _06116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12143" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[43];
  assign _06118_ = _06117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12143" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[44];
  assign _06119_ = _06118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12144" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[45];
  assign _06120_ = _06119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12144" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[46];
  assign _06121_ = _06120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12145" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[47];
  assign _06122_ = _06121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12145" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[48];
  assign _06123_ = _06122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12146" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[49];
  assign _06124_ = _06123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12146" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[50];
  assign _06125_ = _06124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12147" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[51];
  assign _06126_ = _06125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12147" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[52];
  assign _06127_ = _06126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12148" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[53];
  assign _06128_ = _06127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12148" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[54];
  assign _06129_ = _06128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12149" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[55];
  assign _06130_ = _06129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12149" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[56];
  assign _06131_ = _06130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12150" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[57];
  assign _06132_ = _06131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12150" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[58];
  assign _06133_ = _06132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12151" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[59];
  assign _06134_ = _06133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12151" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[60];
  assign _06135_ = _06134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12152" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[61];
  assign _06136_ = _06135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12152" *) _04404_;
  assign _04861_ = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12159" *) _04406_;
  assign _06137_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12162" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[1];
  assign _06138_ = _06137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12162" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[2];
  assign _06139_ = _06138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12163" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[3];
  assign _06140_ = _06139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12163" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[4];
  assign _06141_ = _06140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12164" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[5];
  assign _06142_ = _06141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12164" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[6];
  assign _06143_ = _06142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12165" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[7];
  assign _06144_ = _06143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12165" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[8];
  assign _06145_ = _06144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12166" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[9];
  assign _06146_ = _06145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12166" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[10];
  assign _06147_ = _06146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12167" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[11];
  assign _06148_ = _06147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12167" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[12];
  assign _06149_ = _06148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12168" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[13];
  assign _06150_ = _06149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12168" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[14];
  assign _06151_ = _06150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12169" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[15];
  assign _06152_ = _06151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12169" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[16];
  assign _06153_ = _06152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12170" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[17];
  assign _06154_ = _06153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12170" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[18];
  assign _06155_ = _06154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12171" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[19];
  assign _06156_ = _06155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12171" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[20];
  assign _06157_ = _06156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12172" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[21];
  assign _06158_ = _06157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12172" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[22];
  assign _06159_ = _06158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12173" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[23];
  assign _06160_ = _06159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12173" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[24];
  assign _06161_ = _06160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12174" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[25];
  assign _06162_ = _06161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12174" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[26];
  assign _06163_ = _06162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12175" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[27];
  assign _06164_ = _06163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12175" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[28];
  assign _06165_ = _06164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12176" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[29];
  assign _06166_ = _06165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12176" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[30];
  assign _06167_ = _06166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12177" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[31];
  assign _06168_ = _06167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12177" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[32];
  assign _06169_ = _06168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12178" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[33];
  assign _06170_ = _06169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12178" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[34];
  assign _06171_ = _06170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12179" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[35];
  assign _06172_ = _06171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12179" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[36];
  assign _06173_ = _06172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12180" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[37];
  assign _06174_ = _06173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12180" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[38];
  assign _06175_ = _06174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12181" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[39];
  assign _06176_ = _06175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12181" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[40];
  assign _06177_ = _06176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12182" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[41];
  assign _06178_ = _06177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12182" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[42];
  assign _06179_ = _06178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12183" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[43];
  assign _06180_ = _06179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12183" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[44];
  assign _06181_ = _06180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12184" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[45];
  assign _06182_ = _06181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12184" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[46];
  assign _06183_ = _06182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12185" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[47];
  assign _06184_ = _06183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12185" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[48];
  assign _06185_ = _06184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12186" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[49];
  assign _06186_ = _06185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12186" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[50];
  assign _06187_ = _06186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12187" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[51];
  assign _06188_ = _06187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12187" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[52];
  assign _06189_ = _06188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12188" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[53];
  assign _06190_ = _06189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12188" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[54];
  assign _06191_ = _06190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12189" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[55];
  assign _06192_ = _06191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12189" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[56];
  assign _06193_ = _06192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12190" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[57];
  assign _06194_ = _06193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12190" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[58];
  assign _06195_ = _06194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12191" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[59];
  assign _06196_ = _06195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12191" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[60];
  assign _06197_ = _06196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12192" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[61];
  assign _06198_ = _06197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12192" *) _04407_;
  assign _04859_ = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12199" *) _04409_;
  assign _06199_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12210" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[1];
  assign _06200_ = _06199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12210" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[2];
  assign _06201_ = _06200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12211" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[3];
  assign _06202_ = _06201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12211" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[4];
  assign _06203_ = _06202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12212" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[5];
  assign _06204_ = _06203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12212" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[6];
  assign _06205_ = _06204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12213" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[7];
  assign _06206_ = _06205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12213" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[8];
  assign _06207_ = _06206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12214" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[9];
  assign _06208_ = _06207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12214" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[10];
  assign _06209_ = _06208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12215" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[11];
  assign _06210_ = _06209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12215" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[12];
  assign _06211_ = _06210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12216" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[13];
  assign _06212_ = _06211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12216" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[14];
  assign _06213_ = _06212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12217" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[15];
  assign _06214_ = _06213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12217" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[16];
  assign _06215_ = _06214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12218" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[17];
  assign _06216_ = _06215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12218" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[18];
  assign _06217_ = _06216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12219" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[19];
  assign _06218_ = _06217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12219" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[20];
  assign _06219_ = _06218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12220" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[21];
  assign _06220_ = _06219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12220" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[22];
  assign _06221_ = _06220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12221" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[23];
  assign _06222_ = _06221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12221" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[24];
  assign _06223_ = _06222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12222" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[25];
  assign _06224_ = _06223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12222" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[26];
  assign _06225_ = _06224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12223" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[27];
  assign _06226_ = _06225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12223" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[28];
  assign _06227_ = _06226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12224" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[29];
  assign _06228_ = _06227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12224" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[30];
  assign _06229_ = _06228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12225" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[31];
  assign _06230_ = _06229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12225" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[32];
  assign _06231_ = _06230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12226" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[33];
  assign _06232_ = _06231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12226" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[34];
  assign _06233_ = _06232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12227" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[35];
  assign _06234_ = _06233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12227" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[36];
  assign _06235_ = _06234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12228" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[37];
  assign _06236_ = _06235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12228" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[38];
  assign _06237_ = _06236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12229" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[39];
  assign _06238_ = _06237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12229" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[40];
  assign _06239_ = _06238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12230" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[41];
  assign _06240_ = _06239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12230" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[42];
  assign _06241_ = _06240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12231" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[43];
  assign _06242_ = _06241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12231" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[44];
  assign _06243_ = _06242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12232" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[45];
  assign _06244_ = _06243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12232" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[46];
  assign _06245_ = _06244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12233" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[47];
  assign _06246_ = _06245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12233" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[48];
  assign _06247_ = _06246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12234" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[49];
  assign _06248_ = _06247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12234" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[50];
  assign _06249_ = _06248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12235" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[51];
  assign _06250_ = _06249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12235" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[52];
  assign _06251_ = _06250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12236" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[53];
  assign _06252_ = _06251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12236" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[54];
  assign _06253_ = _06252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12237" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[55];
  assign _06254_ = _06253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12237" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[56];
  assign _06255_ = _06254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12238" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[57];
  assign _06256_ = _06255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12238" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[58];
  assign _06257_ = _06256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12239" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[59];
  assign _06258_ = _06257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12239" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[60];
  assign _06259_ = _06258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12240" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[61];
  assign _06260_ = _06259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12240" *) _04410_;
  assign _04864_ = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12247" *) _04412_;
  assign _06261_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12258" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[1];
  assign _06262_ = _06261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12258" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[2];
  assign _06263_ = _06262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12259" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[3];
  assign _06264_ = _06263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12259" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[4];
  assign _06265_ = _06264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12260" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[5];
  assign _06266_ = _06265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12260" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[6];
  assign _06267_ = _06266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12261" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[7];
  assign _06268_ = _06267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12261" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[8];
  assign _06269_ = _06268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12262" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[9];
  assign _06270_ = _06269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12262" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[10];
  assign _06271_ = _06270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12263" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[11];
  assign _06272_ = _06271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12263" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[12];
  assign _06273_ = _06272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12264" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[13];
  assign _06274_ = _06273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12264" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[14];
  assign _06275_ = _06274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12265" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[15];
  assign _06276_ = _06275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12265" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[16];
  assign _06277_ = _06276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12266" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[17];
  assign _06278_ = _06277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12266" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[18];
  assign _06279_ = _06278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12267" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[19];
  assign _06280_ = _06279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12267" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[20];
  assign _06281_ = _06280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12268" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[21];
  assign _06282_ = _06281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12268" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[22];
  assign _06283_ = _06282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12269" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[23];
  assign _06284_ = _06283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12269" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[24];
  assign _06285_ = _06284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12270" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[25];
  assign _06286_ = _06285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12270" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[26];
  assign _06287_ = _06286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12271" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[27];
  assign _06288_ = _06287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12271" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[28];
  assign _06289_ = _06288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12272" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[29];
  assign _06290_ = _06289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12272" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[30];
  assign _06291_ = _06290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12273" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[31];
  assign _06292_ = _06291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12273" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[32];
  assign _06293_ = _06292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12274" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[33];
  assign _06294_ = _06293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12274" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[34];
  assign _06295_ = _06294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12275" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[35];
  assign _06296_ = _06295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12275" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[36];
  assign _06297_ = _06296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12276" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[37];
  assign _06298_ = _06297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12276" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[38];
  assign _06299_ = _06298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12277" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[39];
  assign _06300_ = _06299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12277" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[40];
  assign _06301_ = _06300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12278" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[41];
  assign _06302_ = _06301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12278" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[42];
  assign _06303_ = _06302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12279" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[43];
  assign _06304_ = _06303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12279" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[44];
  assign _06305_ = _06304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12280" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[45];
  assign _06306_ = _06305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12280" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[46];
  assign _06307_ = _06306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12281" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[47];
  assign _06308_ = _06307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12281" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[48];
  assign _06309_ = _06308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12282" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[49];
  assign _06310_ = _06309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12282" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[50];
  assign _06311_ = _06310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12283" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[51];
  assign _06312_ = _06311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12283" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[52];
  assign _06313_ = _06312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12284" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[53];
  assign _06314_ = _06313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12284" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[54];
  assign _06315_ = _06314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12285" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[55];
  assign _06316_ = _06315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12285" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[56];
  assign _06317_ = _06316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12286" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[57];
  assign _06318_ = _06317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12286" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[58];
  assign _06319_ = _06318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12287" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[59];
  assign _06320_ = _06319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12287" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[60];
  assign _06321_ = _06320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12288" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[61];
  assign _06322_ = _06321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12288" *) _04413_;
  assign _04866_ = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12295" *) _04415_;
  assign _06323_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12298" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[1];
  assign _06324_ = _06323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12298" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[2];
  assign _06325_ = _06324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12299" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[3];
  assign _06326_ = _06325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12299" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[4];
  assign _06327_ = _06326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12300" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[5];
  assign _06328_ = _06327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12300" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[6];
  assign _06329_ = _06328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12301" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[7];
  assign _06330_ = _06329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12301" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[8];
  assign _06331_ = _06330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12302" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[9];
  assign _06332_ = _06331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12302" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[10];
  assign _06333_ = _06332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12303" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[11];
  assign _06334_ = _06333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12303" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[12];
  assign _06335_ = _06334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12304" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[13];
  assign _06336_ = _06335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12304" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[14];
  assign _06337_ = _06336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12305" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[15];
  assign _06338_ = _06337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12305" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[16];
  assign _06339_ = _06338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12306" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[17];
  assign _06340_ = _06339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12306" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[18];
  assign _06341_ = _06340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12307" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[19];
  assign _06342_ = _06341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12307" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[20];
  assign _06343_ = _06342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12308" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[21];
  assign _06344_ = _06343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12308" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[22];
  assign _06345_ = _06344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12309" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[23];
  assign _06346_ = _06345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12309" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[24];
  assign _06347_ = _06346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12310" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[25];
  assign _06348_ = _06347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12310" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[26];
  assign _06349_ = _06348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12311" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[27];
  assign _06350_ = _06349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12311" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[28];
  assign _06351_ = _06350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12312" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[29];
  assign _06352_ = _06351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12312" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[30];
  assign _06353_ = _06352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12313" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[31];
  assign _06354_ = _06353_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12313" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[32];
  assign _06355_ = _06354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12314" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[33];
  assign _06356_ = _06355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12314" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[34];
  assign _06357_ = _06356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12315" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[35];
  assign _06358_ = _06357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12315" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[36];
  assign _06359_ = _06358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12316" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[37];
  assign _06360_ = _06359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12316" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[38];
  assign _06361_ = _06360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12317" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[39];
  assign _06362_ = _06361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12317" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[40];
  assign _06363_ = _06362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12318" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[41];
  assign _06364_ = _06363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12318" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[42];
  assign _06365_ = _06364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12319" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[43];
  assign _06366_ = _06365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12319" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[44];
  assign _06367_ = _06366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12320" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[45];
  assign _06368_ = _06367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12320" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[46];
  assign _06369_ = _06368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12321" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[47];
  assign _06370_ = _06369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12321" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[48];
  assign _06371_ = _06370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12322" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[49];
  assign _06372_ = _06371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12322" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[50];
  assign _06373_ = _06372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12323" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[51];
  assign _06374_ = _06373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12323" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[52];
  assign _06375_ = _06374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12324" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[53];
  assign _06376_ = _06375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12324" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[54];
  assign _06377_ = _06376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12325" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[55];
  assign _06378_ = _06377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12325" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[56];
  assign _06379_ = _06378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12326" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[57];
  assign _06380_ = _06379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12326" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[58];
  assign _06381_ = _06380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12327" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[59];
  assign _06382_ = _06381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12327" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[60];
  assign _06383_ = _06382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12328" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[61];
  assign _06384_ = _06383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12328" *) _04416_;
  assign _04865_ = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12335" *) _04418_;
  assign _06385_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12346" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[1];
  assign _06386_ = _06385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12346" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[2];
  assign _06387_ = _06386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12347" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[3];
  assign _06388_ = _06387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12347" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[4];
  assign _06389_ = _06388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12348" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[5];
  assign _06390_ = _06389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12348" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[6];
  assign _06391_ = _06390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12349" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[7];
  assign _06392_ = _06391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12349" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[8];
  assign _06393_ = _06392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12350" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[9];
  assign _06394_ = _06393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12350" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[10];
  assign _06395_ = _06394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12351" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[11];
  assign _06396_ = _06395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12351" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[12];
  assign _06397_ = _06396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12352" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[13];
  assign _06398_ = _06397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12352" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[14];
  assign _06399_ = _06398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12353" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[15];
  assign _06400_ = _06399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12353" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[16];
  assign _06401_ = _06400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12354" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[17];
  assign _06402_ = _06401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12354" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[18];
  assign _06403_ = _06402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12355" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[19];
  assign _06404_ = _06403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12355" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[20];
  assign _06405_ = _06404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12356" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[21];
  assign _06406_ = _06405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12356" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[22];
  assign _06407_ = _06406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12357" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[23];
  assign _06408_ = _06407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12357" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[24];
  assign _06409_ = _06408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12358" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[25];
  assign _06410_ = _06409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12358" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[26];
  assign _06411_ = _06410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12359" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[27];
  assign _06412_ = _06411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12359" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[28];
  assign _06413_ = _06412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12360" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[29];
  assign _06414_ = _06413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12360" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[30];
  assign _06415_ = _06414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12361" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[31];
  assign _06416_ = _06415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12361" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[32];
  assign _06417_ = _06416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12362" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[33];
  assign _06418_ = _06417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12362" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[34];
  assign _06419_ = _06418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12363" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[35];
  assign _06420_ = _06419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12363" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[36];
  assign _06421_ = _06420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12364" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[37];
  assign _06422_ = _06421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12364" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[38];
  assign _06423_ = _06422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12365" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[39];
  assign _06424_ = _06423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12365" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[40];
  assign _06425_ = _06424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12366" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[41];
  assign _06426_ = _06425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12366" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[42];
  assign _06427_ = _06426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12367" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[43];
  assign _06428_ = _06427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12367" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[44];
  assign _06429_ = _06428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12368" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[45];
  assign _06430_ = _06429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12368" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[46];
  assign _06431_ = _06430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12369" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[47];
  assign _06432_ = _06431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12369" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[48];
  assign _06433_ = _06432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12370" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[49];
  assign _06434_ = _06433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12370" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[50];
  assign _06435_ = _06434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12371" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[51];
  assign _06436_ = _06435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12371" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[52];
  assign _06437_ = _06436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12372" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[53];
  assign _06438_ = _06437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12372" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[54];
  assign _06439_ = _06438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12373" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[55];
  assign _06440_ = _06439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12373" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[56];
  assign _06441_ = _06440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12374" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[57];
  assign _06442_ = _06441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12374" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[58];
  assign _06443_ = _06442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12375" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[59];
  assign _06444_ = _06443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12375" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[60];
  assign _06445_ = _06444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12376" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[61];
  assign _06446_ = _06445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12376" *) _04419_;
  assign _04869_ = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12383" *) _04421_;
  assign _06447_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12394" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[1];
  assign _06448_ = _06447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12394" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[2];
  assign _06449_ = _06448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12395" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[3];
  assign _06450_ = _06449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12395" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[4];
  assign _06451_ = _06450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12396" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[5];
  assign _06452_ = _06451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12396" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[6];
  assign _06453_ = _06452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12397" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[7];
  assign _06454_ = _06453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12397" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[8];
  assign _06455_ = _06454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12398" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[9];
  assign _06456_ = _06455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12398" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[10];
  assign _06457_ = _06456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12399" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[11];
  assign _06458_ = _06457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12399" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[12];
  assign _06459_ = _06458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12400" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[13];
  assign _06460_ = _06459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12400" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[14];
  assign _06461_ = _06460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12401" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[15];
  assign _06462_ = _06461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12401" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[16];
  assign _06463_ = _06462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12402" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[17];
  assign _06464_ = _06463_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12402" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[18];
  assign _06465_ = _06464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12403" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[19];
  assign _06466_ = _06465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12403" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[20];
  assign _06467_ = _06466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12404" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[21];
  assign _06468_ = _06467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12404" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[22];
  assign _06469_ = _06468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12405" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[23];
  assign _06470_ = _06469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12405" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[24];
  assign _06471_ = _06470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12406" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[25];
  assign _06472_ = _06471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12406" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[26];
  assign _06473_ = _06472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12407" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[27];
  assign _06474_ = _06473_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12407" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[28];
  assign _06475_ = _06474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12408" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[29];
  assign _06476_ = _06475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12408" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[30];
  assign _06477_ = _06476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12409" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[31];
  assign _06478_ = _06477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12409" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[32];
  assign _06479_ = _06478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12410" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[33];
  assign _06480_ = _06479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12410" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[34];
  assign _06481_ = _06480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12411" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[35];
  assign _06482_ = _06481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12411" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[36];
  assign _06483_ = _06482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12412" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[37];
  assign _06484_ = _06483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12412" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[38];
  assign _06485_ = _06484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12413" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[39];
  assign _06486_ = _06485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12413" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[40];
  assign _06487_ = _06486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12414" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[41];
  assign _06488_ = _06487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12414" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[42];
  assign _06489_ = _06488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12415" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[43];
  assign _06490_ = _06489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12415" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[44];
  assign _06491_ = _06490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12416" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[45];
  assign _06492_ = _06491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12416" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[46];
  assign _06493_ = _06492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12417" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[47];
  assign _06494_ = _06493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12417" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[48];
  assign _06495_ = _06494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12418" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[49];
  assign _06496_ = _06495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12418" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[50];
  assign _06497_ = _06496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12419" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[51];
  assign _06498_ = _06497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12419" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[52];
  assign _06499_ = _06498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12420" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[53];
  assign _06500_ = _06499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12420" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[54];
  assign _06501_ = _06500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12421" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[55];
  assign _06502_ = _06501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12421" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[56];
  assign _06503_ = _06502_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12422" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[57];
  assign _06504_ = _06503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12422" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[58];
  assign _06505_ = _06504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12423" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[59];
  assign _06506_ = _06505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12423" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[60];
  assign _06507_ = _06506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12424" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[61];
  assign _06508_ = _06507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12424" *) _04422_;
  assign _04873_ = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12431" *) _04424_;
  assign _06509_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12434" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[1];
  assign _06510_ = _06509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12434" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[2];
  assign _06511_ = _06510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12435" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[3];
  assign _06512_ = _06511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12435" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[4];
  assign _06513_ = _06512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12436" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[5];
  assign _06514_ = _06513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12436" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[6];
  assign _06515_ = _06514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12437" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[7];
  assign _06516_ = _06515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12437" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[8];
  assign _06517_ = _06516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12438" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[9];
  assign _06518_ = _06517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12438" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[10];
  assign _06519_ = _06518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12439" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[11];
  assign _06520_ = _06519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12439" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[12];
  assign _06521_ = _06520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12440" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[13];
  assign _06522_ = _06521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12440" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[14];
  assign _06523_ = _06522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12441" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[15];
  assign _06524_ = _06523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12441" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[16];
  assign _06525_ = _06524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12442" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[17];
  assign _06526_ = _06525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12442" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[18];
  assign _06527_ = _06526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12443" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[19];
  assign _06528_ = _06527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12443" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[20];
  assign _06529_ = _06528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12444" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[21];
  assign _06530_ = _06529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12444" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[22];
  assign _06531_ = _06530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12445" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[23];
  assign _06532_ = _06531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12445" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[24];
  assign _06533_ = _06532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12446" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[25];
  assign _06534_ = _06533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12446" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[26];
  assign _06535_ = _06534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12447" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[27];
  assign _06536_ = _06535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12447" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[28];
  assign _06537_ = _06536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12448" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[29];
  assign _06538_ = _06537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12448" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[30];
  assign _06539_ = _06538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12449" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[31];
  assign _06540_ = _06539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12449" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[32];
  assign _06541_ = _06540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12450" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[33];
  assign _06542_ = _06541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12450" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[34];
  assign _06543_ = _06542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12451" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[35];
  assign _06544_ = _06543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12451" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[36];
  assign _06545_ = _06544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12452" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[37];
  assign _06546_ = _06545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12452" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[38];
  assign _06547_ = _06546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12453" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[39];
  assign _06548_ = _06547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12453" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[40];
  assign _06549_ = _06548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12454" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[41];
  assign _06550_ = _06549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12454" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[42];
  assign _06551_ = _06550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12455" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[43];
  assign _06552_ = _06551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12455" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[44];
  assign _06553_ = _06552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12456" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[45];
  assign _06554_ = _06553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12456" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[46];
  assign _06555_ = _06554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12457" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[47];
  assign _06556_ = _06555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12457" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[48];
  assign _06557_ = _06556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12458" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[49];
  assign _06558_ = _06557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12458" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[50];
  assign _06559_ = _06558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12459" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[51];
  assign _06560_ = _06559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12459" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[52];
  assign _06561_ = _06560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12460" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[53];
  assign _06562_ = _06561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12460" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[54];
  assign _06563_ = _06562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12461" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[55];
  assign _06564_ = _06563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12461" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[56];
  assign _06565_ = _06564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12462" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[57];
  assign _06566_ = _06565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12462" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[58];
  assign _06567_ = _06566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12463" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[59];
  assign _06568_ = _06567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12463" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[60];
  assign _06569_ = _06568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12464" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[61];
  assign _06570_ = _06569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12464" *) _04425_;
  assign _04871_ = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12471" *) _04427_;
  assign _06571_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12474" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[1];
  assign _06572_ = _06571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12474" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[2];
  assign _06573_ = _06572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12475" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[3];
  assign _06574_ = _06573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12475" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[4];
  assign _06575_ = _06574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12476" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[5];
  assign _06576_ = _06575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12476" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[6];
  assign _06577_ = _06576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12477" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[7];
  assign _06578_ = _06577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12477" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[8];
  assign _06579_ = _06578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12478" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[9];
  assign _06580_ = _06579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12478" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[10];
  assign _06581_ = _06580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12479" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[11];
  assign _06582_ = _06581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12479" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[12];
  assign _06583_ = _06582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12480" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[13];
  assign _06584_ = _06583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12480" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[14];
  assign _06585_ = _06584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12481" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[15];
  assign _06586_ = _06585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12481" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[16];
  assign _06587_ = _06586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12482" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[17];
  assign _06588_ = _06587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12482" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[18];
  assign _06589_ = _06588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12483" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[19];
  assign _06590_ = _06589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12483" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[20];
  assign _06591_ = _06590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12484" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[21];
  assign _06592_ = _06591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12484" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[22];
  assign _06593_ = _06592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12485" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[23];
  assign _06594_ = _06593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12485" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[24];
  assign _06595_ = _06594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12486" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[25];
  assign _06596_ = _06595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12486" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[26];
  assign _06597_ = _06596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12487" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[27];
  assign _06598_ = _06597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12487" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[28];
  assign _06599_ = _06598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12488" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[29];
  assign _06600_ = _06599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12488" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[30];
  assign _06601_ = _06600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12489" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[31];
  assign _06602_ = _06601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12489" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[32];
  assign _06603_ = _06602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12490" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[33];
  assign _06604_ = _06603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12490" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[34];
  assign _06605_ = _06604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12491" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[35];
  assign _06606_ = _06605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12491" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[36];
  assign _06607_ = _06606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12492" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[37];
  assign _06608_ = _06607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12492" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[38];
  assign _06609_ = _06608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12493" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[39];
  assign _06610_ = _06609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12493" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[40];
  assign _06611_ = _06610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12494" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[41];
  assign _06612_ = _06611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12494" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[42];
  assign _06613_ = _06612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12495" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[43];
  assign _06614_ = _06613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12495" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[44];
  assign _06615_ = _06614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12496" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[45];
  assign _06616_ = _06615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12496" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[46];
  assign _06617_ = _06616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12497" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[47];
  assign _06618_ = _06617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12497" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[48];
  assign _06619_ = _06618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12498" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[49];
  assign _06620_ = _06619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12498" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[50];
  assign _06621_ = _06620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12499" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[51];
  assign _06622_ = _06621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12499" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[52];
  assign _06623_ = _06622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12500" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[53];
  assign _06624_ = _06623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12500" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[54];
  assign _06625_ = _06624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12501" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[55];
  assign _06626_ = _06625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12501" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[56];
  assign _06627_ = _06626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12502" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[57];
  assign _06628_ = _06627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12502" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[58];
  assign _06629_ = _06628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12503" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[59];
  assign _06630_ = _06629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12503" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[60];
  assign _06631_ = _06630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12504" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[61];
  assign _06632_ = _06631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12504" *) _04428_;
  assign _04868_ = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12511" *) _04430_;
  assign _06633_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12514" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[1];
  assign _06634_ = _06633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12514" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[2];
  assign _06635_ = _06634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12515" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[3];
  assign _06636_ = _06635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12515" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[4];
  assign _06637_ = _06636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12516" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[5];
  assign _06638_ = _06637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12516" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[6];
  assign _06639_ = _06638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12517" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[7];
  assign _06640_ = _06639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12517" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[8];
  assign _06641_ = _06640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12518" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[9];
  assign _06642_ = _06641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12518" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[10];
  assign _06643_ = _06642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12519" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[11];
  assign _06644_ = _06643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12519" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[12];
  assign _06645_ = _06644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12520" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[13];
  assign _06646_ = _06645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12520" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[14];
  assign _06647_ = _06646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12521" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[15];
  assign _06648_ = _06647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12521" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[16];
  assign _06649_ = _06648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12522" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[17];
  assign _06650_ = _06649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12522" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[18];
  assign _06651_ = _06650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12523" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[19];
  assign _06652_ = _06651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12523" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[20];
  assign _06653_ = _06652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12524" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[21];
  assign _06654_ = _06653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12524" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[22];
  assign _06655_ = _06654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12525" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[23];
  assign _06656_ = _06655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12525" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[24];
  assign _06657_ = _06656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12526" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[25];
  assign _06658_ = _06657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12526" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[26];
  assign _06659_ = _06658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12527" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[27];
  assign _06660_ = _06659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12527" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[28];
  assign _06661_ = _06660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12528" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[29];
  assign _06662_ = _06661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12528" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[30];
  assign _06663_ = _06662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12529" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[31];
  assign _06664_ = _06663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12529" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[32];
  assign _06665_ = _06664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12530" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[33];
  assign _06666_ = _06665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12530" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[34];
  assign _06667_ = _06666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12531" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[35];
  assign _06668_ = _06667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12531" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[36];
  assign _06669_ = _06668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12532" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[37];
  assign _06670_ = _06669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12532" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[38];
  assign _06671_ = _06670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12533" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[39];
  assign _06672_ = _06671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12533" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[40];
  assign _06673_ = _06672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12534" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[41];
  assign _06674_ = _06673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12534" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[42];
  assign _06675_ = _06674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12535" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[43];
  assign _06676_ = _06675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12535" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[44];
  assign _06677_ = _06676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12536" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[45];
  assign _06678_ = _06677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12536" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[46];
  assign _06679_ = _06678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12537" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[47];
  assign _06680_ = _06679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12537" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[48];
  assign _06681_ = _06680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12538" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[49];
  assign _06682_ = _06681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12538" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[50];
  assign _06683_ = _06682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12539" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[51];
  assign _06684_ = _06683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12539" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[52];
  assign _06685_ = _06684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12540" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[53];
  assign _06686_ = _06685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12540" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[54];
  assign _06687_ = _06686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12541" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[55];
  assign _06688_ = _06687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12541" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[56];
  assign _06689_ = _06688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12542" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[57];
  assign _06690_ = _06689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12542" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[58];
  assign _06691_ = _06690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12543" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[59];
  assign _06692_ = _06691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12543" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[60];
  assign _06693_ = _06692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12544" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[61];
  assign _06694_ = _06693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12544" *) _04431_;
  assign _05324_ = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12551" *) _04433_;
  assign _06695_ = IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12554" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[1];
  assign _06696_ = _06695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12554" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[2];
  assign _06697_ = _06696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12555" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[3];
  assign _06698_ = _06697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12555" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[4];
  assign _06699_ = _06698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12556" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[5];
  assign _06700_ = _06699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12556" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[6];
  assign _06701_ = _06700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12557" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[7];
  assign _06702_ = _06701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12557" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[8];
  assign _06703_ = _06702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12558" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[9];
  assign _06704_ = _06703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12558" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[10];
  assign _06705_ = _06704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12559" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[11];
  assign _06706_ = _06705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12559" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[12];
  assign _06707_ = _06706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12560" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[13];
  assign _06708_ = _06707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12560" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[14];
  assign _06709_ = _06708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12561" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[15];
  assign _06710_ = _06709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12561" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[16];
  assign _06711_ = _06710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12562" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[17];
  assign _06712_ = _06711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12562" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[18];
  assign _06713_ = _06712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12563" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[19];
  assign _06714_ = _06713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12563" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[20];
  assign _06715_ = _06714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12564" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[21];
  assign _06716_ = _06715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12564" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[22];
  assign _06717_ = _06716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12565" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[23];
  assign _06718_ = _06717_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12565" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[24];
  assign _06719_ = _06718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12566" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[25];
  assign _06720_ = _06719_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12566" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[26];
  assign _06721_ = _06720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12567" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[27];
  assign _06722_ = _06721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12567" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[28];
  assign _06723_ = _06722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12568" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[29];
  assign _06724_ = _06723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12568" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[30];
  assign _06725_ = _06724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12569" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[31];
  assign _06726_ = _06725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12569" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[32];
  assign _06727_ = _06726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12570" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[33];
  assign _06728_ = _06727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12570" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[34];
  assign _06729_ = _06728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12571" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[35];
  assign _06730_ = _06729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12571" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[36];
  assign _06731_ = _06730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12572" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[37];
  assign _06732_ = _06731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12572" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[38];
  assign _06733_ = _06732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12573" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[39];
  assign _06734_ = _06733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12573" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[40];
  assign _06735_ = _06734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12574" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[41];
  assign _06736_ = _06735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12574" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[42];
  assign _06737_ = _06736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12575" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[43];
  assign _06738_ = _06737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12575" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[44];
  assign _06739_ = _06738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12576" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[45];
  assign _06740_ = _06739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12576" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[46];
  assign _06741_ = _06740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12577" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[47];
  assign _06742_ = _06741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12577" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[48];
  assign _06743_ = _06742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12578" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[49];
  assign _06744_ = _06743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12578" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[50];
  assign _06745_ = _06744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12579" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[51];
  assign _06746_ = _06745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12579" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[52];
  assign _06747_ = _06746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12580" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[53];
  assign _06748_ = _06747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12580" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[54];
  assign _06749_ = _06748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12581" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[55];
  assign _06750_ = _06749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12581" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[56];
  assign _06751_ = _06750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12582" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[57];
  assign _06752_ = _06751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12582" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[58];
  assign _06753_ = _06752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12583" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[59];
  assign _06754_ = _06753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12583" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[60];
  assign _06755_ = _06754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12584" *) IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[61];
  assign _06756_ = _06755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12584" *) _04434_;
  assign _05318_ = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12591" *) _04436_;
  assign _06757_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12594" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[1];
  assign _06758_ = _06757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12594" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[2];
  assign _06759_ = _06758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12595" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[3];
  assign _06760_ = _06759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12595" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[4];
  assign _06761_ = _06760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12596" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[5];
  assign _06762_ = _06761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12596" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[6];
  assign _06763_ = _06762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12597" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[7];
  assign _06764_ = _06763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12597" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[8];
  assign _06765_ = _06764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12598" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[9];
  assign _06766_ = _06765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12598" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[10];
  assign _06767_ = _06766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12599" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[11];
  assign _06768_ = _06767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12599" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[12];
  assign _06769_ = _06768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12600" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[13];
  assign _06770_ = _06769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12600" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[14];
  assign _06771_ = _06770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12601" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[15];
  assign _06772_ = _06771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12601" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[16];
  assign _06773_ = _06772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12602" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[17];
  assign _06774_ = _06773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12602" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[18];
  assign _06775_ = _06774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12603" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[19];
  assign _06776_ = _06775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12603" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[20];
  assign _06777_ = _06776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12604" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[21];
  assign _06778_ = _06777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12604" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[22];
  assign _06779_ = _06778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12605" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[23];
  assign _06780_ = _06779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12605" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[24];
  assign _06781_ = _06780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12606" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[25];
  assign _06782_ = _06781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12606" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[26];
  assign _06783_ = _06782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12607" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[27];
  assign _06784_ = _06783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12607" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[28];
  assign _06785_ = _06784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12608" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[29];
  assign _06786_ = _06785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12608" *) _04437_;
  assign _06787_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12615" *) _04439_;
  assign _06788_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12622" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[1];
  assign _06789_ = _06788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12622" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[2];
  assign _06790_ = _06789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12623" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[3];
  assign _06791_ = _06790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12623" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[4];
  assign _06792_ = _06791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12624" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[5];
  assign _06793_ = _06792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12624" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[6];
  assign _06794_ = _06793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12625" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[7];
  assign _06795_ = _06794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12625" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[8];
  assign _06796_ = _06795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12626" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[9];
  assign _06797_ = _06796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12626" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[10];
  assign _06798_ = _06797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12627" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[11];
  assign _06799_ = _06798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12627" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[12];
  assign _06800_ = _06799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12628" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[13];
  assign _06801_ = _06800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12628" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[14];
  assign _06802_ = _06801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12629" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[15];
  assign _06803_ = _06802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12629" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[16];
  assign _06804_ = _06803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12630" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[17];
  assign _06805_ = _06804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12630" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[18];
  assign _06806_ = _06805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12631" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[19];
  assign _06807_ = _06806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12631" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[20];
  assign _06808_ = _06807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12632" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[21];
  assign _06809_ = _06808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12632" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[22];
  assign _06810_ = _06809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12633" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[23];
  assign _06811_ = _06810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12633" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[24];
  assign _06812_ = _06811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12634" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[25];
  assign _06813_ = _06812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12634" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[26];
  assign _06814_ = _06813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12635" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[27];
  assign _06815_ = _06814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12635" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[28];
  assign _06816_ = _06815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12636" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[29];
  assign _06817_ = _06816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12636" *) _04440_;
  assign _06818_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12643" *) _04442_;
  assign _06819_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12650" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[1];
  assign _06820_ = _06819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12650" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[2];
  assign _06821_ = _06820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12651" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[3];
  assign _06822_ = _06821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12651" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[4];
  assign _06823_ = _06822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12652" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[5];
  assign _06824_ = _06823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12652" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[6];
  assign _06825_ = _06824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12653" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[7];
  assign _06826_ = _06825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12653" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[8];
  assign _06827_ = _06826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12654" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[9];
  assign _06828_ = _06827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12654" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[10];
  assign _06829_ = _06828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12655" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[11];
  assign _06830_ = _06829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12655" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[12];
  assign _06831_ = _06830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12656" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[13];
  assign _06832_ = _06831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12656" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[14];
  assign _06833_ = _06832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12657" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[15];
  assign _06834_ = _06833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12657" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[16];
  assign _06835_ = _06834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12658" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[17];
  assign _06836_ = _06835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12658" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[18];
  assign _06837_ = _06836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12659" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[19];
  assign _06838_ = _06837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12659" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[20];
  assign _06839_ = _06838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12660" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[21];
  assign _06840_ = _06839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12660" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[22];
  assign _06841_ = _06840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12661" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[23];
  assign _06842_ = _06841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12661" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[24];
  assign _06843_ = _06842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12662" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[25];
  assign _06844_ = _06843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12662" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[26];
  assign _06845_ = _06844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12663" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[27];
  assign _06846_ = _06845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12663" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[28];
  assign _06847_ = _06846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12664" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[29];
  assign _06848_ = _06847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12664" *) _04443_;
  assign _06849_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12671" *) _04445_;
  assign _06850_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12678" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[1];
  assign _06851_ = _06850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12678" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[2];
  assign _06852_ = _06851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12679" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[3];
  assign _06853_ = _06852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12679" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[4];
  assign _06854_ = _06853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12680" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[5];
  assign _06855_ = _06854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12680" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[6];
  assign _06856_ = _06855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12681" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[7];
  assign _06857_ = _06856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12681" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[8];
  assign _06858_ = _06857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12682" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[9];
  assign _06859_ = _06858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12682" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[10];
  assign _06860_ = _06859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12683" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[11];
  assign _06861_ = _06860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12683" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[12];
  assign _06862_ = _06861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12684" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[13];
  assign _06863_ = _06862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12684" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[14];
  assign _06864_ = _06863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12685" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[15];
  assign _06865_ = _06864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12685" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[16];
  assign _06866_ = _06865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12686" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[17];
  assign _06867_ = _06866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12686" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[18];
  assign _06868_ = _06867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12687" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[19];
  assign _06869_ = _06868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12687" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[20];
  assign _06870_ = _06869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12688" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[21];
  assign _06871_ = _06870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12688" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[22];
  assign _06872_ = _06871_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12689" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[23];
  assign _06873_ = _06872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12689" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[24];
  assign _06874_ = _06873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12690" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[25];
  assign _06875_ = _06874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12690" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[26];
  assign _06876_ = _06875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12691" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[27];
  assign _06877_ = _06876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12691" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[28];
  assign _06878_ = _06877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12692" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[29];
  assign _06879_ = _06878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12692" *) _04446_;
  assign _06880_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12699" *) _04448_;
  assign _06881_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12706" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[1];
  assign _06882_ = _06881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12706" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[2];
  assign _06883_ = _06882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12707" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[3];
  assign _06884_ = _06883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12707" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[4];
  assign _06885_ = _06884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12708" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[5];
  assign _06886_ = _06885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12708" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[6];
  assign _06887_ = _06886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12709" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[7];
  assign _06888_ = _06887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12709" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[8];
  assign _06889_ = _06888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12710" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[9];
  assign _06890_ = _06889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12710" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[10];
  assign _06891_ = _06890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12711" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[11];
  assign _06892_ = _06891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12711" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[12];
  assign _06893_ = _06892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12712" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[13];
  assign _06894_ = _06893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12712" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[14];
  assign _06895_ = _06894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12713" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[15];
  assign _06896_ = _06895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12713" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[16];
  assign _06897_ = _06896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12714" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[17];
  assign _06898_ = _06897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12714" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[18];
  assign _06899_ = _06898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12715" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[19];
  assign _06900_ = _06899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12715" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[20];
  assign _06901_ = _06900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12716" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[21];
  assign _06902_ = _06901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12716" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[22];
  assign _06903_ = _06902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12717" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[23];
  assign _06904_ = _06903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12717" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[24];
  assign _06905_ = _06904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12718" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[25];
  assign _06906_ = _06905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12718" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[26];
  assign _06907_ = _06906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12719" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[27];
  assign _06908_ = _06907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12719" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[28];
  assign _06909_ = _06908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12720" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[29];
  assign _06910_ = _06909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12720" *) _04449_;
  assign _06911_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12727" *) _04451_;
  assign _06912_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12734" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[1];
  assign _06913_ = _06912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12734" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[2];
  assign _06914_ = _06913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12735" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[3];
  assign _06915_ = _06914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12735" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[4];
  assign _06916_ = _06915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12736" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[5];
  assign _06917_ = _06916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12736" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[6];
  assign _06918_ = _06917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12737" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[7];
  assign _06919_ = _06918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12737" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[8];
  assign _06920_ = _06919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12738" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[9];
  assign _06921_ = _06920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12738" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[10];
  assign _06922_ = _06921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12739" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[11];
  assign _06923_ = _06922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12739" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[12];
  assign _06924_ = _06923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12740" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[13];
  assign _06925_ = _06924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12740" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[14];
  assign _06926_ = _06925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12741" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[15];
  assign _06927_ = _06926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12741" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[16];
  assign _06928_ = _06927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12742" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[17];
  assign _06929_ = _06928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12742" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[18];
  assign _06930_ = _06929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12743" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[19];
  assign _06931_ = _06930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12743" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[20];
  assign _06932_ = _06931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12744" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[21];
  assign _06933_ = _06932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12744" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[22];
  assign _06934_ = _06933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12745" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[23];
  assign _06935_ = _06934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12745" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[24];
  assign _06936_ = _06935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12746" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[25];
  assign _06937_ = _06936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12746" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[26];
  assign _06938_ = _06937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12747" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[27];
  assign _06939_ = _06938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12747" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[28];
  assign _06940_ = _06939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12748" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[29];
  assign _06941_ = _06940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12748" *) _04452_;
  assign _06942_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12755" *) _04454_;
  assign _06943_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12762" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[1];
  assign _06944_ = _06943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12762" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[2];
  assign _06945_ = _06944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12763" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[3];
  assign _06946_ = _06945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12763" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[4];
  assign _06947_ = _06946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12764" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[5];
  assign _06948_ = _06947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12764" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[6];
  assign _06949_ = _06948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12765" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[7];
  assign _06950_ = _06949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12765" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[8];
  assign _06951_ = _06950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12766" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[9];
  assign _06952_ = _06951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12766" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[10];
  assign _06953_ = _06952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12767" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[11];
  assign _06954_ = _06953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12767" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[12];
  assign _06955_ = _06954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12768" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[13];
  assign _06956_ = _06955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12768" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[14];
  assign _06957_ = _06956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12769" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[15];
  assign _06958_ = _06957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12769" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[16];
  assign _06959_ = _06958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12770" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[17];
  assign _06960_ = _06959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12770" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[18];
  assign _06961_ = _06960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12771" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[19];
  assign _06962_ = _06961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12771" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[20];
  assign _06963_ = _06962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12772" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[21];
  assign _06964_ = _06963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12772" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[22];
  assign _06965_ = _06964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12773" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[23];
  assign _06966_ = _06965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12773" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[24];
  assign _06967_ = _06966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12774" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[25];
  assign _06968_ = _06967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12774" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[26];
  assign _06969_ = _06968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12775" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[27];
  assign _06970_ = _06969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12775" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[28];
  assign _06971_ = _06970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12776" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[29];
  assign _06972_ = _06971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12776" *) _04455_;
  assign _06973_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12783" *) _04457_;
  assign _06974_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12790" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[1];
  assign _06975_ = _06974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12790" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[2];
  assign _06976_ = _06975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12791" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[3];
  assign _06977_ = _06976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12791" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[4];
  assign _06978_ = _06977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12792" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[5];
  assign _06979_ = _06978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12792" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[6];
  assign _06980_ = _06979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12793" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[7];
  assign _06981_ = _06980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12793" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[8];
  assign _06982_ = _06981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12794" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[9];
  assign _06983_ = _06982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12794" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[10];
  assign _06984_ = _06983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12795" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[11];
  assign _06985_ = _06984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12795" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[12];
  assign _06986_ = _06985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12796" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[13];
  assign _06987_ = _06986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12796" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[14];
  assign _06988_ = _06987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12797" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[15];
  assign _06989_ = _06988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12797" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[16];
  assign _06990_ = _06989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12798" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[17];
  assign _06991_ = _06990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12798" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[18];
  assign _06992_ = _06991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12799" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[19];
  assign _06993_ = _06992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12799" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[20];
  assign _06994_ = _06993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12800" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[21];
  assign _06995_ = _06994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12800" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[22];
  assign _06996_ = _06995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12801" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[23];
  assign _06997_ = _06996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12801" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[24];
  assign _06998_ = _06997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12802" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[25];
  assign _06999_ = _06998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12802" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[26];
  assign _07000_ = _06999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12803" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[27];
  assign _07001_ = _07000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12803" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[28];
  assign _07002_ = _07001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12804" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[29];
  assign _07003_ = _07002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12804" *) _04458_;
  assign _07004_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12811" *) _04460_;
  assign _07005_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12818" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[1];
  assign _07006_ = _07005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12818" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[2];
  assign _07007_ = _07006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12819" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[3];
  assign _07008_ = _07007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12819" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[4];
  assign _07009_ = _07008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12820" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[5];
  assign _07010_ = _07009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12820" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[6];
  assign _07011_ = _07010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12821" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[7];
  assign _07012_ = _07011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12821" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[8];
  assign _07013_ = _07012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12822" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[9];
  assign _07014_ = _07013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12822" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[10];
  assign _07015_ = _07014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12823" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[11];
  assign _07016_ = _07015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12823" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[12];
  assign _07017_ = _07016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12824" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[13];
  assign _07018_ = _07017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12824" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[14];
  assign _07019_ = _07018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12825" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[15];
  assign _07020_ = _07019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12825" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[16];
  assign _07021_ = _07020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12826" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[17];
  assign _07022_ = _07021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12826" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[18];
  assign _07023_ = _07022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12827" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[19];
  assign _07024_ = _07023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12827" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[20];
  assign _07025_ = _07024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12828" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[21];
  assign _07026_ = _07025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12828" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[22];
  assign _07027_ = _07026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12829" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[23];
  assign _07028_ = _07027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12829" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[24];
  assign _07029_ = _07028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12830" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[25];
  assign _07030_ = _07029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12830" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[26];
  assign _07031_ = _07030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12831" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[27];
  assign _07032_ = _07031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12831" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[28];
  assign _07033_ = _07032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12832" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[29];
  assign _07034_ = _07033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12832" *) _04461_;
  assign _07035_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12839" *) _04463_;
  assign _07036_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12846" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[1];
  assign _07037_ = _07036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12846" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[2];
  assign _07038_ = _07037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12847" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[3];
  assign _07039_ = _07038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12847" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[4];
  assign _07040_ = _07039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12848" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[5];
  assign _07041_ = _07040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12848" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[6];
  assign _07042_ = _07041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12849" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[7];
  assign _07043_ = _07042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12849" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[8];
  assign _07044_ = _07043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12850" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[9];
  assign _07045_ = _07044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12850" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[10];
  assign _07046_ = _07045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12851" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[11];
  assign _07047_ = _07046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12851" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[12];
  assign _07048_ = _07047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12852" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[13];
  assign _07049_ = _07048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12852" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[14];
  assign _07050_ = _07049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12853" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[15];
  assign _07051_ = _07050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12853" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[16];
  assign _07052_ = _07051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12854" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[17];
  assign _07053_ = _07052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12854" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[18];
  assign _07054_ = _07053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12855" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[19];
  assign _07055_ = _07054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12855" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[20];
  assign _07056_ = _07055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12856" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[21];
  assign _07057_ = _07056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12856" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[22];
  assign _07058_ = _07057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12857" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[23];
  assign _07059_ = _07058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12857" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[24];
  assign _07060_ = _07059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12858" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[25];
  assign _07061_ = _07060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12858" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[26];
  assign _07062_ = _07061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12859" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[27];
  assign _07063_ = _07062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12859" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[28];
  assign _07064_ = _07063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12860" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[29];
  assign _07065_ = _07064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12860" *) _04464_;
  assign _07066_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12867" *) _04466_;
  assign _07067_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12874" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[1];
  assign _07068_ = _07067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12874" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[2];
  assign _07069_ = _07068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12875" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[3];
  assign _07070_ = _07069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12875" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[4];
  assign _07071_ = _07070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12876" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[5];
  assign _07072_ = _07071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12876" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[6];
  assign _07073_ = _07072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12877" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[7];
  assign _07074_ = _07073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12877" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[8];
  assign _07075_ = _07074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12878" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[9];
  assign _07076_ = _07075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12878" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[10];
  assign _07077_ = _07076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12879" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[11];
  assign _07078_ = _07077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12879" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[12];
  assign _07079_ = _07078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12880" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[13];
  assign _07080_ = _07079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12880" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[14];
  assign _07081_ = _07080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12881" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[15];
  assign _07082_ = _07081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12881" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[16];
  assign _07083_ = _07082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12882" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[17];
  assign _07084_ = _07083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12882" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[18];
  assign _07085_ = _07084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12883" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[19];
  assign _07086_ = _07085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12883" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[20];
  assign _07087_ = _07086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12884" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[21];
  assign _07088_ = _07087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12884" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[22];
  assign _07089_ = _07088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12885" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[23];
  assign _07090_ = _07089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12885" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[24];
  assign _07091_ = _07090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12886" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[25];
  assign _07092_ = _07091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12886" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[26];
  assign _07093_ = _07092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12887" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[27];
  assign _07094_ = _07093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12887" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[28];
  assign _07095_ = _07094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12888" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[29];
  assign _07096_ = _07095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12888" *) _04467_;
  assign _07097_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12895" *) _04469_;
  assign _07098_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12902" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[1];
  assign _07099_ = _07098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12902" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[2];
  assign _07100_ = _07099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12903" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[3];
  assign _07101_ = _07100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12903" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[4];
  assign _07102_ = _07101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12904" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[5];
  assign _07103_ = _07102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12904" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[6];
  assign _07104_ = _07103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12905" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[7];
  assign _07105_ = _07104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12905" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[8];
  assign _07106_ = _07105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12906" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[9];
  assign _07107_ = _07106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12906" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[10];
  assign _07108_ = _07107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12907" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[11];
  assign _07109_ = _07108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12907" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[12];
  assign _07110_ = _07109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12908" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[13];
  assign _07111_ = _07110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12908" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[14];
  assign _07112_ = _07111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12909" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[15];
  assign _07113_ = _07112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12909" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[16];
  assign _07114_ = _07113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12910" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[17];
  assign _07115_ = _07114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12910" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[18];
  assign _07116_ = _07115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12911" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[19];
  assign _07117_ = _07116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12911" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[20];
  assign _07118_ = _07117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12912" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[21];
  assign _07119_ = _07118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12912" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[22];
  assign _07120_ = _07119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12913" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[23];
  assign _07121_ = _07120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12913" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[24];
  assign _07122_ = _07121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12914" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[25];
  assign _07123_ = _07122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12914" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[26];
  assign _07124_ = _07123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12915" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[27];
  assign _07125_ = _07124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12915" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[28];
  assign _07126_ = _07125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12916" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[29];
  assign _07127_ = _07126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12916" *) _04470_;
  assign _07128_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12923" *) _04472_;
  assign _07129_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12930" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[1];
  assign _07130_ = _07129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12930" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[2];
  assign _07131_ = _07130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12931" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[3];
  assign _07132_ = _07131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12931" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[4];
  assign _07133_ = _07132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12932" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[5];
  assign _07134_ = _07133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12932" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[6];
  assign _07135_ = _07134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12933" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[7];
  assign _07136_ = _07135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12933" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[8];
  assign _07137_ = _07136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12934" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[9];
  assign _07138_ = _07137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12934" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[10];
  assign _07139_ = _07138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12935" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[11];
  assign _07140_ = _07139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12935" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[12];
  assign _07141_ = _07140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12936" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[13];
  assign _07142_ = _07141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12936" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[14];
  assign _07143_ = _07142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12937" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[15];
  assign _07144_ = _07143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12937" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[16];
  assign _07145_ = _07144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12938" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[17];
  assign _07146_ = _07145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12938" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[18];
  assign _07147_ = _07146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12939" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[19];
  assign _07148_ = _07147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12939" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[20];
  assign _07149_ = _07148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12940" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[21];
  assign _07150_ = _07149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12940" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[22];
  assign _07151_ = _07150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12941" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[23];
  assign _07152_ = _07151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12941" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[24];
  assign _07153_ = _07152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12942" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[25];
  assign _07154_ = _07153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12942" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[26];
  assign _07155_ = _07154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12943" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[27];
  assign _07156_ = _07155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12943" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[28];
  assign _07157_ = _07156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12944" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[29];
  assign _07158_ = _07157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12944" *) _04473_;
  assign _07159_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12951" *) _04475_;
  assign _07160_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12958" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[1];
  assign _07161_ = _07160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12958" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[2];
  assign _07162_ = _07161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12959" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[3];
  assign _07163_ = _07162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12959" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[4];
  assign _07164_ = _07163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12960" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[5];
  assign _07165_ = _07164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12960" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[6];
  assign _07166_ = _07165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12961" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[7];
  assign _07167_ = _07166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12961" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[8];
  assign _07168_ = _07167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12962" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[9];
  assign _07169_ = _07168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12962" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[10];
  assign _07170_ = _07169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12963" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[11];
  assign _07171_ = _07170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12963" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[12];
  assign _07172_ = _07171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12964" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[13];
  assign _07173_ = _07172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12964" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[14];
  assign _07174_ = _07173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12965" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[15];
  assign _07175_ = _07174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12965" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[16];
  assign _07176_ = _07175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12966" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[17];
  assign _07177_ = _07176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12966" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[18];
  assign _07178_ = _07177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12967" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[19];
  assign _07179_ = _07178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12967" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[20];
  assign _07180_ = _07179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12968" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[21];
  assign _07181_ = _07180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12968" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[22];
  assign _07182_ = _07181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12969" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[23];
  assign _07183_ = _07182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12969" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[24];
  assign _07184_ = _07183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12970" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[25];
  assign _07185_ = _07184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12970" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[26];
  assign _07186_ = _07185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12971" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[27];
  assign _07187_ = _07186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12971" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[28];
  assign _07188_ = _07187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12972" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[29];
  assign _07189_ = _07188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12972" *) _04476_;
  assign _07190_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12979" *) _04478_;
  assign _07191_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12986" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[1];
  assign _07192_ = _07191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12986" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[2];
  assign _07193_ = _07192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12987" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[3];
  assign _07194_ = _07193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12987" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[4];
  assign _07195_ = _07194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12988" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[5];
  assign _07196_ = _07195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12988" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[6];
  assign _07197_ = _07196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12989" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[7];
  assign _07198_ = _07197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12989" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[8];
  assign _07199_ = _07198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12990" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[9];
  assign _07200_ = _07199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12990" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[10];
  assign _07201_ = _07200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12991" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[11];
  assign _07202_ = _07201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12991" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[12];
  assign _07203_ = _07202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12992" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[13];
  assign _07204_ = _07203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12992" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[14];
  assign _07205_ = _07204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12993" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[15];
  assign _07206_ = _07205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12993" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[16];
  assign _07207_ = _07206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12994" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[17];
  assign _07208_ = _07207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12994" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[18];
  assign _07209_ = _07208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12995" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[19];
  assign _07210_ = _07209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12995" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[20];
  assign _07211_ = _07210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12996" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[21];
  assign _07212_ = _07211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12996" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[22];
  assign _07213_ = _07212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12997" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[23];
  assign _07214_ = _07213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12997" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[24];
  assign _07215_ = _07214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12998" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[25];
  assign _07216_ = _07215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12998" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[26];
  assign _07217_ = _07216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12999" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[27];
  assign _07218_ = _07217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:12999" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[28];
  assign _07219_ = _07218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13000" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[29];
  assign _07220_ = _07219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13000" *) _04479_;
  assign _07221_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13007" *) _04481_;
  assign _07222_ = IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13014" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[1];
  assign _07223_ = _07222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13014" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[2];
  assign _07224_ = _07223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13015" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[3];
  assign _07225_ = _07224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13015" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[4];
  assign _07226_ = _07225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13016" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[5];
  assign _07227_ = _07226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13016" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[6];
  assign _07228_ = _07227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13017" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[7];
  assign _07229_ = _07228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13017" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[8];
  assign _07230_ = _07229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13018" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[9];
  assign _07231_ = _07230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13018" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[10];
  assign _07232_ = _07231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13019" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[11];
  assign _07233_ = _07232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13019" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[12];
  assign _07234_ = _07233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13020" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[13];
  assign _07235_ = _07234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13020" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[14];
  assign _07236_ = _07235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13021" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[15];
  assign _07237_ = _07236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13021" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[16];
  assign _07238_ = _07237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13022" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[17];
  assign _07239_ = _07238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13022" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[18];
  assign _07240_ = _07239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13023" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[19];
  assign _07241_ = _07240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13023" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[20];
  assign _07242_ = _07241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13024" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[21];
  assign _07243_ = _07242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13024" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[22];
  assign _07244_ = _07243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13025" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[23];
  assign _07245_ = _07244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13025" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[24];
  assign _07246_ = _07245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13026" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[25];
  assign _07247_ = _07246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13026" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[26];
  assign _07248_ = _07247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13027" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[27];
  assign _07249_ = _07248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13027" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[28];
  assign _07250_ = _07249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13028" *) IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[29];
  assign _07251_ = _07250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13028" *) _04482_;
  assign _07252_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13035" *) _04484_;
  assign _07253_ = FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13047" *) FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[1];
  assign _07254_ = _07253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13047" *) FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[2];
  assign _07255_ = _07254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13048" *) FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[3];
  assign _07256_ = _07255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13048" *) FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[4];
  assign _07257_ = _07256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13048" *) FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[6];
  assign _07258_ = FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13056" *) FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[1];
  assign _07259_ = _07258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13056" *) FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[2];
  assign _07260_ = _07259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13057" *) FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[3];
  assign _07261_ = _07260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13057" *) FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[4];
  assign _07262_ = _07261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13057" *) FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[6];
  assign _07263_ = cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13065" *) cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[1];
  assign _07264_ = _07263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13065" *) cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[2];
  assign _07265_ = _07264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13066" *) cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[3];
  assign _07266_ = _07265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13066" *) cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[4];
  assign _07267_ = _07266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13066" *) cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[6];
  assign _07268_ = cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13074" *) cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1];
  assign _07269_ = _07268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13074" *) cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2];
  assign _07270_ = _07269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13075" *) cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3];
  assign _07271_ = _07270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13075" *) cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4];
  assign _07272_ = _07271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13075" *) cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6];
  assign _07273_ = cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13083" *) cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[1];
  assign _07274_ = _07273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13083" *) cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[2];
  assign _07275_ = _07274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13084" *) cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[3];
  assign _07276_ = _07275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13084" *) cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[4];
  assign _07277_ = _07276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13084" *) cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[6];
  assign _07278_ = cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13092" *) cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1];
  assign _07279_ = _07278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13092" *) cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2];
  assign _07280_ = _07279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13093" *) cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3];
  assign _07281_ = _07280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13093" *) cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4];
  assign _07282_ = _07281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13093" *) cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6];
  assign _07283_ = cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13101" *) cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1];
  assign _07284_ = _07283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13101" *) cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2];
  assign _07285_ = _07284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13102" *) cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3];
  assign _07286_ = _07285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13102" *) cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4];
  assign _07287_ = _07286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13102" *) cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6];
  assign _07288_ = cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13110" *) cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1];
  assign _07289_ = _07288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13110" *) cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2];
  assign _07290_ = _07289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13111" *) cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3];
  assign _07291_ = _07290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13111" *) cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4];
  assign _07292_ = _07291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13111" *) cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6];
  assign _07293_ = FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13119" *) FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[1];
  assign _07294_ = _07293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13119" *) FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[2];
  assign _07295_ = _07294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13120" *) FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[3];
  assign _07296_ = _07295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13120" *) FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[4];
  assign _07297_ = _07296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13120" *) FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[6];
  assign _07298_ = cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13128" *) cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1];
  assign _07299_ = _07298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13128" *) cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2];
  assign _07300_ = _07299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13129" *) cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3];
  assign _07301_ = _07300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13129" *) cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4];
  assign _07302_ = _07301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13129" *) cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6];
  assign _07303_ = cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13137" *) cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1];
  assign _07304_ = _07303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13137" *) cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2];
  assign _07305_ = _07304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13138" *) cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3];
  assign _07306_ = _07305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13138" *) cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4];
  assign _07307_ = _07306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13138" *) cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6];
  assign _07308_ = cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13146" *) cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1];
  assign _07309_ = _07308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13146" *) cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2];
  assign _07310_ = _07309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13147" *) cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3];
  assign _07311_ = _07310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13147" *) cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4];
  assign _07312_ = _07311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13147" *) cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6];
  assign _07313_ = cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13155" *) cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1];
  assign _07314_ = _07313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13155" *) cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2];
  assign _07315_ = _07314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13156" *) cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3];
  assign _07316_ = _07315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13156" *) cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4];
  assign _07317_ = _07316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13156" *) cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6];
  assign _07318_ = cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13164" *) cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1];
  assign _07319_ = _07318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13164" *) cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2];
  assign _07320_ = _07319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13165" *) cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3];
  assign _07321_ = _07320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13165" *) cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4];
  assign _07322_ = _07321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13165" *) cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6];
  assign _07323_ = cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13173" *) cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1];
  assign _07324_ = _07323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13173" *) cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2];
  assign _07325_ = _07324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13174" *) cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3];
  assign _07326_ = _07325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13174" *) cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4];
  assign _07327_ = _07326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13174" *) cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6];
  assign _07328_ = cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13182" *) cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[1];
  assign _07329_ = _07328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13182" *) cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[2];
  assign _07330_ = _07329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13183" *) cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[3];
  assign _07331_ = _07330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13183" *) cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[4];
  assign _07332_ = _07331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13183" *) cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[6];
  assign _07333_ = cvt_1_IntSaturation_17U_8U_else_if_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13193" *) FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  assign _07334_ = cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13207" *) FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  assign _07335_ = cvt_else_equal_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13214" *) cvt_else_equal_tmp_1;
  assign _07336_ = _07335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13214" *) and_2136_cse;
  assign _07337_ = cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13225" *) FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  assign _07338_ = cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13238" *) FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  assign _07339_ = cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13252" *) FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  assign _07340_ = cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13266" *) FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  assign _07341_ = cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13280" *) FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  assign _07342_ = cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13294" *) FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  assign _07343_ = cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13308" *) FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  assign _07344_ = cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13322" *) FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  assign _07345_ = cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13336" *) FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  assign _07346_ = cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13350" *) FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  assign _07347_ = cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13364" *) FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  assign _07348_ = cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13373" *) cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1;
  assign _07349_ = cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13387" *) FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  assign _07350_ = cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13401" *) FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  assign _07351_ = _04102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13528" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[23];
  assign _07352_ = _04103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13530" *) _04104_;
  assign _07353_ = _07352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13530" *) FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva[23];
  assign _07354_ = _04105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13544" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[23];
  assign _07355_ = _04106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13546" *) _04107_;
  assign _07356_ = _07355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13546" *) FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva[23];
  assign _07357_ = _04108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13560" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[23];
  assign _07358_ = _04109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13562" *) _04110_;
  assign _07359_ = _07358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13562" *) FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva[23];
  assign _07360_ = _04111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13576" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva[23];
  assign _07361_ = _04112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13578" *) _04113_;
  assign _07362_ = _07361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13578" *) FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva[23];
  assign _07363_ = _04114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13592" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva[23];
  assign _07364_ = _04115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13594" *) _04116_;
  assign _07365_ = _07364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13594" *) FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva[23];
  assign _07366_ = _04117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13608" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva[23];
  assign _07367_ = _04118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13610" *) _04119_;
  assign _07368_ = _07367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13610" *) FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva[23];
  assign _07369_ = _04120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13624" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva[23];
  assign _07370_ = _04121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13626" *) _04122_;
  assign _07371_ = _07370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13626" *) FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva[23];
  assign _07372_ = _04123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13640" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva[23];
  assign _07373_ = _04124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13642" *) _04125_;
  assign _07374_ = _07373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13642" *) FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva[23];
  assign _07375_ = _04126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13656" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva[23];
  assign _07376_ = _04127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13658" *) _04128_;
  assign _07377_ = _07376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13658" *) FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva[23];
  assign _07378_ = _04129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13672" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva[23];
  assign _07379_ = _04130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13674" *) _04131_;
  assign _07380_ = _07379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13674" *) FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva[23];
  assign _07381_ = _04132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13688" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva[23];
  assign _07382_ = _04133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13690" *) _04134_;
  assign _07383_ = _07382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13690" *) FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva[23];
  assign _07384_ = _04135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13704" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva[23];
  assign _07385_ = _04136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13706" *) _04137_;
  assign _07386_ = _07385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13706" *) FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva[23];
  assign _07387_ = _04138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13720" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva[23];
  assign _07388_ = _04139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13722" *) _04140_;
  assign _07389_ = _07388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13722" *) FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva[23];
  assign _07390_ = _04141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13736" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva[23];
  assign _07391_ = _04142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13738" *) _04143_;
  assign _07392_ = _07391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13738" *) FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva[23];
  assign _07393_ = _04144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13752" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva[23];
  assign _07394_ = _04145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13754" *) _04146_;
  assign _07395_ = _07394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13754" *) FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva[23];
  assign _07396_ = _04147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13768" *) FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[23];
  assign _07397_ = _04148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13770" *) _04149_;
  assign _07398_ = _07397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13770" *) FpMantDecShiftRight_23U_8U_10U_least_mask_sva[23];
  assign _04385_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13786" *) nand_133_cse;
  assign _04382_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13794" *) nand_135_cse;
  assign _04379_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13802" *) nand_137_cse;
  assign _04376_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13810" *) nand_139_cse;
  assign _04373_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13818" *) nand_141_cse;
  assign _04370_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13826" *) nand_143_cse;
  assign _04367_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13834" *) nand_145_cse;
  assign _04364_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13842" *) nand_147_cse;
  assign _04361_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13850" *) nand_149_cse;
  assign _04358_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13858" *) nand_151_cse;
  assign _04355_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13866" *) nand_153_cse;
  assign _04352_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13874" *) nand_156_cse;
  assign _04349_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13882" *) nand_158_cse;
  assign _04346_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13890" *) nand_160_cse;
  assign _04343_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13898" *) nand_162_cse;
  assign _04340_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13906" *) nand_164_cse;
  assign _07399_ = cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13976" *) IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0;
  assign _07400_ = cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13978" *) IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0;
  assign _07401_ = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13980" *) IsNaN_5U_10U_land_3_lpi_1_dfm_4;
  assign _07402_ = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13982" *) IsNaN_5U_10U_land_4_lpi_1_dfm_4;
  assign _07403_ = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13984" *) IsNaN_5U_10U_land_5_lpi_1_dfm_4;
  assign _07404_ = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13986" *) IsNaN_5U_10U_land_6_lpi_1_dfm_4;
  assign _07405_ = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13988" *) IsNaN_5U_10U_land_7_lpi_1_dfm_5;
  assign _07406_ = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13990" *) IsNaN_5U_10U_land_8_lpi_1_dfm_4;
  assign _07407_ = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13992" *) IsNaN_5U_10U_land_9_lpi_1_dfm_4;
  assign _07408_ = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13994" *) IsNaN_5U_10U_land_10_lpi_1_dfm_4;
  assign _07409_ = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13996" *) IsNaN_5U_10U_land_11_lpi_1_dfm_4;
  assign _07410_ = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:13998" *) IsNaN_5U_10U_land_12_lpi_1_dfm_4;
  assign _07411_ = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14000" *) IsNaN_5U_10U_land_13_lpi_1_dfm_4;
  assign _07412_ = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14002" *) IsNaN_5U_10U_land_14_lpi_1_dfm_5;
  assign _07413_ = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14004" *) IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0;
  assign _07414_ = cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14006" *) IsNaN_5U_10U_land_lpi_1_dfm_4;
  assign _07415_ = cvt_if_unequal_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14071" *) cfg_mode_eql_1_sva_6;
  assign _07416_ = _07415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14071" *) cvt_unequal_tmp_21;
  assign or_tmp_19 = cfg_proc_precision_rsci_d[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14107" *) _04567_;
  assign or_23_nl = _04185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14108" *) or_4550_cse;
  assign _07417_ = nor_2040_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14110" *) cfg_proc_precision_rsci_d[0];
  assign or_tmp_24 = _07417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14110" *) _04567_;
  assign _07418_ = _04568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14113" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2;
  assign _07419_ = _07418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14113" *) _04185_;
  assign or_86_nl = _07419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14113" *) or_4550_cse;
  assign _07420_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14121" *) _04569_;
  assign or_tmp_213 = or_2242_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14124" *) _00065_;
  assign _07421_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14125" *) and_dcpl_3;
  assign or_tmp_218 = cfg_out_precision_1_sva_st_154[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14128" *) not_tmp_119;
  assign _07422_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14131" *) _04570_;
  assign _07423_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14134" *) _04188_;
  assign _07424_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14136" *) _04571_;
  assign _07425_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14139" *) _04572_;
  assign or_tmp_306 = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14142" *) or_4862_cse;
  assign _07426_ = cfg_proc_precision_1_sva_st_64[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14143" *) _04573_;
  assign or_378_nl = _04185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14146" *) cfg_mode_eql_1_sva_4;
  assign or_tmp_378 = _05427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14150" *) or_4862_cse;
  assign _07427_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14151" *) _00058_;
  assign _07428_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14153" *) _04575_;
  assign or_tmp_389 = cfg_proc_precision_1_sva_st_89[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14156" *) _04576_;
  assign _07429_ = cfg_proc_precision_1_sva_st_64[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14157" *) _04185_;
  assign _07430_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14159" *) _00058_;
  assign _07431_ = cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14162" *) or_2251_nl;
  assign or_429_nl = _07431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14162" *) _00066_;
  assign _07432_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14164" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign or_431_nl = _07432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14164" *) nor_50_cse;
  assign _07433_ = nor_2040_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14167" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp;
  assign _07434_ = _07433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14167" *) or_2251_nl;
  assign or_434_nl = _07434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14167" *) _00066_;
  assign _07435_ = IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14171" *) cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  assign or_448_nl = cfg_proc_precision_1_sva_st_64[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14174" *) _04577_;
  assign or_445_nl = _01547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14180" *) cfg_out_precision_1_sva_st_154[0];
  assign _07436_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14184" *) _04578_;
  assign _07437_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14186" *) _04579_;
  assign _07438_ = _04185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *) or_2251_nl;
  assign _07439_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  assign or_2688_nl = _07439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14189" *) _04580_;
  assign _07440_ = nor_2219_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14190" *) _00058_;
  assign _07441_ = _07440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14191" *) or_578_cse;
  assign _07442_ = _07441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14191" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign or_2691_nl = _07442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14192" *) nor_50_cse;
  assign _07443_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14195" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  assign or_2696_nl = _07443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14195" *) _04580_;
  assign _07444_ = _07441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14197" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign or_2699_nl = _07444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14198" *) nor_50_cse;
  assign or_510_cse = IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14201" *) cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign _07445_ = _01549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14204" *) cfg_out_precision_1_sva_st_154[0];
  assign _07446_ = _07445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14204" *) _04581_;
  assign _07447_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14206" *) _04579_;
  assign or_520_nl = _01550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14210" *) cfg_out_precision_1_sva_st_149[0];
  assign _07448_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14212" *) _04581_;
  assign or_451_cse = _04582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14214" *) cfg_mode_eql_1_sva_5;
  assign or_423_cse = or_451_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14215" *) or_425_cse;
  assign or_tmp_533 = or_423_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14215" *) _00058_;
  assign _07449_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14225" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign or_2705_nl = _07449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14225" *) _04583_;
  assign _07450_ = nor_151_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14226" *) nor_2219_cse;
  assign _07451_ = _07450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14226" *) _00058_;
  assign _07452_ = _07451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14227" *) or_578_cse;
  assign _07453_ = _07452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14227" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign or_2709_nl = _07453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14227" *) nor_50_cse;
  assign _07454_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14229" *) _04584_;
  assign _07455_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14234" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  assign or_2714_nl = _07455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14234" *) _04580_;
  assign _07456_ = _07441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14236" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign or_2717_nl = _07456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14237" *) nor_50_cse;
  assign _07457_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14239" *) nor_151_cse;
  assign _07458_ = _01552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14242" *) cfg_out_precision_1_sva_st_154[0];
  assign _07459_ = _07458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14242" *) _04581_;
  assign or_600_cse = IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14244" *) cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign or_599_nl = _01553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14247" *) cfg_out_precision_1_sva_st_149[0];
  assign _07460_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14252" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign or_2723_nl = _07460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14252" *) _04580_;
  assign _07461_ = _07452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14254" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign or_2727_nl = _07461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14254" *) nor_50_cse;
  assign _07462_ = _01554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14258" *) cfg_out_precision_1_sva_st_154[0];
  assign _07463_ = _07462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14258" *) _04581_;
  assign or_645_nl = _01555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14262" *) cfg_out_precision_1_sva_st_149[0];
  assign _07464_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14267" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign or_2733_nl = _07464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14267" *) _04580_;
  assign _07465_ = _07452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14269" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign or_2737_nl = _07465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14269" *) nor_50_cse;
  assign _07466_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14273" *) _04585_;
  assign _07467_ = _01556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14276" *) cfg_out_precision_1_sva_st_154[0];
  assign _07468_ = _07467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14276" *) _04581_;
  assign _07469_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14278" *) _04586_;
  assign or_690_nl = _01557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14282" *) cfg_out_precision_1_sva_st_149[0];
  assign _07470_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14284" *) _04587_;
  assign _07471_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14286" *) _04588_;
  assign _07472_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14288" *) _04589_;
  assign _07473_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14290" *) _04590_;
  assign _07474_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14293" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign or_2744_nl = _07474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14293" *) _04580_;
  assign _07475_ = _07452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14295" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign or_2749_nl = _07475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14295" *) nor_50_cse;
  assign _07476_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14299" *) nor_50_cse;
  assign _07477_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14303" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  assign or_2754_nl = _07477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14303" *) _04580_;
  assign _07478_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14305" *) or_578_cse;
  assign _07479_ = _07478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14305" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign or_2758_nl = _07479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14306" *) _04591_;
  assign _07480_ = _01560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14309" *) cfg_out_precision_1_sva_st_154[0];
  assign _07481_ = _07480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14309" *) _04581_;
  assign or_784_nl = _01561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14313" *) cfg_out_precision_1_sva_st_149[0];
  assign or_795_nl = _04592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14317" *) IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm;
  assign _07482_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14320" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign or_2764_nl = _07482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14321" *) _04583_;
  assign _07483_ = nor_151_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14322" *) _00058_;
  assign _07484_ = _07483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14323" *) or_578_cse;
  assign _07485_ = _07484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14323" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign or_2768_nl = _07485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14323" *) _04591_;
  assign _07486_ = _01562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14326" *) cfg_out_precision_1_sva_st_154[0];
  assign _07487_ = _07486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14326" *) _04581_;
  assign or_828_nl = _01563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14330" *) cfg_out_precision_1_sva_st_149[0];
  assign _07488_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14337" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign or_2774_nl = _07488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14338" *) _04583_;
  assign _07489_ = _07484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14340" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign or_2778_nl = _07489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14340" *) _04591_;
  assign _07490_ = _01564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14343" *) cfg_out_precision_1_sva_st_154[0];
  assign _07491_ = _07490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14343" *) _04588_;
  assign _07492_ = _01565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14347" *) cfg_out_precision_1_sva_st_149[0];
  assign or_871_nl = _04593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14347" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2;
  assign _07493_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14349" *) _04594_;
  assign _07494_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14354" *) _04595_;
  assign _07495_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14356" *) _04596_;
  assign _07496_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14358" *) _04597_;
  assign _07497_ = cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14361" *) or_2251_nl;
  assign or_894_nl = _07497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14361" *) _00064_;
  assign _07498_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14363" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign _07499_ = _07498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14363" *) cfg_out_precision_1_sva_st_149[0];
  assign or_898_nl = _07499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14364" *) _04598_;
  assign _07500_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14368" *) _04599_;
  assign _07501_ = cfg_proc_precision_1_sva_st_64[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14370" *) _04600_;
  assign _07502_ = _01567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14374" *) cfg_out_precision_1_sva_st_149[0];
  assign or_921_nl = _04601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14374" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2;
  assign _07503_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14376" *) _04602_;
  assign _07504_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14378" *) _04603_;
  assign _07505_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14382" *) _04604_;
  assign _07506_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14384" *) _04605_;
  assign _07507_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14387" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign or_2784_nl = _07507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14388" *) _04583_;
  assign _07508_ = _07478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14390" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign or_2789_nl = _07508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14390" *) _04606_;
  assign _07509_ = cfg_proc_precision_1_sva_st_64[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14392" *) _04607_;
  assign _07510_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14397" *) _04608_;
  assign _07511_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14399" *) _04609_;
  assign _07512_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14401" *) _04610_;
  assign _07513_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14404" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign or_2796_nl = _07513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14405" *) _04583_;
  assign _07514_ = _07478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14407" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign or_2802_nl = _07514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14407" *) _04611_;
  assign _07515_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14409" *) _00058_;
  assign _07516_ = _01568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14413" *) cfg_out_precision_1_sva_st_149[0];
  assign or_1015_nl = _04612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14413" *) IsNaN_5U_10U_nor_14_itm_2;
  assign _07517_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14415" *) _04613_;
  assign _07518_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14417" *) _04614_;
  assign _07519_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14419" *) _04615_;
  assign _07520_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14423" *) _04616_;
  assign _07521_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14425" *) _04617_;
  assign _07522_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14427" *) _04618_;
  assign _07523_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14430" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign or_2809_nl = _07523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14431" *) _04583_;
  assign _07524_ = _07478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14433" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign or_2815_nl = _07524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14433" *) _04611_;
  assign _07525_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14435" *) _04607_;
  assign _07526_ = cfg_proc_precision_1_sva_st_64[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14437" *) _04619_;
  assign _07527_ = _01569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14441" *) cfg_out_precision_1_sva_st_149[0];
  assign or_1072_nl = _04620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14441" *) IsNaN_5U_10U_nor_itm_2;
  assign _07528_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14443" *) _04621_;
  assign _07529_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14445" *) _04622_;
  assign _07530_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14447" *) _04623_;
  assign _07531_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14449" *) _04624_;
  assign _07532_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14453" *) _04625_;
  assign _07533_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14455" *) _04626_;
  assign _07534_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14457" *) _04627_;
  assign _07535_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14459" *) _04628_;
  assign _07536_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14462" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp;
  assign or_2823_nl = _07536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14463" *) _04580_;
  assign _07537_ = _07478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14465" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign or_2830_nl = _07537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14465" *) _04611_;
  assign _07538_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14467" *) _04629_;
  assign _07539_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14469" *) _04630_;
  assign _07540_ = nor_1672_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14471" *) _04631_;
  assign or_tmp_1375 = _07540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14471" *) cfg_mode_eql_1_sva_6;
  assign _07541_ = cfg_proc_precision_1_sva_st_102[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14485" *) nor_1672_cse;
  assign _07542_ = cfg_proc_precision_1_sva_st_90[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14488" *) nor_1672_cse;
  assign _07543_ = cfg_proc_precision_1_sva_st_102[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14490" *) _04632_;
  assign _07544_ = cfg_out_precision_1_sva_st_144[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14498" *) _04566_;
  assign _07545_ = cfg_out_precision_1_sva_st_156[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14500" *) _04634_;
  assign _07546_ = _04566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14501" *) cfg_mode_eql_1_sva_6;
  assign _07547_ = _07546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14502" *) _04150_;
  assign or_1644_nl = _07547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14502" *) cfg_out_precision_1_sva_st_156[0];
  assign or_5189_cse = _04635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14505" *) chn_out_rsci_bawt;
  assign _07548_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14505" *) _04631_;
  assign mux_tmp_1047 = _07548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14505" *) mux_tmp_1038;
  assign _07549_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14507" *) _01573_;
  assign _07550_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14509" *) _04582_;
  assign _07551_ = _07550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14509" *) cfg_mode_eql_1_sva_5;
  assign or_1643_nl = _07551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14509" *) or_1198_cse;
  assign or_tmp_1650 = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14513" *) _04637_;
  assign _07552_ = cfg_out_precision_1_sva_6[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14522" *) _04638_;
  assign or_1918_nl = _04566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14525" *) _04151_;
  assign _07553_ = cfg_out_precision_1_sva_st_156[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14527" *) _04639_;
  assign _07554_ = cfg_mode_eql_1_sva_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14528" *) _04150_;
  assign or_1745_nl = _07554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14529" *) cfg_out_precision_1_sva_st_156[0];
  assign _07555_ = nor_1589_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14534" *) _04566_;
  assign _07556_ = _07555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14535" *) cfg_mode_eql_1_sva_6;
  assign _07557_ = _07556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14535" *) _04150_;
  assign or_1774_nl = _07557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14535" *) cfg_out_precision_1_sva_st_156[0];
  assign mux_tmp_1109 = _07548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14538" *) mux_tmp_1100;
  assign _07558_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14540" *) _01574_;
  assign or_4667_nl = nor_151_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14541" *) or_578_cse;
  assign _07559_ = or_4667_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14542" *) _04582_;
  assign _07560_ = _07559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14542" *) cfg_mode_eql_1_sva_5;
  assign or_1773_nl = _07560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14542" *) or_1198_cse;
  assign or_tmp_1780 = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14546" *) _04641_;
  assign _07561_ = cfg_proc_precision_1_sva_st_102[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14557" *) nor_213_cse;
  assign _07562_ = cfg_proc_precision_1_sva_st_66[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14559" *) _04642_;
  assign or_tmp_1981 = or_1431_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14562" *) nand_202_cse;
  assign or_tmp_1992 = or_1157_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14563" *) nand_202_cse;
  assign _07563_ = cfg_proc_precision_1_sva_st_66[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14564" *) _04631_;
  assign _07564_ = cfg_proc_precision_1_sva_st_90[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14566" *) _04643_;
  assign _07565_ = cfg_proc_precision_1_sva_st_102[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14568" *) _04644_;
  assign or_513_cse = _04186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14571" *) cfg_mode_eql_1_sva_4;
  assign or_2289_cse = or_513_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14572" *) or_2251_nl;
  assign or_tmp_2136 = or_2289_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14572" *) _04185_;
  assign or_tmp_2139 = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14573" *) _00042_;
  assign or_2140_cse = nor_50_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14576" *) cfg_out_precision_1_sva_st_149[0];
  assign or_2232_nl = nor_151_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14601" *) cfg_out_precision_1_sva_st_149[0];
  assign _07566_ = _04645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14608" *) _04635_;
  assign or_2245_nl = _07566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14608" *) chn_out_rsci_bawt;
  assign _07567_ = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14612" *) _04635_;
  assign or_2246_nl = _07567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14612" *) chn_out_rsci_bawt;
  assign _07568_ = nor_8_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14614" *) nor_2150_cse;
  assign or_4569_nl = _07568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14615" *) or_2251_nl;
  assign _07569_ = or_4569_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14615" *) mux_tmp_1419;
  assign _07570_ = cvt_5_FpMantRNE_17U_11U_else_and_1_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14624" *) _00058_;
  assign or_2306_nl = _04647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14626" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign or_tmp_2432 = _00063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14628" *) cfg_mode_eql_rsci_d;
  assign or_tmp_2466 = IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14629" *) IsNaN_8U_23U_nor_4_tmp;
  assign or_tmp_2469 = IsNaN_8U_23U_nor_4_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14630" *) IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2;
  assign _07571_ = _04221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14633" *) _04635_;
  assign _07572_ = _07571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14633" *) chn_out_rsci_bawt;
  assign _07573_ = _07572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14633" *) _04185_;
  assign or_tmp_2569 = _07573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14633" *) or_4550_cse;
  assign _07574_ = _04220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14636" *) _04635_;
  assign _07575_ = _07574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14636" *) chn_out_rsci_bawt;
  assign _07576_ = _07575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14636" *) _04185_;
  assign or_tmp_2571 = _07576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14636" *) or_4550_cse;
  assign _07577_ = _04219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14639" *) _04635_;
  assign _07578_ = _07577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14639" *) chn_out_rsci_bawt;
  assign _07579_ = _07578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14639" *) _04185_;
  assign or_tmp_2573 = _07579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14639" *) or_4550_cse;
  assign _07580_ = _04218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14642" *) _04635_;
  assign _07581_ = _07580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14642" *) chn_out_rsci_bawt;
  assign _07582_ = _07581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14642" *) _04185_;
  assign or_tmp_2575 = _07582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14642" *) or_4550_cse;
  assign _07583_ = _04217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14645" *) _04635_;
  assign _07584_ = _07583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14645" *) chn_out_rsci_bawt;
  assign _07585_ = _07584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14645" *) _04185_;
  assign or_tmp_2577 = _07585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14645" *) or_4550_cse;
  assign _07586_ = _04216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14648" *) _04635_;
  assign _07587_ = _07586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14648" *) chn_out_rsci_bawt;
  assign _07588_ = _07587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14648" *) _04185_;
  assign or_tmp_2579 = _07588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14648" *) or_4550_cse;
  assign _07589_ = _04214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14651" *) _04635_;
  assign _07590_ = _07589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14651" *) chn_out_rsci_bawt;
  assign _07591_ = _07590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14651" *) _04185_;
  assign or_tmp_2588 = _07591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14651" *) or_4550_cse;
  assign _07592_ = _04213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14654" *) _04635_;
  assign _07593_ = _07592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14654" *) chn_out_rsci_bawt;
  assign _07594_ = _07593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14654" *) _04185_;
  assign or_tmp_2590 = _07594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14654" *) or_4550_cse;
  assign _07595_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14659" *) _04212_;
  assign _07596_ = _07595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14659" *) _04185_;
  assign or_tmp_2595 = _07596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14659" *) or_4550_cse;
  assign _07597_ = _04210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14662" *) _04635_;
  assign _07598_ = _07597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14662" *) chn_out_rsci_bawt;
  assign _07599_ = _07598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14662" *) _04185_;
  assign or_tmp_2604 = _07599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14662" *) or_4550_cse;
  assign _07600_ = _04209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14665" *) _04635_;
  assign _07601_ = _07600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14665" *) chn_out_rsci_bawt;
  assign _07602_ = _07601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14665" *) _04185_;
  assign or_tmp_2606 = _07602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14665" *) or_4550_cse;
  assign _07603_ = _04208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14668" *) _04635_;
  assign _07604_ = _07603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14668" *) chn_out_rsci_bawt;
  assign _07605_ = _07604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14668" *) _04185_;
  assign or_tmp_2608 = _07605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14668" *) or_4550_cse;
  assign _07606_ = _04207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14671" *) _04635_;
  assign _07607_ = _07606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14671" *) chn_out_rsci_bawt;
  assign _07608_ = _07607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14671" *) _04185_;
  assign or_tmp_2610 = _07608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14671" *) or_4550_cse;
  assign _07609_ = _04206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14674" *) _04635_;
  assign _07610_ = _07609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14674" *) chn_out_rsci_bawt;
  assign _07611_ = _07610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14674" *) _04185_;
  assign or_tmp_2612 = _07611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14674" *) or_4550_cse;
  assign or_dcpl_4 = and_dcpl_93 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14676" *) _04631_;
  assign or_dcpl_15 = and_dcpl_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14682" *) _03932_;
  assign _07612_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14698" *) _00058_;
  assign or_tmp_2960 = cfg_out_precision_1_sva_st_154[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14703" *) not_tmp_2254;
  assign _07613_ = nor_2219_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14724" *) nor_50_cse;
  assign or_tmp_3025 = _07613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14724" *) cfg_out_precision_1_sva_st_149[0];
  assign or_tmp_3032 = cfg_out_precision_1_sva_st_154[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14725" *) not_tmp_270;
  assign _07614_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14733" *) _00070_;
  assign or_dcpl_147 = or_4862_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14739" *) or_300_cse;
  assign _07615_ = nor_50_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14746" *) cfg_out_precision_1_sva_st_113[0];
  assign _07616_ = nor_1672_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14754" *) _04150_;
  assign or_dcpl_160 = and_1021_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14759" *) cfg_out_precision_1_sva_st_113[0];
  assign or_dcpl_163 = nor_50_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14762" *) and_dcpl_479;
  assign _07617_ = cfg_proc_precision_1_sva_st_102[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14764" *) _04653_;
  assign or_dcpl_181 = or_dcpl_178 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14769" *) and_dcpl_535;
  assign or_dcpl_184 = _04653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14770" *) and_dcpl_535;
  assign or_dcpl_188 = or_dcpl_184 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14772" *) and_1059_cse;
  assign or_dcpl_195 = _04632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14773" *) and_dcpl_535;
  assign or_dcpl_197 = or_dcpl_195 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14774" *) and_1059_cse;
  assign or_3817_cse = _00069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14777" *) and_1021_cse;
  assign _07618_ = or_3817_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14777" *) _00058_;
  assign or_dcpl_243 = and_1021_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14780" *) _00058_;
  assign _07619_ = _00069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14781" *) or_dcpl_243;
  assign _07620_ = _00070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14783" *) or_dcpl_243;
  assign _07621_ = _07450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14785" *) nor_50_cse;
  assign _07622_ = _07621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14786" *) _00058_;
  assign or_tmp_3379 = _07622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14786" *) or_578_cse;
  assign or_dcpl_277 = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14787" *) cfg_out_precision_1_sva_st_149[0];
  assign _07623_ = _04655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14789" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7];
  assign or_dcpl_320 = _07623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14789" *) _04656_;
  assign _07624_ = _04657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14791" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign or_dcpl_322 = _07624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14791" *) _04658_;
  assign _07625_ = _04659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14793" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign or_dcpl_324 = _07625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14793" *) _04660_;
  assign _07626_ = _04661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14795" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign or_dcpl_326 = _07626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14795" *) _04662_;
  assign _07627_ = _04663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14797" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign or_dcpl_328 = _07627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14797" *) _04664_;
  assign _07628_ = _04665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14799" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign or_dcpl_330 = _07628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14799" *) _04666_;
  assign _07629_ = _04667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14801" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign or_dcpl_332 = _07629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14801" *) _04668_;
  assign _07630_ = _04669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14803" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign or_dcpl_334 = _07630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14803" *) _04670_;
  assign _07631_ = _04671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14805" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign or_dcpl_336 = _07631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14805" *) _04672_;
  assign _07632_ = _04673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14807" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign or_dcpl_338 = _07632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14807" *) _04674_;
  assign _07633_ = _04675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14809" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign or_dcpl_340 = _07633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14809" *) _04676_;
  assign _07634_ = _04677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14811" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign or_dcpl_342 = _07634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14811" *) _04678_;
  assign _07635_ = _04679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14813" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign or_dcpl_344 = _07635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14813" *) _04680_;
  assign _07636_ = _04681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14815" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign or_dcpl_346 = _07636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14815" *) _04682_;
  assign _07637_ = _04683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14817" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign or_dcpl_348 = _07637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14817" *) _04684_;
  assign _07638_ = _04685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14819" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7];
  assign or_dcpl_350 = _07638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14819" *) _04686_;
  assign or_dcpl_353 = _04584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14820" *) and_1021_cse;
  assign or_dcpl_386 = and_dcpl_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14821" *) _04185_;
  assign or_dcpl_389 = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14822" *) or_1198_cse;
  assign or_dcpl_399 = and_dcpl_93 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14824" *) _00058_;
  assign _07639_ = nand_190_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14828" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign or_dcpl_420 = _07639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14828" *) cfg_out_precision_1_sva_st_149[0];
  assign _07640_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14832" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign or_dcpl_439 = _07640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14832" *) or_578_cse;
  assign _07641_ = nand_190_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14835" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign or_dcpl_448 = _07641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14835" *) cfg_out_precision_1_sva_st_149[0];
  assign or_dcpl_480 = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14839" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign _07642_ = nand_190_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14841" *) cfg_out_precision_1_sva_st_149[0];
  assign or_dcpl_490 = _07642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14841" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign or_dcpl_511 = and_dcpl_93 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14844" *) and_1021_cse;
  assign _07643_ = _00063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14850" *) _04687_;
  assign or_dcpl_612 = _07643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14850" *) and_dcpl_93;
  assign chn_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14852" *) fsm_output[0];
  assign _07644_ = _04689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14860" *) or_309_cse;
  assign _07645_ = _07644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14860" *) or_4862_cse;
  assign _07646_ = or_dcpl_353 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14879" *) cfg_out_precision_1_sva_st_113[0];
  assign _07647_ = _04692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14884" *) or_309_cse;
  assign _07648_ = _07647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14884" *) or_4862_cse;
  assign _07649_ = _07613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14969" *) nor_151_cse;
  assign _07650_ = _07649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14970" *) cfg_out_precision_1_sva_st_149[0];
  assign or_tmp_3763 = _07650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14970" *) nand_190_cse;
  assign or_tmp_3768 = _07613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14971" *) or_578_cse;
  assign or_tmp_3826 = cfg_proc_precision_1_sva_st_101[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14972" *) fsm_output[1];
  assign _07651_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *) cfg_proc_precision_1_sva_st_101[0];
  assign _07652_ = _07651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *) fsm_output[1];
  assign _07653_ = _04694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *) _04635_;
  assign or_tmp_3832 = _07653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14982" *) chn_out_rsci_bawt;
  assign _07654_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14983" *) cfg_proc_precision_1_sva_st_101[1];
  assign _07655_ = _04695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *) _00058_;
  assign _07656_ = _07655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *) cfg_proc_precision_1_sva_st_101[0];
  assign _07657_ = _07656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14984" *) fsm_output[1];
  assign _07658_ = _04696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14985" *) _04635_;
  assign or_4675_nl = _07658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14985" *) chn_out_rsci_bawt;
  assign _07659_ = _07613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14989" *) _00058_;
  assign _07660_ = _07659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14990" *) cfg_out_precision_1_sva_st_149[0];
  assign or_tmp_3840 = _07660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14990" *) _04697_;
  assign or_tmp_3849 = or_tmp_3768 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14992" *) _04698_;
  assign _07661_ = cvt_else_nor_dfs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14999" *) FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  assign or_tmp = _07661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:14999" *) cvt_else_equal_tmp_5;
  assign _07662_ = cvt_else_nor_dfs_10 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15003" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7;
  assign or_tmp_4080 = _07662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15003" *) cvt_else_equal_tmp_9;
  assign _07663_ = cvt_else_nor_dfs_10 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15009" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  assign or_tmp_4081 = _07663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15009" *) cvt_else_equal_tmp_16;
  assign _07664_ = cvt_else_nor_dfs_10 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15015" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  assign or_tmp_4082 = _07664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15015" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  assign _07665_ = cvt_else_nor_dfs_11 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15020" *) cvt_else_equal_tmp_33;
  assign or_tmp_4084 = _07665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15020" *) cvt_else_equal_tmp_34;
  assign _07666_ = reg_cvt_else_nor_dfs_9_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15027" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7;
  assign or_tmp_4086 = _07666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15027" *) cvt_else_equal_tmp_28;
  assign _07667_ = cvt_else_nor_dfs_10 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15032" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  assign or_tmp_4087 = _07667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15032" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  assign _07668_ = reg_cvt_else_nor_dfs_9_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15041" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7;
  assign or_tmp_4092 = _07668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15041" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  assign _07669_ = cvt_else_nor_dfs_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15045" *) cvt_else_equal_tmp_45;
  assign or_tmp_4095 = _07669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15045" *) cvt_else_equal_tmp_46;
  assign _07670_ = cvt_else_nor_dfs_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15051" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  assign or_tmp_4097 = _07670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15051" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  assign or_tmp_4102 = _01623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15057" *) cvt_asn_321;
  assign or_5174_tmp = _01625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15059" *) cvt_asn_321;
  assign or_5175_tmp = _01627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15061" *) cvt_asn_321;
  assign or_5176_tmp = _01629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15063" *) cvt_asn_321;
  assign or_5177_tmp = _01631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15065" *) cvt_asn_321;
  assign or_5178_tmp = _01633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15067" *) cvt_asn_321;
  assign or_5179_tmp = _01635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15069" *) cvt_asn_321;
  assign or_5180_tmp = _01637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15071" *) cvt_asn_321;
  assign or_5181_tmp = _01639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15073" *) cvt_asn_321;
  assign or_5182_tmp = _01641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15075" *) cvt_asn_321;
  assign or_5183_tmp = _01643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15077" *) cvt_asn_321;
  assign or_5184_tmp = _01645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15079" *) cvt_asn_321;
  assign or_5185_tmp = _01647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15081" *) cvt_asn_321;
  assign or_5186_tmp = _01649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15083" *) cvt_asn_321;
  assign or_5187_tmp = _01651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15085" *) cvt_asn_321;
  assign or_5188_tmp = _01653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15087" *) cvt_asn_321;
  assign _07671_ = _04733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15369" *) _04566_;
  assign _07672_ = _07671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15369" *) cfg_mode_eql_1_sva_6;
  assign _07673_ = _04734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15383" *) _04566_;
  assign _07674_ = _07673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15383" *) cfg_mode_eql_1_sva_6;
  assign _07675_ = _04735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15396" *) _04566_;
  assign _07676_ = _07675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15396" *) cfg_mode_eql_1_sva_6;
  assign _07677_ = _04736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15410" *) _04566_;
  assign _07678_ = _07677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15410" *) cfg_mode_eql_1_sva_6;
  assign _07679_ = _04737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15424" *) _04566_;
  assign _07680_ = _07679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15424" *) cfg_mode_eql_1_sva_6;
  assign _07681_ = _04738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15438" *) _04566_;
  assign _07682_ = _07681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15438" *) cfg_mode_eql_1_sva_6;
  assign _07683_ = _04739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15452" *) _04566_;
  assign _07684_ = _07683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15452" *) cfg_mode_eql_1_sva_6;
  assign _07685_ = _04740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15466" *) _04566_;
  assign _07686_ = _07685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15466" *) cfg_mode_eql_1_sva_6;
  assign _07687_ = _04741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15480" *) _04566_;
  assign _07688_ = _07687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15480" *) cfg_mode_eql_1_sva_6;
  assign _07689_ = mux_2362_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15514" *) _04566_;
  assign _07690_ = _07689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15514" *) cfg_mode_eql_1_sva_6;
  assign _07691_ = and_dcpl_103 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15621" *) and_dcpl_105;
  assign _07692_ = or_tmp_3487 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15629" *) main_stage_v_1_mx0c1;
  assign _07693_ = and_550_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16448" *) _01791_;
  assign _07694_ = _07693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16448" *) IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1;
  assign _07695_ = and_dcpl_114 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16522" *) main_stage_v_2_mx0c1;
  assign _07696_ = _04814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16668" *) _04815_;
  assign _07697_ = _04817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16670" *) _04818_;
  assign _07698_ = _04820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16672" *) _04821_;
  assign _07699_ = _04823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16674" *) _04824_;
  assign _07700_ = _04826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16676" *) _04827_;
  assign _07701_ = _04829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16678" *) _04830_;
  assign _07702_ = _04832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16680" *) _04833_;
  assign _07703_ = _04835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16682" *) _04836_;
  assign _07704_ = _04838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16684" *) _04839_;
  assign _07705_ = _04841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16686" *) _04842_;
  assign _07706_ = _04844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16688" *) _04845_;
  assign _07707_ = _04847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16690" *) _04848_;
  assign _07708_ = _04850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16692" *) _04851_;
  assign _07709_ = _01809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16717" *) and_637_rgt;
  assign _07710_ = _01813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16736" *) and_639_rgt;
  assign _07711_ = _01816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16759" *) and_641_rgt;
  assign _07712_ = _01819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16770" *) and_643_rgt;
  assign _07713_ = _01822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16781" *) and_646_rgt;
  assign _07714_ = _01826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16800" *) and_648_rgt;
  assign _07715_ = _01829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16831" *) and_650_rgt;
  assign _07716_ = _01832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16842" *) and_652_rgt;
  assign _07717_ = _01835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16853" *) and_654_rgt;
  assign _07718_ = _01838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16876" *) and_656_rgt;
  assign _07719_ = _01841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16887" *) and_658_rgt;
  assign _07720_ = _01844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16898" *) and_660_rgt;
  assign _07721_ = _01847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16909" *) and_662_rgt;
  assign _07722_ = _01850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16920" *) and_664_rgt;
  assign _07723_ = _01853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16931" *) and_666_rgt;
  assign _07724_ = _01857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16950" *) and_668_rgt;
  assign _07725_ = _01880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *) and_704_rgt;
  assign _07726_ = mux_2176_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17257" *) nor_2040_cse;
  assign _07727_ = _01889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *) and_719_rgt;
  assign _07728_ = _01898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *) and_734_rgt;
  assign _07729_ = _01906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *) and_749_rgt;
  assign _07730_ = mux_2186_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17443" *) nor_2040_cse;
  assign _07731_ = _01914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *) and_766_rgt;
  assign _07732_ = _01928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *) and_787_rgt;
  assign _07733_ = _01936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *) and_801_rgt;
  assign _07734_ = _01944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *) and_816_rgt;
  assign _07735_ = _01952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *) and_830_rgt;
  assign _07736_ = mux_2214_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17782" *) fsm_output[0];
  assign _07737_ = _01963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *) and_849_rgt;
  assign _07738_ = mux_2218_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17838" *) nor_2040_cse;
  assign _07739_ = _01972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *) and_866_rgt;
  assign _07740_ = mux_2223_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17894" *) nor_2040_cse;
  assign _07741_ = _01981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *) and_881_rgt;
  assign _07742_ = and_dcpl_401 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17954" *) main_stage_v_3_mx0c1;
  assign _07743_ = and_896_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18029" *) and_900_rgt;
  assign _07744_ = _07743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18029" *) and_dcpl_420;
  assign _07745_ = cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18136" *) cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  assign _07746_ = _07745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18136" *) and_dcpl_420;
  assign _07747_ = _01995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *) and_2360_cse;
  assign _07748_ = _07747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *) cvt_unequal_tmp_20;
  assign _07749_ = cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18186" *) cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  assign _07750_ = _07749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18186" *) and_dcpl_420;
  assign _07751_ = cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18283" *) cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _07752_ = _07751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18283" *) and_dcpl_420;
  assign _07753_ = and_dcpl_408 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18305" *) FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1;
  assign _07754_ = _07753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18305" *) FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2;
  assign _07755_ = and_954_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18349" *) and_956_rgt;
  assign _07756_ = _07755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18349" *) and_dcpl_420;
  assign _07757_ = and_dcpl_407 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18369" *) and_957_rgt;
  assign _07758_ = cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18381" *) cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1;
  assign _07759_ = _07758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18381" *) and_dcpl_420;
  assign _07760_ = cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18425" *) cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _07761_ = _07760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18425" *) and_dcpl_420;
  assign _07762_ = and_984_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18473" *) and_986_rgt;
  assign _07763_ = _07762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18473" *) and_dcpl_420;
  assign _07764_ = _02015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18486" *) cvt_unequal_tmp_20;
  assign _07765_ = _03933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18494" *) cvt_unequal_tmp_20;
  assign _07766_ = _07765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18494" *) and_2360_cse;
  assign _07767_ = and_987_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18512" *) and_989_rgt;
  assign _07768_ = _07767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18512" *) and_dcpl_420;
  assign _07769_ = cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18544" *) cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  assign _07770_ = _07769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18544" *) and_dcpl_420;
  assign _07771_ = mux_2239_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18575" *) and_2360_cse;
  assign _07772_ = and_1009_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18592" *) and_1011_rgt;
  assign _07773_ = _07772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18592" *) and_dcpl_420;
  assign _07774_ = cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18615" *) cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _07775_ = _07774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18615" *) and_dcpl_420;
  assign _07776_ = cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18639" *) cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  assign _07777_ = _07776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18639" *) and_dcpl_420;
  assign _07778_ = cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18663" *) cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  assign _07779_ = _07778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18663" *) and_dcpl_420;
  assign _07780_ = cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18687" *) cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _07781_ = _07780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18687" *) and_dcpl_420;
  assign _07782_ = cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18703" *) cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  assign _07783_ = _07782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18703" *) and_dcpl_420;
  assign _07784_ = _03964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18755" *) IntShiftRightSat_49U_6U_17U_oelse_mux_24_nl;
  assign _07785_ = _03965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18760" *) IntShiftRightSat_49U_6U_17U_oelse_mux_26_nl;
  assign _07786_ = _03966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18763" *) IntShiftRightSat_49U_6U_17U_oelse_mux_22_nl;
  assign _07787_ = _03967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18766" *) IntShiftRightSat_49U_6U_17U_oelse_mux_28_nl;
  assign _07788_ = _03968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18769" *) IntShiftRightSat_49U_6U_17U_oelse_mux_18_nl;
  assign _07789_ = _03969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18772" *) IntShiftRightSat_49U_6U_17U_oelse_mux_20_nl;
  assign _07790_ = _03970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18775" *) IntShiftRightSat_49U_6U_17U_oelse_mux_16_nl;
  assign _07791_ = _03971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18778" *) IntShiftRightSat_49U_6U_17U_oelse_mux_30_nl;
  assign _07792_ = _03972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18781" *) IntShiftRightSat_49U_6U_17U_oelse_mux_10_nl;
  assign _07793_ = _03973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18784" *) IntShiftRightSat_49U_6U_17U_oelse_mux_12_nl;
  assign _07794_ = _03974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18787" *) IntShiftRightSat_49U_6U_17U_oelse_mux_8_nl;
  assign _07795_ = _03975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18790" *) IntShiftRightSat_49U_6U_17U_oelse_mux_14_nl;
  assign _07796_ = _03976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18793" *) IntShiftRightSat_49U_6U_17U_oelse_mux_4_nl;
  assign _07797_ = _03977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18796" *) IntShiftRightSat_49U_6U_17U_oelse_mux_6_nl;
  assign _07798_ = _03978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18799" *) IntShiftRightSat_49U_6U_17U_oelse_mux_2_nl;
  assign _07799_ = _03979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18802" *) IntShiftRightSat_49U_6U_17U_oelse_mux_32_nl;
  assign _07800_ = or_dcpl_181 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18882" *) _04631_;
  assign _07801_ = or_dcpl_184 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18899" *) _04631_;
  assign _07802_ = or_dcpl_195 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18959" *) or_dcpl_4;
  assign _07803_ = _02056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18990" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  assign _07804_ = _02071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19027" *) and_1077_rgt;
  assign _07805_ = _02090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19062" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _07806_ = _02092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19065" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _07807_ = _02109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19103" *) and_1091_rgt;
  assign _07808_ = _02197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19261" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _07809_ = or_4862_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19576" *) cfg_out_precision_1_sva_st_113[0];
  assign _07810_ = _04952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19577" *) cfg_out_precision_1_sva_st_113[1];
  assign _07811_ = _04953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19577" *) cfg_mode_eql_1_sva_5;
  assign _07812_ = _04954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19586" *) cfg_mode_eql_1_sva_5;
  assign _07813_ = _02344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19609" *) and_1213_rgt;
  assign _07814_ = and_1249_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19663" *) and_1250_rgt;
  assign FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse = and_1249_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19700" *) and_1247_rgt;
  assign _07815_ = _02387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *) and_1321_rgt;
  assign _07816_ = _02393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20098" *) and_1325_rgt;
  assign _07817_ = _02399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20117" *) and_1329_rgt;
  assign _07818_ = _02405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20136" *) and_1333_rgt;
  assign _07819_ = _02411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20155" *) and_1337_rgt;
  assign _07820_ = _02417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20174" *) and_1341_rgt;
  assign _07821_ = _02423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20193" *) and_1345_rgt;
  assign _07822_ = _02429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20212" *) and_1349_rgt;
  assign _07823_ = _02435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20231" *) and_1353_rgt;
  assign _07824_ = _02441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20250" *) and_1357_rgt;
  assign _07825_ = _02447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20269" *) and_1361_rgt;
  assign _07826_ = _02453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20288" *) and_1365_rgt;
  assign _07827_ = _02459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20307" *) and_1369_rgt;
  assign _07828_ = _02465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20326" *) and_1373_rgt;
  assign _07829_ = _02471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20345" *) and_1377_rgt;
  assign _07830_ = _02477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20364" *) and_1381_rgt;
  assign _07831_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20374" *) IntSaturation_17U_16U_and_31_rgt;
  assign _07832_ = _07831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20374" *) IntSaturation_17U_16U_o_and_31_rgt;
  assign _07833_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20386" *) IntSaturation_17U_16U_and_29_rgt;
  assign _07834_ = _07833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20386" *) IntSaturation_17U_16U_o_and_29_rgt;
  assign _07835_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20398" *) IntSaturation_17U_16U_and_27_rgt;
  assign _07836_ = _07835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20398" *) IntSaturation_17U_16U_o_and_27_rgt;
  assign _07837_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20410" *) IntSaturation_17U_16U_and_25_rgt;
  assign _07838_ = _07837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20410" *) IntSaturation_17U_16U_o_and_25_rgt;
  assign _07839_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20422" *) IntSaturation_17U_16U_and_23_rgt;
  assign _07840_ = _07839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20422" *) IntSaturation_17U_16U_o_and_23_rgt;
  assign _07841_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20434" *) IntSaturation_17U_16U_and_21_rgt;
  assign _07842_ = _07841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20434" *) IntSaturation_17U_16U_o_and_21_rgt;
  assign _07843_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20446" *) IntSaturation_17U_16U_and_19_rgt;
  assign _07844_ = _07843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20446" *) IntSaturation_17U_16U_o_and_19_rgt;
  assign _07845_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20458" *) IntSaturation_17U_16U_and_17_rgt;
  assign _07846_ = _07845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20458" *) IntSaturation_17U_16U_o_and_17_rgt;
  assign _07847_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20470" *) IntSaturation_17U_16U_and_15_rgt;
  assign _07848_ = _07847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20470" *) IntSaturation_17U_16U_o_and_15_rgt;
  assign _07849_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20482" *) IntSaturation_17U_16U_and_13_rgt;
  assign _07850_ = _07849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20482" *) IntSaturation_17U_16U_o_and_13_rgt;
  assign _07851_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20494" *) IntSaturation_17U_16U_and_11_rgt;
  assign _07852_ = _07851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20494" *) IntSaturation_17U_16U_o_and_11_rgt;
  assign _07853_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20506" *) IntSaturation_17U_16U_and_9_rgt;
  assign _07854_ = _07853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20506" *) IntSaturation_17U_16U_o_and_9_rgt;
  assign _07855_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20518" *) IntSaturation_17U_16U_and_7_rgt;
  assign _07856_ = _07855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20518" *) IntSaturation_17U_16U_o_and_7_rgt;
  assign _07857_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20530" *) IntSaturation_17U_16U_and_5_rgt;
  assign _07858_ = _07857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20530" *) IntSaturation_17U_16U_o_and_5_rgt;
  assign _07859_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20542" *) IntSaturation_17U_16U_and_3_rgt;
  assign _07860_ = _07859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20542" *) IntSaturation_17U_16U_o_and_3_rgt;
  assign _07861_ = IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20554" *) IntSaturation_17U_16U_and_1_rgt;
  assign _07862_ = _07861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20554" *) IntSaturation_17U_16U_o_and_1_rgt;
  assign _07863_ = _02512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20581" *) cvt_9_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _07864_ = _02513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20583" *) cvt_5_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _07865_ = _02514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20585" *) cvt_3_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _07866_ = _02515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20587" *) cvt_1_IntSaturation_17U_16U_if_acc_nl[2];
  assign _07867_ = _02516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20589" *) cvt_16_IntSaturation_17U_16U_if_acc_4_nl[2];
  assign _07868_ = _02517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20591" *) cvt_15_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _07869_ = _02518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20593" *) cvt_13_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _07870_ = _02519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20595" *) cvt_12_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _07871_ = _02520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20597" *) cvt_11_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _07872_ = _02521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20599" *) cvt_10_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _07873_ = _02522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20601" *) cvt_8_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _07874_ = _02523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20603" *) cvt_7_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _07875_ = _02524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20605" *) cvt_6_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _07876_ = _02525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20607" *) cvt_4_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _07877_ = _02526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20609" *) cvt_2_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign _07878_ = _02544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20819" *) and_1467_rgt;
  assign _07879_ = and_dcpl_942 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20830" *) nor_50_cse;
  assign _07880_ = _07879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20830" *) and_dcpl_93;
  assign _07881_ = _07880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign _07882_ = _07881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *) or_dcpl_389;
  assign _07883_ = nor_50_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign _07884_ = _07883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *) or_dcpl_389;
  assign _07885_ = and_dcpl_946 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20848" *) or_dcpl_151;
  assign _07886_ = _07885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20848" *) or_dcpl_399;
  assign _07887_ = _07886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07888_ = _07887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *) or_578_cse;
  assign _07889_ = or_dcpl_151 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20857" *) _00058_;
  assign _07890_ = _07889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07891_ = _07890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *) or_578_cse;
  assign _07892_ = and_dcpl_950 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20866" *) _04584_;
  assign _07893_ = _07892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20866" *) or_dcpl_399;
  assign _07894_ = _07893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07895_ = _07894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *) or_578_cse;
  assign _07896_ = _04584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20875" *) _00058_;
  assign _07897_ = _07896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07898_ = _07897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *) or_578_cse;
  assign _07899_ = and_dcpl_954 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20884" *) _04584_;
  assign _07900_ = _07899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20884" *) and_1021_cse;
  assign _07901_ = _07900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *) and_dcpl_93;
  assign _07902_ = _07901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *) or_dcpl_420;
  assign _07903_ = or_dcpl_353 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *) or_dcpl_420;
  assign _07904_ = and_dcpl_958 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20902" *) or_dcpl_163;
  assign _07905_ = _07904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20902" *) or_dcpl_399;
  assign _07906_ = _07905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20903" *) or_578_cse;
  assign _07907_ = _07906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20903" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07908_ = or_dcpl_163 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20912" *) _00058_;
  assign _07909_ = _07908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20913" *) or_578_cse;
  assign _07910_ = _07909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20913" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07911_ = and_dcpl_962 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20922" *) or_dcpl_163;
  assign _07912_ = _07911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20922" *) and_1021_cse;
  assign _07913_ = _07912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *) and_dcpl_93;
  assign _07914_ = _07913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *) or_dcpl_439;
  assign _07915_ = or_3774_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *) or_dcpl_439;
  assign _07916_ = and_dcpl_966 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20940" *) or_dcpl_163;
  assign _07917_ = _07916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20940" *) and_1021_cse;
  assign _07918_ = _07917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *) and_dcpl_93;
  assign _07919_ = _07918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *) or_dcpl_448;
  assign _07920_ = or_3774_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *) or_dcpl_448;
  assign _07921_ = and_dcpl_970 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20958" *) nor_50_cse;
  assign _07922_ = _07921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20958" *) and_dcpl_479;
  assign _07923_ = _07922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20959" *) and_1021_cse;
  assign _07924_ = _07923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20959" *) and_dcpl_93;
  assign _07925_ = _07924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20959" *) _00058_;
  assign _07926_ = _07925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *) or_578_cse;
  assign _07927_ = _07926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign _07928_ = or_3774_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20968" *) _00058_;
  assign _07929_ = _07928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *) or_578_cse;
  assign _07930_ = _07929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign _07931_ = and_dcpl_974 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20977" *) _00069_;
  assign _07932_ = _07931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20977" *) or_dcpl_399;
  assign _07933_ = _07932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20978" *) or_578_cse;
  assign _07934_ = _07933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20978" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07935_ = _00069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20987" *) _00058_;
  assign _07936_ = _07935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20988" *) or_578_cse;
  assign _07937_ = _07936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20988" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _07938_ = and_dcpl_978 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20997" *) _00069_;
  assign _07939_ = _07938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20997" *) and_1021_cse;
  assign _07940_ = _07939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *) or_dcpl_480;
  assign _07941_ = _07940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *) and_dcpl_93;
  assign _07942_ = _07941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *) or_578_cse;
  assign _07943_ = or_3817_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *) or_dcpl_480;
  assign _07944_ = _07943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21006" *) or_578_cse;
  assign _07945_ = and_dcpl_982 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21015" *) _00069_;
  assign _07946_ = _07945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21015" *) and_1021_cse;
  assign _07947_ = _07946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *) and_dcpl_93;
  assign _07948_ = _07947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *) or_dcpl_490;
  assign _07949_ = or_3817_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *) or_dcpl_490;
  assign _07950_ = and_dcpl_987 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21033" *) nor_50_cse;
  assign _07951_ = _07950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21033" *) and_dcpl_479;
  assign _07952_ = _07951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21034" *) and_1021_cse;
  assign _07953_ = _07952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21034" *) or_578_cse;
  assign _07954_ = _07953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign _07955_ = _07954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *) _00058_;
  assign _07956_ = _07955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *) and_dcpl_93;
  assign _07957_ = or_3817_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *) or_578_cse;
  assign _07958_ = _07957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign _07959_ = _07958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21044" *) _00058_;
  assign _07960_ = and_dcpl_991 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21053" *) _00069_;
  assign _07961_ = _07960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *) or_578_cse;
  assign _07962_ = _07961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign _07963_ = _07962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *) _00058_;
  assign _07964_ = _07963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21054" *) or_dcpl_511;
  assign _07965_ = or_tmp_3025 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *) _04947_;
  assign _07966_ = _07965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign _07967_ = _07966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *) _00058_;
  assign _07968_ = _07967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21064" *) and_1021_cse;
  assign _07969_ = and_dcpl_995 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21073" *) nor_50_cse;
  assign _07970_ = _07969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21073" *) and_dcpl_479;
  assign _07971_ = _07970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *) or_578_cse;
  assign _07972_ = _07971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *) _00058_;
  assign _07973_ = _07972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign _07974_ = _07973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21074" *) or_dcpl_511;
  assign or_3151_cse = _00071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21083" *) or_578_cse;
  assign _07975_ = or_3151_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *) _00058_;
  assign _07976_ = _07975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign _07977_ = and_dcpl_999 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21092" *) nor_50_cse;
  assign _07978_ = _07977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21092" *) and_dcpl_479;
  assign _07979_ = _07978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *) or_578_cse;
  assign _07980_ = _07979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *) and_dcpl_93;
  assign _07981_ = _07980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *) and_1021_cse;
  assign _07982_ = _07981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *) _00058_;
  assign _07983_ = _07982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21093" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign _07984_ = _00070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21102" *) or_578_cse;
  assign _07985_ = _07984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *) _00058_;
  assign _07986_ = _07985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign _07987_ = and_dcpl_1003 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21111" *) _00069_;
  assign _07988_ = _07987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21111" *) or_dcpl_277;
  assign _07989_ = _07988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *) _04947_;
  assign _07990_ = _07989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign _07991_ = _07990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *) or_dcpl_511;
  assign _07992_ = _00069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21120" *) or_dcpl_277;
  assign _07993_ = _07992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *) _04947_;
  assign _07994_ = _07993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *) and_1021_cse;
  assign _07995_ = _07994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21121" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign _07996_ = or_dcpl_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21179" *) nand_171_cse;
  assign _07997_ = _07996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21179" *) cfg_out_precision_1_sva_st_154[0];
  assign _07998_ = or_dcpl_612 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21260" *) cfg_proc_precision_rsci_d[0];
  assign _07999_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21261" *) _04685_;
  assign _08000_ = _07999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21261" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7];
  assign _08001_ = _08000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *) _04686_;
  assign _08002_ = _08001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *) fsm_output[0];
  assign _08003_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21271" *) _04683_;
  assign _08004_ = _08003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21271" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08005_ = _08004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *) _04684_;
  assign _08006_ = _08005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *) fsm_output[0];
  assign _08007_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21281" *) _04681_;
  assign _08008_ = _08007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21281" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08009_ = _08008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *) _04682_;
  assign _08010_ = _08009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *) fsm_output[0];
  assign _08011_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21291" *) _04679_;
  assign _08012_ = _08011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21291" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08013_ = _08012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *) _04680_;
  assign _08014_ = _08013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *) fsm_output[0];
  assign _08015_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21301" *) _04677_;
  assign _08016_ = _08015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21301" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08017_ = _08016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *) _04678_;
  assign _08018_ = _08017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *) fsm_output[0];
  assign _08019_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21311" *) _04675_;
  assign _08020_ = _08019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21311" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08021_ = _08020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *) _04676_;
  assign _08022_ = _08021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *) fsm_output[0];
  assign _08023_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21321" *) _04673_;
  assign _08024_ = _08023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21321" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08025_ = _08024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *) _04674_;
  assign _08026_ = _08025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *) fsm_output[0];
  assign _08027_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21331" *) _04671_;
  assign _08028_ = _08027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21331" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08029_ = _08028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *) _04672_;
  assign _08030_ = _08029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *) fsm_output[0];
  assign _08031_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21341" *) _04669_;
  assign _08032_ = _08031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21341" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08033_ = _08032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *) _04670_;
  assign _08034_ = _08033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *) fsm_output[0];
  assign _08035_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21351" *) _04667_;
  assign _08036_ = _08035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21351" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08037_ = _08036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *) _04668_;
  assign _08038_ = _08037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *) fsm_output[0];
  assign _08039_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21361" *) _04665_;
  assign _08040_ = _08039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21361" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08041_ = _08040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *) _04666_;
  assign _08042_ = _08041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *) fsm_output[0];
  assign _08043_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21371" *) _04663_;
  assign _08044_ = _08043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21371" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08045_ = _08044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *) _04664_;
  assign _08046_ = _08045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *) fsm_output[0];
  assign _08047_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21381" *) _04661_;
  assign _08048_ = _08047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21381" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08049_ = _08048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *) _04662_;
  assign _08050_ = _08049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *) fsm_output[0];
  assign _08051_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21391" *) _04659_;
  assign _08052_ = _08051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21391" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08053_ = _08052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *) _04660_;
  assign _08054_ = _08053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *) fsm_output[0];
  assign _08055_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21401" *) _04657_;
  assign _08056_ = _08055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21401" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08057_ = _08056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *) _04658_;
  assign _08058_ = _08057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *) fsm_output[0];
  assign _08059_ = _07998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21411" *) _04655_;
  assign _08060_ = _08059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21411" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7];
  assign _08061_ = _08060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *) _04656_;
  assign _08062_ = _08061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *) fsm_output[0];
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_nl = _02625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21429" *) FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_1_nl = _02626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21431" *) FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_2_nl = _02627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21433" *) FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_3_nl = _02628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21435" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_4_nl = _02629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21437" *) FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_5_nl = _02630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21439" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_6_nl = _02631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21441" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_7_nl = _02632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21443" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_8_nl = _02633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21445" *) FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_9_nl = _02634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21447" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_10_nl = _02635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21449" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_11_nl = _02636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21451" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_12_nl = _02637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21453" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_13_nl = _02638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21455" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_14_nl = _02639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21457" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_15_nl = _02640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21459" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  assign cvt_or_48_nl = cvt_asn_321 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21460" *) cfg_mode_eql_1_sva_6;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_nl = _02641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21547" *) FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_1_nl = _02642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21574" *) FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_2_nl = _02643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21600" *) FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_3_nl = _02644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21627" *) FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_4_nl = _02645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21654" *) FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_5_nl = _02646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21681" *) FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_6_nl = _02647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21708" *) FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_7_nl = _02648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21735" *) FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_8_nl = _02649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21762" *) FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_9_nl = _02650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21789" *) FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_10_nl = _02651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21816" *) FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_11_nl = _02652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21843" *) FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_12_nl = _02653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21870" *) FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_14_nl = _02654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21920" *) FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_15_nl = _02655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21935" *) FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  assign _08063_ = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21960" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7];
  assign _08064_ = _08063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *) _04686_;
  assign _08065_ = _08064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *) or_4524_cse;
  assign _08066_ = _08065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21961" *) _00063_;
  assign _08067_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21964" *) _05071_;
  assign _08068_ = _08067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21965" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2;
  assign _08069_ = _08068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21965" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2;
  assign or_9_nl = _05072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21967" *) cfg_mode_eql_rsci_d;
  assign _08070_ = _02657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21970" *) or_4524_cse;
  assign or_11_nl = _05073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21970" *) cfg_mode_eql_rsci_d;
  assign _08071_ = cvt_1_FpMantRNE_24U_11U_else_and_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21971" *) or_4524_cse;
  assign or_13_nl = _05074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21972" *) cfg_mode_eql_rsci_d;
  assign or_17_nl = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21974" *) _04686_;
  assign _08072_ = _02660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21982" *) or_4550_cse;
  assign _08073_ = _05076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21982" *) cfg_mode_eql_1_sva_4;
  assign or_14_nl = _05071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21984" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2;
  assign _08074_ = nor_8_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21986" *) cfg_mode_eql_1_sva_4;
  assign _08075_ = IsNaN_8U_23U_land_1_lpi_1_dfm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21987" *) _04206_;
  assign _08076_ = or_14_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21992" *) _04635_;
  assign _08077_ = _08076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21992" *) chn_out_rsci_bawt;
  assign _08078_ = _08077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21993" *) _04185_;
  assign or_19_nl = _08078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21993" *) or_4550_cse;
  assign _08079_ = _05071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22001" *) _04635_;
  assign _08080_ = _08079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22001" *) chn_out_rsci_bawt;
  assign _08081_ = _08080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22002" *) _04185_;
  assign or_28_nl = _08081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22002" *) or_4550_cse;
  assign _08082_ = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22005" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08083_ = _08082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22006" *) _04683_;
  assign _08084_ = _08083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22006" *) or_4524_cse;
  assign _08085_ = _08084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22006" *) _00063_;
  assign _08086_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22009" *) _05077_;
  assign _08087_ = _08086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22010" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2;
  assign _08088_ = _08087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22010" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08089_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22013" *) _05077_;
  assign _08090_ = _08089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22017" *) _04635_;
  assign _08091_ = _08090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22017" *) chn_out_rsci_bawt;
  assign _08092_ = _08091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22018" *) _04185_;
  assign or_35_nl = _08092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22018" *) or_4550_cse;
  assign _08093_ = _05077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22024" *) _04635_;
  assign _08094_ = _08093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22024" *) chn_out_rsci_bawt;
  assign _08095_ = _08094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22025" *) _04185_;
  assign or_37_nl = _08095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22025" *) or_4550_cse;
  assign _08096_ = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22028" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08097_ = _08096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22029" *) _04681_;
  assign _08098_ = _08097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22029" *) or_4524_cse;
  assign _08099_ = _08098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22029" *) _00063_;
  assign _08100_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22032" *) _05078_;
  assign _08101_ = _08100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22033" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2;
  assign _08102_ = _08101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22033" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08103_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22036" *) _05078_;
  assign _08104_ = _08103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22040" *) _04635_;
  assign _08105_ = _08104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22040" *) chn_out_rsci_bawt;
  assign _08106_ = _08105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22041" *) _04185_;
  assign or_43_nl = _08106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22041" *) or_4550_cse;
  assign _08107_ = _05078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22047" *) _04635_;
  assign _08108_ = _08107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22047" *) chn_out_rsci_bawt;
  assign _08109_ = _08108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22048" *) _04185_;
  assign or_45_nl = _08109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22048" *) or_4550_cse;
  assign _08110_ = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22051" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08111_ = _08110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22052" *) _04679_;
  assign _08112_ = _08111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22052" *) or_4524_cse;
  assign _08113_ = _08112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22052" *) _00063_;
  assign _08114_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22055" *) _05079_;
  assign _08115_ = _08114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22056" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2;
  assign _08116_ = _08115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22056" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08117_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22059" *) _05079_;
  assign _08118_ = _08117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22063" *) _04635_;
  assign _08119_ = _08118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22063" *) chn_out_rsci_bawt;
  assign _08120_ = _08119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22064" *) _04185_;
  assign or_51_nl = _08120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22064" *) or_4550_cse;
  assign _08121_ = _05079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22070" *) _04635_;
  assign _08122_ = _08121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22070" *) chn_out_rsci_bawt;
  assign _08123_ = _08122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22071" *) _04185_;
  assign or_53_nl = _08123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22071" *) or_4550_cse;
  assign _08124_ = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22075" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2;
  assign _08125_ = _08124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22076" *) _05080_;
  assign _08126_ = _08125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22076" *) _04185_;
  assign or_56_nl = _08126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22076" *) or_4550_cse;
  assign _08127_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22079" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08128_ = _08127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22080" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2;
  assign _08129_ = _08128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22081" *) _05080_;
  assign _08130_ = _08129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22081" *) _04185_;
  assign or_58_nl = _08130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22081" *) or_4550_cse;
  assign _08131_ = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22083" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08132_ = _08131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22083" *) _04677_;
  assign _08133_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22087" *) _05080_;
  assign _08134_ = _08133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22087" *) _04185_;
  assign or_61_nl = _08134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22087" *) or_4550_cse;
  assign _08135_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22090" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2;
  assign _08136_ = _08135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22091" *) _05080_;
  assign _08137_ = _08136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22091" *) _04185_;
  assign or_63_nl = _08137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22091" *) or_4550_cse;
  assign _08138_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22100" *) _05080_;
  assign _08139_ = _08138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22100" *) _04185_;
  assign or_68_nl = _08139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22100" *) or_4550_cse;
  assign _08140_ = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22104" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2;
  assign _08141_ = _08140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22105" *) _05081_;
  assign _08142_ = _08141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22105" *) _04185_;
  assign or_71_nl = _08142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22105" *) or_4550_cse;
  assign _08143_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22108" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08144_ = _08143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22109" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2;
  assign _08145_ = _08144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22110" *) _05081_;
  assign _08146_ = _08145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22110" *) _04185_;
  assign or_73_nl = _08146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22110" *) or_4550_cse;
  assign _08147_ = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22112" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08148_ = _08147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22112" *) _04675_;
  assign _08149_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22116" *) _05081_;
  assign _08150_ = _08149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22116" *) _04185_;
  assign or_76_nl = _08150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22116" *) or_4550_cse;
  assign _08151_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22119" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2;
  assign _08152_ = _08151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22120" *) _05081_;
  assign _08153_ = _08152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22120" *) _04185_;
  assign or_78_nl = _08153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22120" *) or_4550_cse;
  assign _08154_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22129" *) _05081_;
  assign _08155_ = _08154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22129" *) _04185_;
  assign or_83_nl = _08155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22129" *) or_4550_cse;
  assign _08156_ = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22133" *) _04635_;
  assign _08157_ = _08156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22133" *) chn_out_rsci_bawt;
  assign _08158_ = _08157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22134" *) _04568_;
  assign _08159_ = _08158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22135" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2;
  assign _08160_ = _08159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22135" *) _04185_;
  assign or_88_nl = _08160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22135" *) or_4550_cse;
  assign _08161_ = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22137" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08162_ = _08161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22137" *) _04673_;
  assign _08163_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22141" *) _04568_;
  assign _08164_ = _08163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22142" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2;
  assign _08165_ = _08164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22142" *) _04185_;
  assign or_90_nl = _08165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22142" *) or_4550_cse;
  assign _08166_ = _08163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22151" *) _04185_;
  assign or_95_nl = _08166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22151" *) or_4550_cse;
  assign _08167_ = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22154" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08168_ = _08167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22155" *) _04671_;
  assign _08169_ = _08168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22155" *) or_4524_cse;
  assign _08170_ = _08169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22155" *) _00063_;
  assign _08171_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22158" *) _05082_;
  assign _08172_ = _08171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22159" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2;
  assign _08173_ = _08172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22159" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08174_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22162" *) _05082_;
  assign _08175_ = _08174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22166" *) _04635_;
  assign _08176_ = _08175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22166" *) chn_out_rsci_bawt;
  assign _08177_ = _08176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22167" *) _04185_;
  assign or_101_nl = _08177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22167" *) or_4550_cse;
  assign _08178_ = _05082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22173" *) _04635_;
  assign _08179_ = _08178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22173" *) chn_out_rsci_bawt;
  assign _08180_ = _08179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22174" *) _04185_;
  assign or_103_nl = _08180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22174" *) or_4550_cse;
  assign _08181_ = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22177" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08182_ = _08181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22178" *) _04669_;
  assign _08183_ = _08182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22178" *) or_4524_cse;
  assign _08184_ = _08183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22178" *) _00063_;
  assign _08185_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22181" *) _05083_;
  assign _08186_ = _08185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22182" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2;
  assign _08187_ = _08186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22182" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08188_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22185" *) _05083_;
  assign _08189_ = _08188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22189" *) _04635_;
  assign _08190_ = _08189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22189" *) chn_out_rsci_bawt;
  assign _08191_ = _08190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22190" *) _04185_;
  assign or_109_nl = _08191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22190" *) or_4550_cse;
  assign _08192_ = _05083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22196" *) _04635_;
  assign _08193_ = _08192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22196" *) chn_out_rsci_bawt;
  assign _08194_ = _08193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22197" *) _04185_;
  assign or_111_nl = _08194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22197" *) or_4550_cse;
  assign _08195_ = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22201" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2;
  assign _08196_ = _08195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22202" *) _05084_;
  assign _08197_ = _08196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22202" *) _04185_;
  assign or_114_nl = _08197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22202" *) or_4550_cse;
  assign _08198_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22206" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08199_ = _08198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22207" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2;
  assign _08200_ = _08199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22208" *) _05084_;
  assign _08201_ = _08200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22208" *) _04185_;
  assign or_116_nl = _08201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22208" *) or_4550_cse;
  assign _08202_ = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22210" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08203_ = _08202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22210" *) _04667_;
  assign _08204_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22214" *) _05084_;
  assign _08205_ = _08204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22214" *) _04185_;
  assign or_119_nl = _08205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22214" *) or_4550_cse;
  assign _08206_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22218" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2;
  assign _08207_ = _08206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22219" *) _05084_;
  assign _08208_ = _08207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22219" *) _04185_;
  assign or_121_nl = _08208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22219" *) or_4550_cse;
  assign _08209_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22228" *) _05084_;
  assign _08210_ = _08209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22228" *) _04185_;
  assign or_126_nl = _08210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22228" *) or_4550_cse;
  assign _08211_ = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22231" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08212_ = _08211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22232" *) _04665_;
  assign _08213_ = _08212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22232" *) or_4524_cse;
  assign _08214_ = _08213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22232" *) _00063_;
  assign _08215_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22235" *) _05085_;
  assign _08216_ = _08215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22236" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2;
  assign _08217_ = _08216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22236" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08218_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22239" *) _05085_;
  assign _08219_ = _08218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22243" *) _04635_;
  assign _08220_ = _08219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22243" *) chn_out_rsci_bawt;
  assign _08221_ = _08220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22244" *) _04185_;
  assign or_132_nl = _08221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22244" *) or_4550_cse;
  assign _08222_ = _05085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22250" *) _04635_;
  assign _08223_ = _08222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22250" *) chn_out_rsci_bawt;
  assign _08224_ = _08223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22251" *) _04185_;
  assign or_134_nl = _08224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22251" *) or_4550_cse;
  assign _08225_ = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22254" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08226_ = _08225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22255" *) _04663_;
  assign _08227_ = _08226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22255" *) or_4524_cse;
  assign _08228_ = _08227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22255" *) _00063_;
  assign _08229_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22258" *) _05086_;
  assign _08230_ = _08229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22259" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2;
  assign _08231_ = _08230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22259" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08232_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22262" *) _05086_;
  assign _08233_ = _08232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22266" *) _04635_;
  assign _08234_ = _08233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22266" *) chn_out_rsci_bawt;
  assign _08235_ = _08234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22267" *) _04185_;
  assign or_140_nl = _08235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22267" *) or_4550_cse;
  assign _08236_ = _05086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22273" *) _04635_;
  assign _08237_ = _08236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22273" *) chn_out_rsci_bawt;
  assign _08238_ = _08237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22274" *) _04185_;
  assign or_142_nl = _08238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22274" *) or_4550_cse;
  assign _08239_ = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22278" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2;
  assign _08240_ = _08239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22279" *) _05087_;
  assign _08241_ = _08240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22279" *) _04185_;
  assign or_145_nl = _08241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22279" *) or_4550_cse;
  assign _08242_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22283" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08243_ = _08242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22284" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2;
  assign _08244_ = _08243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22285" *) _05087_;
  assign _08245_ = _08244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22285" *) _04185_;
  assign or_147_nl = _08245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22285" *) or_4550_cse;
  assign _08246_ = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22287" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08247_ = _08246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22287" *) _04661_;
  assign _08248_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22291" *) _05087_;
  assign _08249_ = _08248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22291" *) _04185_;
  assign or_150_nl = _08249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22291" *) or_4550_cse;
  assign _08250_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22295" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2;
  assign _08251_ = _08250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22296" *) _05087_;
  assign _08252_ = _08251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22296" *) _04185_;
  assign or_152_nl = _08252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22296" *) or_4550_cse;
  assign _08253_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22305" *) _05087_;
  assign _08254_ = _08253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22305" *) _04185_;
  assign or_157_nl = _08254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22305" *) or_4550_cse;
  assign _08255_ = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22308" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08256_ = _08255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22309" *) _04659_;
  assign _08257_ = _08256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22309" *) or_4524_cse;
  assign _08258_ = _08257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22309" *) _00063_;
  assign _08259_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22312" *) _05088_;
  assign _08260_ = _08259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22313" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2;
  assign _08261_ = _08260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22313" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08262_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22316" *) _05088_;
  assign _08263_ = _08262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22320" *) _04635_;
  assign _08264_ = _08263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22320" *) chn_out_rsci_bawt;
  assign _08265_ = _08264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22321" *) _04185_;
  assign or_163_nl = _08265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22321" *) or_4550_cse;
  assign _08266_ = _05088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22327" *) _04635_;
  assign _08267_ = _08266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22327" *) chn_out_rsci_bawt;
  assign _08268_ = _08267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22328" *) _04185_;
  assign or_165_nl = _08268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22328" *) or_4550_cse;
  assign _08269_ = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22331" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08270_ = _08269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22332" *) _04657_;
  assign _08271_ = _08270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22332" *) or_4524_cse;
  assign _08272_ = _08271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22332" *) _00063_;
  assign _08273_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22335" *) _05089_;
  assign _08274_ = _08273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22336" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2;
  assign _08275_ = _08274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22336" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08276_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22339" *) _05089_;
  assign _08277_ = _08276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22343" *) _04635_;
  assign _08278_ = _08277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22343" *) chn_out_rsci_bawt;
  assign _08279_ = _08278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22344" *) _04185_;
  assign or_171_nl = _08279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22344" *) or_4550_cse;
  assign _08280_ = _05089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22350" *) _04635_;
  assign _08281_ = _08280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22350" *) chn_out_rsci_bawt;
  assign _08282_ = _08281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22351" *) _04185_;
  assign or_173_nl = _08282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22351" *) or_4550_cse;
  assign _08283_ = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22354" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7];
  assign _08284_ = _08283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22355" *) _04655_;
  assign _08285_ = _08284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22355" *) or_4524_cse;
  assign _08286_ = _08285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22355" *) _00063_;
  assign _08287_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22358" *) _05090_;
  assign _08288_ = _08287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22359" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2;
  assign _08289_ = _08288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22359" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2;
  assign _08290_ = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22362" *) _05090_;
  assign _08291_ = _08290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22366" *) _04635_;
  assign _08292_ = _08291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22366" *) chn_out_rsci_bawt;
  assign _08293_ = _08292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22367" *) _04185_;
  assign or_179_nl = _08293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22367" *) or_4550_cse;
  assign _08294_ = _05090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22373" *) _04635_;
  assign _08295_ = _08294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22373" *) chn_out_rsci_bawt;
  assign _08296_ = _08295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22374" *) _04185_;
  assign or_181_nl = _08296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22374" *) or_4550_cse;
  assign _08297_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22486" *) cfg_out_precision_1_sva_st_149[1];
  assign _08298_ = _08297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22486" *) cfg_proc_precision_1_sva_st_65[0];
  assign _08299_ = _08298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22486" *) nand_219_cse;
  assign _08300_ = or_961_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22543" *) _04578_;
  assign _08301_ = or_2251_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22550" *) _00066_;
  assign _08302_ = nor_2040_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22552" *) or_2251_nl;
  assign _08303_ = _08302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22553" *) _00066_;
  assign _08304_ = IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22579" *) cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  assign _08305_ = nor_2040_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22586" *) cfg_out_precision_1_sva_st_154[0];
  assign _08306_ = _08305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22586" *) not_tmp_270;
  assign _08307_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22590" *) _05091_;
  assign _08308_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22594" *) _05092_;
  assign _08309_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22597" *) _05093_;
  assign _08310_ = IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22615" *) cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  assign _08311_ = nor_2150_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22620" *) or_2251_nl;
  assign _08312_ = _08305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22625" *) not_tmp_119;
  assign _08313_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22634" *) _05094_;
  assign _08314_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22637" *) _05095_;
  assign _08315_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22650" *) _05096_;
  assign _08316_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22653" *) _05097_;
  assign _08317_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22666" *) _05098_;
  assign _08318_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22669" *) _05099_;
  assign _08319_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22702" *) _05100_;
  assign _08320_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22705" *) _05101_;
  assign _08321_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22720" *) _05102_;
  assign _08322_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22723" *) _05103_;
  assign _08323_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22738" *) _05104_;
  assign _08324_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22741" *) _05105_;
  assign _08325_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22747" *) _05106_;
  assign _08326_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22753" *) _05107_;
  assign _08327_ = _02690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22758" *) cfg_out_precision_1_sva_st_154[0];
  assign _08328_ = _08327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22758" *) _05108_;
  assign _08329_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22761" *) _05109_;
  assign _08330_ = or_961_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22765" *) _05108_;
  assign _08331_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22768" *) _05110_;
  assign _08332_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22781" *) _05111_;
  assign _08333_ = _02693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22798" *) cfg_out_precision_1_sva_st_154[0];
  assign _08334_ = _08333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22798" *) _05112_;
  assign _08335_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22801" *) _05113_;
  assign _08336_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22807" *) _05114_;
  assign _08337_ = cfg_out_precision_1_sva_st_154[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22811" *) _05115_;
  assign _08338_ = _02695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22823" *) cfg_out_precision_1_sva_st_154[0];
  assign _08339_ = _08338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22823" *) _05116_;
  assign _08340_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22826" *) _05117_;
  assign _08341_ = or_961_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22830" *) _05116_;
  assign _08342_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22833" *) _05118_;
  assign _08343_ = cfg_out_precision_1_sva_st_154[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22837" *) _05119_;
  assign _08344_ = nor_1056_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22879" *) chn_idata_data_sva_2_47_31_1[0];
  assign _08345_ = _05120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22880" *) or_300_cse;
  assign _08346_ = _08345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22880" *) _00058_;
  assign _08347_ = _08346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22880" *) cfg_mode_eql_1_sva_5;
  assign _08348_ = _05121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22883" *) _00058_;
  assign _08349_ = _08348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22883" *) cfg_mode_eql_1_sva_5;
  assign _08350_ = cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22887" *) chn_idata_data_sva_3_47_31_1[0];
  assign or_4532_nl = _05122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22890" *) or_1159_cse;
  assign or_1383_nl = _04631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22893" *) cfg_mode_eql_1_sva_6;
  assign _08351_ = or_1383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22893" *) mux_810_nl;
  assign _08352_ = _05123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22896" *) or_4862_cse;
  assign _08353_ = _08352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22896" *) or_300_cse;
  assign _08354_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22899" *) mux_812_nl;
  assign _08355_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22899" *) _05124_;
  assign _08356_ = _04689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22906" *) or_4862_cse;
  assign _08357_ = _08356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22906" *) or_300_cse;
  assign _08358_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22909" *) mux_819_nl;
  assign _08359_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22909" *) _05126_;
  assign _08360_ = cvt_1_FpMantRNE_17U_11U_else_and_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22916" *) or_1198_cse;
  assign or_1201_nl = _08360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22916" *) _05127_;
  assign _08361_ = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl[4] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *) _05128_;
  assign _08362_ = _05129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22918" *) or_1198_cse;
  assign _08363_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22923" *) cfg_mode_eql_1_sva_5;
  assign _08364_ = _08363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22923" *) mux_826_nl;
  assign _08365_ = _04165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22925" *) FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6;
  assign _08366_ = _08365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22925" *) cfg_out_precision_1_sva_6[0];
  assign or_1209_nl = _08366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22925" *) nand_207_cse;
  assign _08367_ = or_1383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22927" *) mux_828_nl;
  assign _08368_ = nor_2219_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22929" *) or_1198_cse;
  assign _08369_ = _05131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22932" *) or_4862_cse;
  assign _08370_ = _08369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22932" *) or_300_cse;
  assign _08371_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22935" *) mux_830_nl;
  assign _08372_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22935" *) _05132_;
  assign _08373_ = _05133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22948" *) or_4862_cse;
  assign _08374_ = _08373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22948" *) or_300_cse;
  assign _08375_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22951" *) mux_834_nl;
  assign _08376_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22951" *) _05134_;
  assign _08377_ = _05137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22966" *) or_4862_cse;
  assign _08378_ = _08377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22966" *) or_300_cse;
  assign _08379_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22969" *) mux_838_nl;
  assign _08380_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22969" *) _05138_;
  assign _08381_ = _05139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22976" *) or_300_cse;
  assign _08382_ = _08381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22976" *) _00058_;
  assign _08383_ = _08382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22976" *) cfg_mode_eql_1_sva_5;
  assign _08384_ = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22977" *) chn_idata_data_sva_2_175_159_1[0];
  assign _08385_ = _05140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22978" *) or_300_cse;
  assign _08386_ = _08385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22978" *) _00058_;
  assign _08387_ = _08386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22978" *) cfg_mode_eql_1_sva_5;
  assign _08388_ = _05139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22982" *) _00058_;
  assign _08389_ = _08388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22982" *) cfg_mode_eql_1_sva_5;
  assign _08390_ = cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22986" *) chn_idata_data_sva_3_175_159_1[0];
  assign or_4530_nl = _05141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22989" *) or_1159_cse;
  assign _08391_ = or_1383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22992" *) mux_848_nl;
  assign _08392_ = _05142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22995" *) or_4862_cse;
  assign _08393_ = _08392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22995" *) or_300_cse;
  assign _08394_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22998" *) mux_850_nl;
  assign _08395_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22998" *) _05143_;
  assign _08396_ = cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *) chn_idata_data_sva_2_511_1;
  assign _08397_ = _08396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *) _00058_;
  assign _08398_ = _08397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *) cvt_unequal_tmp_20;
  assign _08399_ = _08398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23005" *) cfg_mode_eql_1_sva_5;
  assign _08400_ = nor_1629_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23009" *) _04631_;
  assign _08401_ = _08400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23009" *) cvt_unequal_tmp_21;
  assign _08402_ = _08401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23010" *) cfg_mode_eql_1_sva_6;
  assign or_1280_nl = cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23013" *) IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3;
  assign _08403_ = _05144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23017" *) or_4862_cse;
  assign _08404_ = _08403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23017" *) or_300_cse;
  assign _08405_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23020" *) mux_860_nl;
  assign _08406_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23020" *) _05145_;
  assign _08407_ = _05146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23027" *) or_4862_cse;
  assign _08408_ = _08407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23027" *) or_300_cse;
  assign _08409_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23030" *) mux_864_nl;
  assign _08410_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23030" *) _05147_;
  assign _08411_ = _05148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23037" *) or_300_cse;
  assign _08412_ = _08411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23037" *) _00058_;
  assign _08413_ = _08412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23037" *) cfg_mode_eql_1_sva_5;
  assign _08414_ = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23038" *) chn_idata_data_sva_2_495_479_1[0];
  assign _08415_ = _05149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23039" *) or_300_cse;
  assign _08416_ = _08415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23039" *) _00058_;
  assign _08417_ = _08416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23039" *) cfg_mode_eql_1_sva_5;
  assign _08418_ = _05148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23043" *) _00058_;
  assign _08419_ = _08418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23043" *) cfg_mode_eql_1_sva_5;
  assign _08420_ = cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23047" *) chn_idata_data_sva_3_495_479_1[0];
  assign or_4528_nl = _05150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23050" *) or_1159_cse;
  assign _08421_ = or_1383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23053" *) mux_874_nl;
  assign _08422_ = _05151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23056" *) or_4862_cse;
  assign _08423_ = _08422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23056" *) or_300_cse;
  assign _08424_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23059" *) mux_876_nl;
  assign _08425_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23059" *) _05152_;
  assign _08426_ = _05153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23066" *) or_300_cse;
  assign _08427_ = _08426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23066" *) _00058_;
  assign _08428_ = _08427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23066" *) cfg_mode_eql_1_sva_5;
  assign _08429_ = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23067" *) chn_idata_data_sva_2_239_223_1[0];
  assign _08430_ = _05154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23068" *) or_300_cse;
  assign _08431_ = _08430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23068" *) _00058_;
  assign _08432_ = _08431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23068" *) cfg_mode_eql_1_sva_5;
  assign _08433_ = _05153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23072" *) _00058_;
  assign _08434_ = _08433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23072" *) cfg_mode_eql_1_sva_5;
  assign _08435_ = cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23076" *) chn_idata_data_sva_3_239_223_1[0];
  assign or_4526_nl = _05155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23079" *) or_1159_cse;
  assign _08436_ = or_1383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23082" *) mux_886_nl;
  assign _08437_ = _05156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23085" *) or_4862_cse;
  assign _08438_ = _08437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23085" *) or_300_cse;
  assign _08439_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23088" *) mux_888_nl;
  assign _08440_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23088" *) _05157_;
  assign _08441_ = cvt_6_FpMantRNE_17U_11U_else_and_2_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *) _05158_;
  assign _08442_ = _08441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23096" *) or_578_cse;
  assign _08443_ = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23098" *) _05160_;
  assign _08444_ = _05162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *) or_578_cse;
  assign or_1374_nl = _05161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23099" *) _05164_;
  assign or_1375_nl = _08363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23105" *) mux_895_nl;
  assign _08445_ = _04151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  assign _08446_ = _08445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *) nor_183_cse;
  assign _08447_ = _08446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *) nor_213_cse;
  assign _08448_ = _08447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *) _04150_;
  assign or_1379_nl = _08448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23107" *) or_tmp_1375;
  assign or_1196_cse = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23112" *) or_300_cse;
  assign _08449_ = _05165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23113" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _08450_ = _05166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23114" *) or_1198_cse;
  assign or_1393_nl = _08450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23114" *) _05167_;
  assign _08451_ = or_5069_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23117" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _08452_ = _05168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23118" *) or_1198_cse;
  assign or_1399_nl = _08452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23118" *) _05167_;
  assign or_1396_nl = _05169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23119" *) cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign _08453_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23122" *) mux_904_nl;
  assign or_1402_nl = cvt_unequal_tmp_21 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23125" *) or_1157_cse;
  assign _08454_ = _04151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  assign _08455_ = _08454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *) nor_183_cse;
  assign _08456_ = _08455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *) nor_213_cse;
  assign _08457_ = _08456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *) nor_1589_cse;
  assign or_1409_nl = _08457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23127" *) _04150_;
  assign _08458_ = or_1383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23129" *) mux_908_nl;
  assign or_4793_nl = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23132" *) _05170_;
  assign _08459_ = _05171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23135" *) or_4862_cse;
  assign _08460_ = _08459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23135" *) or_300_cse;
  assign _08461_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23138" *) mux_910_nl;
  assign _08462_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23138" *) _05172_;
  assign _08463_ = _05173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23145" *) or_300_cse;
  assign _08464_ = _08463_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23145" *) _00058_;
  assign _08465_ = _08464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23145" *) cfg_mode_eql_1_sva_5;
  assign _08466_ = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23146" *) chn_idata_data_sva_2_271_255_1[0];
  assign _08467_ = _05174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23147" *) or_300_cse;
  assign _08468_ = _08467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23147" *) _00058_;
  assign _08469_ = _08468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23147" *) cfg_mode_eql_1_sva_5;
  assign _08470_ = or_425_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23151" *) _00058_;
  assign _08471_ = _08470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23151" *) cfg_mode_eql_1_sva_5;
  assign _08472_ = _05173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23153" *) _00058_;
  assign _08473_ = _08472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23153" *) cfg_mode_eql_1_sva_5;
  assign _08474_ = cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23160" *) chn_idata_data_sva_3_271_255_1[0];
  assign _08475_ = or_1383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23162" *) mux_920_nl;
  assign _08476_ = _05175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23165" *) or_4862_cse;
  assign _08477_ = _08476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23165" *) or_300_cse;
  assign _08478_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23168" *) mux_922_nl;
  assign _08479_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23168" *) _05176_;
  assign _08480_ = _05177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23175" *) or_4862_cse;
  assign _08481_ = _08480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23175" *) or_300_cse;
  assign _08482_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23178" *) mux_926_nl;
  assign _08483_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23178" *) _05178_;
  assign _08484_ = _05179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23185" *) or_4862_cse;
  assign _08485_ = _08484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23185" *) or_300_cse;
  assign _08486_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23188" *) mux_930_nl;
  assign _08487_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23188" *) _05180_;
  assign _08488_ = _05181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23195" *) or_4862_cse;
  assign _08489_ = _08488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23195" *) or_300_cse;
  assign _08490_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23198" *) mux_934_nl;
  assign _08491_ = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23198" *) _05182_;
  assign _08492_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23300" *) _04582_;
  assign or_1483_nl = _08492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23300" *) cfg_mode_eql_1_sva_5;
  assign _08493_ = cvt_1_IntSaturation_17U_8U_if_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23302" *) _00058_;
  assign _08494_ = _08493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23302" *) _04582_;
  assign or_1484_nl = _08494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23302" *) cfg_mode_eql_1_sva_5;
  assign _08495_ = cfg_out_precision_1_sva_st_113[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23304" *) mux_939_nl;
  assign _08496_ = _04631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23306" *) _04566_;
  assign _08497_ = _08496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23307" *) cfg_mode_eql_1_sva_6;
  assign _08498_ = _08497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23307" *) cfg_out_precision_1_sva_6[0];
  assign _08499_ = _04166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23308" *) cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2;
  assign _08500_ = _05183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23309" *) cfg_out_precision_1_sva_6[1];
  assign _08501_ = _08498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23309" *) _05184_;
  assign _08502_ = cfg_proc_precision_1_sva_st_90[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23316" *) _05185_;
  assign _08503_ = or_1483_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23322" *) cfg_out_precision_1_sva_st_113[0];
  assign _08504_ = or_461_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *) cvt_3_IntSaturation_17U_8U_if_acc_1_nl[10];
  assign _08505_ = _08504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *) nor_2219_cse;
  assign _08506_ = cfg_out_precision_1_sva_st_113[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *) _05186_;
  assign _08507_ = _08503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23324" *) _05187_;
  assign _08508_ = _04167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *) cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  assign _08509_ = _08508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *) nor_213_cse;
  assign _08510_ = cfg_out_precision_1_sva_6[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *) _05188_;
  assign _08511_ = _08498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23328" *) _05189_;
  assign _08512_ = or_461_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *) cvt_5_IntSaturation_17U_8U_if_acc_1_nl[10];
  assign _08513_ = _08512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *) nor_2219_cse;
  assign _08514_ = cfg_out_precision_1_sva_st_113[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *) _05190_;
  assign _08515_ = _08503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23334" *) _05191_;
  assign _08516_ = _04167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *) cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  assign _08517_ = _08516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *) nor_213_cse;
  assign _08518_ = cfg_out_precision_1_sva_6[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *) _05192_;
  assign _08519_ = _08498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23338" *) _05193_;
  assign _08520_ = or_461_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *) cvt_9_IntSaturation_17U_8U_if_acc_1_nl[10];
  assign _08521_ = _08520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *) nor_2219_cse;
  assign _08522_ = cfg_out_precision_1_sva_st_113[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *) _05194_;
  assign _08523_ = _08503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23344" *) _05195_;
  assign _08524_ = _04167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *) cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  assign _08525_ = _08524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *) nor_213_cse;
  assign _08526_ = cfg_out_precision_1_sva_6[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *) _05196_;
  assign _08527_ = _08498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23348" *) _05197_;
  assign or_3841_nl = and_dcpl_942 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23350" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign _08528_ = or_dcpl_389 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23356" *) _04582_;
  assign _08529_ = _08528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23356" *) cfg_mode_eql_1_sva_5;
  assign _08530_ = _08529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23356" *) nor_50_cse;
  assign _08531_ = _07540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *) _04566_;
  assign _08532_ = _08531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *) cfg_mode_eql_1_sva_6;
  assign _08533_ = _08532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *) _04150_;
  assign _08534_ = _08533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23358" *) _04165_;
  assign _08535_ = _02723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23365" *) or_1198_cse;
  assign _08536_ = _08535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign _08537_ = _08536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  assign _08538_ = _08537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23366" *) _05199_;
  assign _08539_ = _07548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23369" *) _04166_;
  assign _08540_ = _08539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23369" *) nor_1672_cse;
  assign _08541_ = _04631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23371" *) _04166_;
  assign _08542_ = _08541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23371" *) nor_1672_cse;
  assign or_3850_nl = and_dcpl_946 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23374" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _08543_ = _02725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23381" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _08544_ = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23382" *) _05202_;
  assign _08545_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23391" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _08546_ = _08545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23391" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _08547_ = _08546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23392" *) nor_2219_cse;
  assign _08548_ = _02726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *) or_1198_cse;
  assign _08549_ = _08547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23394" *) _05205_;
  assign or_3860_nl = and_dcpl_950 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23396" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign or_3879_nl = and_dcpl_958 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23401" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _08550_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23410" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _08551_ = _08550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23410" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _08552_ = _08551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23411" *) nor_2219_cse;
  assign _08553_ = _02728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *) or_1198_cse;
  assign _08554_ = _08552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23413" *) _05208_;
  assign _08555_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23424" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign _08556_ = _08555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23424" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _08557_ = _08556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23425" *) nor_2219_cse;
  assign _08558_ = _08557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23425" *) nor_151_cse;
  assign _08559_ = _02730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *) or_1198_cse;
  assign _08560_ = _08558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23427" *) _05211_;
  assign _08561_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23433" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _08562_ = _08561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23433" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _08563_ = _08562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23434" *) nor_2219_cse;
  assign _08564_ = _02732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *) or_1198_cse;
  assign _08565_ = _08563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23436" *) _05214_;
  assign _08566_ = _07548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23439" *) _04167_;
  assign _08567_ = _08566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23439" *) _04653_;
  assign _08568_ = _04631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23441" *) _04167_;
  assign _08569_ = _08568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23441" *) _04653_;
  assign _08570_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23451" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign _08571_ = _08570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23451" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _08572_ = _08571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23452" *) nor_2219_cse;
  assign _08573_ = _08572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23452" *) nor_151_cse;
  assign _08574_ = _02734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *) or_1198_cse;
  assign _08575_ = _08573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23454" *) _05217_;
  assign _08576_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23463" *) FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign _08577_ = _08576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23463" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _08578_ = _08577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23464" *) nor_2219_cse;
  assign _08579_ = _08578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23464" *) nor_151_cse;
  assign _08580_ = _02736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *) or_1198_cse;
  assign _08581_ = _08579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23466" *) _05220_;
  assign _08582_ = or_578_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23479" *) FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign _08583_ = _08582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23479" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _08584_ = _08583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23480" *) nor_2219_cse;
  assign _08585_ = _08584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23480" *) nor_151_cse;
  assign _08586_ = _02738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *) or_1198_cse;
  assign _08587_ = _08585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23482" *) _05223_;
  assign or_3920_nl = and_dcpl_974 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23484" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _08588_ = _07478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23490" *) _04582_;
  assign _08589_ = _08588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23490" *) cfg_mode_eql_1_sva_5;
  assign _08590_ = _08589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23491" *) or_1198_cse;
  assign _08591_ = _08590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23491" *) _04591_;
  assign _08592_ = nor_2219_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23496" *) or_578_cse;
  assign _08593_ = _08592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23497" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _08594_ = _08593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23498" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _08595_ = _02740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *) or_1198_cse;
  assign _08596_ = _08594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23500" *) _05226_;
  assign _08597_ = _08592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23508" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign _08598_ = _08597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23509" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _08599_ = _02743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *) or_1198_cse;
  assign _08600_ = _08598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23511" *) _05229_;
  assign _08601_ = _08592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23520" *) FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign _08602_ = _08601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23521" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _08603_ = _02745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *) or_1198_cse;
  assign _08604_ = _08602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23523" *) _05232_;
  assign _08605_ = cfg_proc_precision_1_sva_st_108[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23530" *) _05234_;
  assign _08606_ = _08592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23541" *) FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign _08607_ = _08606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23542" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _08608_ = _02748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *) or_1198_cse;
  assign _08609_ = _08607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23544" *) _05237_;
  assign _08610_ = _08592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23552" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign _08611_ = _08610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _08612_ = _08611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *) or_1198_cse;
  assign _08613_ = _02750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23553" *) _05241_;
  assign _08614_ = _07649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23556" *) or_425_cse;
  assign _08615_ = _07649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23562" *) or_300_cse;
  assign _08616_ = _08592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23573" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign _08617_ = _08616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _08618_ = _08617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *) or_1198_cse;
  assign _08619_ = _02759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23574" *) _05246_;
  assign _08620_ = _08592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23582" *) FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign _08621_ = _08620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _08622_ = _08621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *) or_1198_cse;
  assign _08623_ = _02762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23583" *) _05249_;
  assign _08624_ = _07450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23591" *) or_578_cse;
  assign _08625_ = _08624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23591" *) FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign _08626_ = _08625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2;
  assign _08627_ = _08626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *) or_1198_cse;
  assign _08628_ = _02765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23592" *) _05252_;
  assign _08629_ = cfg_proc_precision_1_sva_st_108[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23595" *) _05253_;
  assign _08630_ = or_5189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23599" *) _05254_;
  assign _08631_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23602" *) _04650_;
  assign or_4857_nl = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23603" *) cfg_proc_precision_1_sva_st_65[0];
  assign _08632_ = _04582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23606" *) or_4862_cse;
  assign or_3623_cse = nor_8_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23619" *) cfg_out_precision_1_sva_st_154[0];
  assign _08633_ = or_3623_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23620" *) _05255_;
  assign _08634_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23622" *) _05256_;
  assign _08635_ = or_2140_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23625" *) _05257_;
  assign or_2433_nl = _04168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23629" *) cfg_proc_precision_rsci_d[0];
  assign _08636_ = _08066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23636" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp;
  assign _08637_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23639" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2;
  assign _08638_ = _08637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23640" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2;
  assign _08639_ = _08638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23640" *) IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  assign _08640_ = _08639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23641" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2;
  assign _08641_ = _08640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23642" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2;
  assign _08642_ = _08641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23642" *) nand_164_cse;
  assign _08643_ = _02769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23645" *) _04685_;
  assign _08644_ = _08643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23646" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7];
  assign _08645_ = _08644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23646" *) _04686_;
  assign _08646_ = _08645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23647" *) or_4524_cse;
  assign _08647_ = _08646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23647" *) _00063_;
  assign _08648_ = _08647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23647" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp;
  assign _08649_ = _08637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23651" *) _05258_;
  assign _08650_ = _08649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23651" *) IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  assign _08651_ = _08650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23652" *) _05259_;
  assign _08652_ = _08651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23653" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2;
  assign _08653_ = _08652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23653" *) nand_164_cse;
  assign _08654_ = _08085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23659" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp;
  assign _08655_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23662" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2;
  assign _08656_ = _08655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23663" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08657_ = _08656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23663" *) IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  assign _08658_ = _08657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23664" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _08659_ = _08658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23665" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2;
  assign _08660_ = _08659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23665" *) nand_162_cse;
  assign _08661_ = _02770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23668" *) _04684_;
  assign _08662_ = _08661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23669" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08663_ = _08662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23669" *) _04683_;
  assign _08664_ = _08663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23670" *) or_4524_cse;
  assign _08665_ = _08664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23670" *) _00063_;
  assign _08666_ = _08665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23670" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp;
  assign _08667_ = _08655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23674" *) _05260_;
  assign _08668_ = _08667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23674" *) IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  assign _08669_ = _08668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23675" *) _05261_;
  assign _08670_ = _08669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23676" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2;
  assign _08671_ = _08670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23676" *) nand_162_cse;
  assign _08672_ = _08099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23682" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp;
  assign _08673_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23685" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2;
  assign _08674_ = _08673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23686" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08675_ = _08674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23686" *) IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  assign _08676_ = _08675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23687" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _08677_ = _08676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23688" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2;
  assign _08678_ = _08677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23688" *) nand_160_cse;
  assign _08679_ = _02771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23691" *) _04682_;
  assign _08680_ = _08679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23692" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08681_ = _08680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23692" *) _04681_;
  assign _08682_ = _08681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23693" *) or_4524_cse;
  assign _08683_ = _08682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23693" *) _00063_;
  assign _08684_ = _08683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23693" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp;
  assign _08685_ = _08673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23697" *) _05262_;
  assign _08686_ = _08685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23697" *) IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  assign _08687_ = _08686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23698" *) _05263_;
  assign _08688_ = _08687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23699" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2;
  assign _08689_ = _08688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23699" *) nand_160_cse;
  assign _08690_ = _08113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23705" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp;
  assign _08691_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23708" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2;
  assign _08692_ = _08691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23709" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08693_ = _08692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23709" *) IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  assign _08694_ = _08693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23710" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _08695_ = _08694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23711" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2;
  assign _08696_ = _08695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23711" *) nand_158_cse;
  assign _08697_ = _02772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23714" *) _04680_;
  assign _08698_ = _08697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23715" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08699_ = _08698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23715" *) _04679_;
  assign _08700_ = _08699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23716" *) or_4524_cse;
  assign _08701_ = _08700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23716" *) _00063_;
  assign _08702_ = _08701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23716" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp;
  assign _08703_ = _08691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23720" *) _05264_;
  assign _08704_ = _08703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23720" *) IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  assign _08705_ = _08704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23721" *) _05265_;
  assign _08706_ = _08705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23722" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2;
  assign _08707_ = _08706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23722" *) nand_158_cse;
  assign _08708_ = _05266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23727" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign _08709_ = _08708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23727" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08710_ = _08709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23728" *) _04677_;
  assign _08711_ = _08710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23728" *) or_4524_cse;
  assign _08712_ = _08711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23728" *) _00063_;
  assign _08713_ = nor_1099_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23729" *) _04185_;
  assign _08714_ = _08713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23730" *) or_4550_cse;
  assign _08715_ = _08714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23731" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2;
  assign _08716_ = _08715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23732" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08717_ = _08716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23733" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _08718_ = _08717_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23734" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2;
  assign _08719_ = _08718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23734" *) nand_156_cse;
  assign _08720_ = _02773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23739" *) _05267_;
  assign _08721_ = _08715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23743" *) _05268_;
  assign _08722_ = _08721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23744" *) _05269_;
  assign _08723_ = _08722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23745" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2;
  assign _08724_ = _08723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23745" *) nand_156_cse;
  assign _08725_ = _08148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23751" *) or_4524_cse;
  assign _08726_ = _08725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23751" *) _00063_;
  assign _08727_ = _08726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23751" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp;
  assign _08728_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23754" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2;
  assign _08729_ = _08728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23755" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08730_ = _08729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23755" *) IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  assign _08731_ = _08730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23756" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _08732_ = _08731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23757" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2;
  assign _08733_ = _08732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23757" *) nand_153_cse;
  assign _08734_ = _02779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23760" *) _04676_;
  assign _08735_ = _08734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23761" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08736_ = _08735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23761" *) _04675_;
  assign _08737_ = _08736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23762" *) or_4524_cse;
  assign _08738_ = _08737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23762" *) _00063_;
  assign _08739_ = _08738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23762" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp;
  assign _08740_ = _08728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23766" *) _05270_;
  assign _08741_ = _08740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23766" *) IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  assign _08742_ = _08741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23767" *) _05271_;
  assign _08743_ = _08742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23768" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2;
  assign _08744_ = _08743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23768" *) nand_153_cse;
  assign _08745_ = _08162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23774" *) or_4524_cse;
  assign _08746_ = _08745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23774" *) _00063_;
  assign _08747_ = _08746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23774" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp;
  assign _08748_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23777" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2;
  assign _08749_ = _08748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23778" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08750_ = _08749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23778" *) IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  assign _08751_ = _08750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23779" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _08752_ = _08751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23780" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2;
  assign _08753_ = _08752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23780" *) nand_151_cse;
  assign _08754_ = _02780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23783" *) _04674_;
  assign _08755_ = _08754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23784" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08756_ = _08755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23784" *) _04673_;
  assign _08757_ = _08756_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23785" *) or_4524_cse;
  assign _08758_ = _08757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23785" *) _00063_;
  assign _08759_ = _08758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23785" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp;
  assign _08760_ = _08748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23789" *) _05272_;
  assign _08761_ = _08760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23789" *) IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  assign _08762_ = _08761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23790" *) _05273_;
  assign _08763_ = _08762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23791" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2;
  assign _08764_ = _08763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23791" *) nand_151_cse;
  assign _08765_ = _08170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23797" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp;
  assign _08766_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23800" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2;
  assign _08767_ = _08766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23801" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08768_ = _08767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23801" *) IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  assign _08769_ = _08768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23802" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _08770_ = _08769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23803" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2;
  assign _08771_ = _08770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23803" *) nand_149_cse;
  assign _08772_ = _02781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23806" *) _04672_;
  assign _08773_ = _08772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23807" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08774_ = _08773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23807" *) _04671_;
  assign _08775_ = _08774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23808" *) or_4524_cse;
  assign _08776_ = _08775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23808" *) _00063_;
  assign _08777_ = _08776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23808" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp;
  assign _08778_ = _08766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23812" *) _05274_;
  assign _08779_ = _08778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23812" *) IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  assign _08780_ = _08779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23813" *) _05275_;
  assign _08781_ = _08780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23814" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2;
  assign _08782_ = _08781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23814" *) nand_149_cse;
  assign _08783_ = _08184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23820" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp;
  assign _08784_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23823" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2;
  assign _08785_ = _08784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23824" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _08786_ = _08785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23824" *) IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  assign _08787_ = _08786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23825" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _08788_ = _08787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23826" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2;
  assign _08789_ = _08788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23826" *) nand_147_cse;
  assign _08790_ = _02782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23829" *) _04670_;
  assign _08791_ = _08790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23830" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08792_ = _08791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23830" *) _04669_;
  assign _08793_ = _08792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23831" *) or_4524_cse;
  assign _08794_ = _08793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23831" *) _00063_;
  assign _08795_ = _08794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23831" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp;
  assign _08796_ = _08784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23835" *) _05276_;
  assign _08797_ = _08796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23835" *) IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  assign _08798_ = _08797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23836" *) _05277_;
  assign _08799_ = _08798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23837" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2;
  assign _08800_ = _08799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23837" *) nand_147_cse;
  assign _08801_ = _08203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23843" *) or_4524_cse;
  assign _08802_ = _08801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23843" *) _00063_;
  assign _08803_ = _08802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23843" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp;
  assign _08804_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23846" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2;
  assign _08805_ = _08804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23847" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08806_ = _08805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23847" *) IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  assign _08807_ = _08806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23848" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _08808_ = _08807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23849" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2;
  assign _08809_ = _08808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23849" *) nand_145_cse;
  assign _08810_ = _02783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23852" *) _04668_;
  assign _08811_ = _08810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23853" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08812_ = _08811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23853" *) _04667_;
  assign _08813_ = _08812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23854" *) or_4524_cse;
  assign _08814_ = _08813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23854" *) _00063_;
  assign _08815_ = _08814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23854" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp;
  assign _08816_ = _08804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23858" *) _05278_;
  assign _08817_ = _08816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23858" *) IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  assign _08818_ = _08817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23859" *) _05279_;
  assign _08819_ = _08818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23860" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2;
  assign _08820_ = _08819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23860" *) nand_145_cse;
  assign _08821_ = _08214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23866" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp;
  assign _08822_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23869" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2;
  assign _08823_ = _08822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23870" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08824_ = _08823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23870" *) IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  assign _08825_ = _08824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23871" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _08826_ = _08825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23872" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2;
  assign _08827_ = _08826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23872" *) nand_143_cse;
  assign _08828_ = _02784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23875" *) _04666_;
  assign _08829_ = _08828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23876" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08830_ = _08829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23876" *) _04665_;
  assign _08831_ = _08830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23877" *) or_4524_cse;
  assign _08832_ = _08831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23877" *) _00063_;
  assign _08833_ = _08832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23877" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp;
  assign _08834_ = _08822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23881" *) _05280_;
  assign _08835_ = _08834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23881" *) IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  assign _08836_ = _08835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23882" *) _05281_;
  assign _08837_ = _08836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23883" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2;
  assign _08838_ = _08837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23883" *) nand_143_cse;
  assign _08839_ = _08228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23889" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp;
  assign _08840_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23892" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2;
  assign _08841_ = _08840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23893" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08842_ = _08841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23893" *) IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  assign _08843_ = _08842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23894" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _08844_ = _08843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23895" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2;
  assign _08845_ = _08844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23895" *) nand_141_cse;
  assign _08846_ = _02785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23898" *) _04664_;
  assign _08847_ = _08846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23899" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08848_ = _08847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23899" *) _04663_;
  assign _08849_ = _08848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23900" *) or_4524_cse;
  assign _08850_ = _08849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23900" *) _00063_;
  assign _08851_ = _08850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23900" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp;
  assign _08852_ = _08840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23904" *) _05282_;
  assign _08853_ = _08852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23904" *) IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  assign _08854_ = _08853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23905" *) _05283_;
  assign _08855_ = _08854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23906" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2;
  assign _08856_ = _08855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23906" *) nand_141_cse;
  assign _08857_ = _08247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23912" *) or_4524_cse;
  assign _08858_ = _08857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23912" *) _00063_;
  assign _08859_ = _08858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23912" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp;
  assign _08860_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23915" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2;
  assign _08861_ = _08860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23916" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _08862_ = _08861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23916" *) IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  assign _08863_ = _08862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23917" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _08864_ = _08863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23918" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2;
  assign _08865_ = _08864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23918" *) nand_139_cse;
  assign _08866_ = _02786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23921" *) _04662_;
  assign _08867_ = _08866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23922" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08868_ = _08867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23922" *) _04661_;
  assign _08869_ = _08868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23923" *) or_4524_cse;
  assign _08870_ = _08869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23923" *) _00063_;
  assign _08871_ = _08870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23923" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp;
  assign _08872_ = _08860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23927" *) _05284_;
  assign _08873_ = _08872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23927" *) IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  assign _08874_ = _08873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23928" *) _05285_;
  assign _08875_ = _08874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23929" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2;
  assign _08876_ = _08875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23929" *) nand_139_cse;
  assign _08877_ = _08258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23935" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp;
  assign _08878_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23938" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2;
  assign _08879_ = _08878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23939" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08880_ = _08879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23939" *) IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  assign _08881_ = _08880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23940" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _08882_ = _08881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23941" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2;
  assign _08883_ = _08882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23941" *) nand_137_cse;
  assign _08884_ = _02787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23944" *) _04660_;
  assign _08885_ = _08884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23945" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08886_ = _08885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23945" *) _04659_;
  assign _08887_ = _08886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23946" *) or_4524_cse;
  assign _08888_ = _08887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23946" *) _00063_;
  assign _08889_ = _08888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23946" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp;
  assign _08890_ = _08878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23950" *) _05286_;
  assign _08891_ = _08890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23950" *) IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  assign _08892_ = _08891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23951" *) _05287_;
  assign _08893_ = _08892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23952" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2;
  assign _08894_ = _08893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23952" *) nand_137_cse;
  assign _08895_ = _08272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23958" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp;
  assign _08896_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23961" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2;
  assign _08897_ = _08896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23962" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _08898_ = _08897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23962" *) IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  assign _08899_ = _08898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23963" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _08900_ = _08899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23964" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2;
  assign _08901_ = _08900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23964" *) nand_135_cse;
  assign _08902_ = _02788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23967" *) _04658_;
  assign _08903_ = _08902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23968" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08904_ = _08903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23968" *) _04657_;
  assign _08905_ = _08904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23969" *) or_4524_cse;
  assign _08906_ = _08905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23969" *) _00063_;
  assign _08907_ = _08906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23969" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp;
  assign _08908_ = _08896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23973" *) _05288_;
  assign _08909_ = _08908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23973" *) IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  assign _08910_ = _08909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23974" *) _05289_;
  assign _08911_ = _08910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23975" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2;
  assign _08912_ = _08911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23975" *) nand_135_cse;
  assign _08913_ = _08286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23981" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp;
  assign _08914_ = or_23_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23984" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2;
  assign _08915_ = _08914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23985" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2;
  assign _08916_ = _08915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23985" *) IsNaN_8U_23U_land_lpi_1_dfm_3;
  assign _08917_ = _08916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23986" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2;
  assign _08918_ = _08917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23987" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2;
  assign _08919_ = _08918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23987" *) nand_133_cse;
  assign _08920_ = _02789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23990" *) _04656_;
  assign _08921_ = _08920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23991" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7];
  assign _08922_ = _08921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23991" *) _04655_;
  assign _08923_ = _08922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23992" *) or_4524_cse;
  assign _08924_ = _08923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23992" *) _00063_;
  assign _08925_ = _08924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23992" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp;
  assign _08926_ = _08914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23996" *) _05290_;
  assign _08927_ = _08926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23996" *) IsNaN_8U_23U_land_lpi_1_dfm_3;
  assign _08928_ = _08927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23997" *) _05291_;
  assign _08929_ = _08928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23998" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2;
  assign _08930_ = _08929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:23998" *) nand_133_cse;
  assign _08931_ = _04656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24003" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7];
  assign _08932_ = _08931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24003" *) _04655_;
  assign _08933_ = _04658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24008" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08934_ = _08933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24008" *) _04657_;
  assign _08935_ = _04660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24013" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08936_ = _08935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24013" *) _04659_;
  assign _08937_ = _04662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24018" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08938_ = _08937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24018" *) _04661_;
  assign _08939_ = _04664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24023" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08940_ = _08939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24023" *) _04663_;
  assign _08941_ = _04666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24028" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08942_ = _08941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24028" *) _04665_;
  assign _08943_ = _04668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24035" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08944_ = _08943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24035" *) _04667_;
  assign _08945_ = _04185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *) cfg_proc_precision_1_sva_st_64[0];
  assign _08946_ = _08945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24038" *) _05292_;
  assign _08947_ = _04670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24043" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08948_ = _08947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24043" *) _04669_;
  assign _08949_ = _04672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24048" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign _08950_ = _08949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24048" *) _04671_;
  assign _08951_ = _04674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24053" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08952_ = _08951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24053" *) _04673_;
  assign _08953_ = _04676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24060" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08954_ = _08953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24060" *) _04675_;
  assign _08955_ = _08945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24063" *) _05293_;
  assign _08956_ = _04678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24068" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08957_ = _08956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24068" *) _04677_;
  assign _08958_ = _04680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24073" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign _08959_ = _08958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24073" *) _04679_;
  assign _08960_ = _04682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24078" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08961_ = _08960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24078" *) _04681_;
  assign _08962_ = _04684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24083" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign _08963_ = _08962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24083" *) _04683_;
  assign _08964_ = or_17_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24088" *) _04685_;
  assign or_724_nl = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24123" *) _05294_;
  assign or_733_nl = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24125" *) _05295_;
  assign or_1118_nl = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24127" *) _05296_;
  assign or_1134_nl = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24129" *) _04572_;
  assign or_1145_nl = cfg_proc_precision_1_sva_st_101[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24132" *) _05297_;
  assign or_236_nl = or_2251_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24226" *) _05294_;
  assign or_263_nl = cfg_out_precision_1_sva_st_154[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24229" *) _05298_;
  assign or_270_nl = or_2251_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24231" *) _04572_;
  assign or_275_nl = or_2251_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24233" *) _05296_;
  assign _08965_ = _02801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02864_;
  assign _08966_ = _02802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02865_;
  assign _08967_ = _02803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02866_;
  assign _08968_ = _02804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02867_;
  assign _08969_ = _02805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02868_;
  assign _08970_ = _02806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02869_;
  assign _08971_ = _02807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02870_;
  assign _08972_ = _02808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02871_;
  assign _08973_ = _02809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02872_;
  assign _08974_ = _02810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02873_;
  assign _08975_ = _02811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02874_;
  assign _08976_ = _02812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02875_;
  assign _08977_ = _02813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02876_;
  assign _08978_ = _02814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02877_;
  assign _08979_ = _02815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02878_;
  assign _08980_ = _02816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02879_;
  assign _08981_ = _02817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02880_;
  assign _08982_ = _02818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02881_;
  assign _08983_ = _02819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02882_;
  assign _08984_ = _02820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02883_;
  assign _08985_ = _02821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02884_;
  assign _08986_ = _02822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02885_;
  assign _08987_ = _02823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02886_;
  assign _08988_ = _02824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02887_;
  assign _08989_ = _02825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02888_;
  assign _08990_ = _02826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02889_;
  assign _08991_ = _02827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02890_;
  assign _08992_ = _02828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02891_;
  assign _08993_ = _02829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02892_;
  assign _08994_ = _02830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02893_;
  assign _08995_ = _02831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02894_;
  assign _08996_ = _02832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02895_;
  assign _08997_ = _02833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02896_;
  assign _08998_ = _02834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02897_;
  assign _08999_ = _02835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02898_;
  assign _09000_ = _02836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02899_;
  assign _09001_ = _02837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02900_;
  assign _09002_ = _02838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02901_;
  assign _09003_ = _02839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02902_;
  assign _09004_ = _02840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02903_;
  assign _09005_ = _02841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02904_;
  assign _09006_ = _02842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02905_;
  assign _09007_ = _02843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02906_;
  assign _09008_ = _02844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02907_;
  assign _09009_ = _02845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02908_;
  assign _09010_ = _02846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02909_;
  assign _09011_ = _02847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02910_;
  assign _09012_ = _02848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02911_;
  assign _09013_ = _02849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02912_;
  assign _09014_ = _02850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02913_;
  assign _09015_ = _02851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02914_;
  assign _09016_ = _02852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02915_;
  assign _09017_ = _02853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02916_;
  assign _09018_ = _02854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02917_;
  assign _09019_ = _02855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02918_;
  assign _09020_ = _02856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02919_;
  assign _09021_ = _02857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02920_;
  assign _09022_ = _02858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02921_;
  assign _09023_ = _02859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02922_;
  assign _09024_ = _02860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02923_;
  assign _09025_ = _02861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02924_;
  assign _09026_ = _02862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02925_;
  assign _09027_ = _02863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24252" *) _02926_;
  assign _09028_ = _08965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02927_;
  assign _09029_ = _08966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02928_;
  assign _09030_ = _08967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02929_;
  assign _09031_ = _08968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02930_;
  assign _09032_ = _08969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02931_;
  assign _09033_ = _08970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02932_;
  assign _09034_ = _08971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02933_;
  assign _09035_ = _08972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02934_;
  assign _09036_ = _08973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02935_;
  assign _09037_ = _08974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02936_;
  assign _09038_ = _08975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02937_;
  assign _09039_ = _08976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02938_;
  assign _09040_ = _08977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02939_;
  assign _09041_ = _08978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02940_;
  assign _09042_ = _08979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02941_;
  assign _09043_ = _08980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02942_;
  assign _09044_ = _08981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02943_;
  assign _09045_ = _08982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02944_;
  assign _09046_ = _08983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02945_;
  assign _09047_ = _08984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02946_;
  assign _09048_ = _08985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02947_;
  assign _09049_ = _08986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02948_;
  assign _09050_ = _08987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02949_;
  assign _09051_ = _08988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02950_;
  assign _09052_ = _08989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02951_;
  assign _09053_ = _08990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02952_;
  assign _09054_ = _08991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02953_;
  assign _09055_ = _08992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02954_;
  assign _09056_ = _08993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02955_;
  assign _09057_ = _08994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02956_;
  assign _09058_ = _08995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02957_;
  assign chn_odata_data_13_0_lpi_1_dfm_1_mx0w0 = _08996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02958_;
  assign cvt_else_mux1h_10_nl = _08997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02959_;
  assign cvt_else_mux1h_8_nl = _08998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02960_;
  assign cvt_else_mux1h_29_nl = _08999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02961_;
  assign cvt_else_mux1h_27_nl = _09000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02962_;
  assign cvt_else_mux1h_48_nl = _09001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02963_;
  assign cvt_else_mux1h_46_nl = _09002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02964_;
  assign cvt_else_mux1h_67_nl = _09003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02965_;
  assign cvt_else_mux1h_65_nl = _09004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02966_;
  assign cvt_else_mux1h_86_nl = _09005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02967_;
  assign cvt_else_mux1h_84_nl = _09006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02968_;
  assign cvt_else_mux1h_105_nl = _09007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02969_;
  assign cvt_else_mux1h_103_nl = _09008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02970_;
  assign cvt_else_mux1h_124_nl = _09009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02971_;
  assign cvt_else_mux1h_122_nl = _09010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02972_;
  assign cvt_else_mux1h_143_nl = _09011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02973_;
  assign cvt_else_mux1h_141_nl = _09012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02974_;
  assign cvt_else_mux1h_162_nl = _09013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02975_;
  assign cvt_else_mux1h_160_nl = _09014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02976_;
  assign cvt_else_mux1h_181_nl = _09015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02977_;
  assign cvt_else_mux1h_179_nl = _09016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02978_;
  assign cvt_else_mux1h_200_nl = _09017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02979_;
  assign cvt_else_mux1h_198_nl = _09018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02980_;
  assign cvt_else_mux1h_219_nl = _09019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02981_;
  assign cvt_else_mux1h_217_nl = _09020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02982_;
  assign cvt_else_mux1h_238_nl = _09021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02983_;
  assign cvt_else_mux1h_236_nl = _09022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02984_;
  assign cvt_else_mux1h_255_nl = _09023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02985_;
  assign cvt_else_mux1h_276_nl = _09024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02986_;
  assign cvt_else_mux1h_274_nl = _09025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02987_;
  assign cvt_else_mux1h_295_nl = _09026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02988_;
  assign cvt_else_mux1h_292_nl = _09027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24253" *) _02989_;
  assign _09059_ = _02990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03006_;
  assign _09060_ = _02991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03007_;
  assign _09061_ = _02992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03008_;
  assign _09062_ = _02993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03009_;
  assign _09063_ = _02994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03010_;
  assign _09064_ = _02995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03011_;
  assign _09065_ = _02996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03012_;
  assign _09066_ = _02997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03013_;
  assign _09067_ = _02998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03014_;
  assign _09068_ = _02999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03015_;
  assign _09069_ = _03000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03016_;
  assign _09070_ = _03001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03017_;
  assign _09071_ = _03002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03018_;
  assign _09072_ = _03003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03019_;
  assign _09073_ = _03004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03020_;
  assign _09074_ = _03005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24267" *) _03021_;
  assign _09075_ = _09059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03022_;
  assign _09076_ = _09060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03023_;
  assign _09077_ = _09061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03024_;
  assign _09078_ = _09062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03025_;
  assign _09079_ = _09063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03026_;
  assign _09080_ = _09064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03027_;
  assign _09081_ = _09065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03028_;
  assign _09082_ = _09066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03029_;
  assign _09083_ = _09067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03030_;
  assign _09084_ = _09068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03031_;
  assign _09085_ = _09069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03032_;
  assign _09086_ = _09070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03033_;
  assign _09087_ = _09071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03034_;
  assign _09088_ = _09072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03035_;
  assign _09089_ = _09073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03036_;
  assign _09090_ = _09074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24268" *) _03037_;
  assign _09091_ = _09075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03038_;
  assign _09092_ = _09076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03039_;
  assign _09093_ = _09077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03040_;
  assign _09094_ = _09078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03041_;
  assign _09095_ = _09079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03042_;
  assign _09096_ = _09080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03043_;
  assign _09097_ = _09081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03044_;
  assign _09098_ = _09082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03045_;
  assign _09099_ = _09083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03046_;
  assign _09100_ = _09084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03047_;
  assign _09101_ = _09085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03048_;
  assign _09102_ = _09086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03049_;
  assign _09103_ = _09087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03050_;
  assign _09104_ = _09088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03051_;
  assign _09105_ = _09089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03052_;
  assign _09106_ = _09090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24269" *) _03053_;
  assign _09107_ = _09091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03054_;
  assign _09108_ = _09092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03055_;
  assign _09109_ = _09093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03056_;
  assign _09110_ = _09094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03057_;
  assign _09111_ = _09095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03058_;
  assign _09112_ = _09096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03059_;
  assign _09113_ = _09097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03060_;
  assign _09114_ = _09098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03061_;
  assign _09115_ = _09099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03062_;
  assign _09116_ = _09100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03063_;
  assign _09117_ = _09101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03064_;
  assign _09118_ = _09102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03065_;
  assign _09119_ = _09103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03066_;
  assign _09120_ = _09104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03067_;
  assign _09121_ = _09105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03068_;
  assign _09122_ = _09106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24270" *) _03069_;
  assign _09123_ = _03070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03098_;
  assign _09124_ = _03071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03099_;
  assign _09125_ = _03072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03100_;
  assign _09126_ = _03073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03101_;
  assign _09127_ = _03074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03102_;
  assign _09128_ = _03075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03103_;
  assign _09129_ = _03076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03104_;
  assign _09130_ = _03077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03105_;
  assign _09131_ = _03078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03106_;
  assign _09132_ = _03079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03107_;
  assign _09133_ = _03080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03108_;
  assign _09134_ = _03081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03109_;
  assign _09135_ = _03082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03110_;
  assign _09136_ = _03083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03111_;
  assign _09137_ = _03084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03112_;
  assign _09138_ = _03085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03113_;
  assign _09139_ = _03086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03114_;
  assign _09140_ = _03087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03115_;
  assign _09141_ = _03088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03116_;
  assign _09142_ = _03089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03117_;
  assign _09143_ = _03090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03118_;
  assign _09144_ = _03091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03119_;
  assign _09145_ = _03092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03120_;
  assign _09146_ = _03093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03121_;
  assign _09147_ = _03094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03122_;
  assign _09148_ = _03095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03123_;
  assign _09149_ = _03096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03124_;
  assign _09150_ = _03097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24282" *) _03125_;
  assign _09151_ = _09123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03126_;
  assign _09152_ = _09124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03127_;
  assign _09153_ = _09125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03128_;
  assign _09154_ = _09126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03129_;
  assign _09155_ = _09127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03130_;
  assign _09156_ = _09128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03131_;
  assign _09157_ = _09129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03132_;
  assign _09158_ = _09130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03133_;
  assign _09159_ = _09131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03134_;
  assign _09160_ = _09132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03135_;
  assign _09161_ = _09133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03136_;
  assign _09162_ = _09134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03137_;
  assign _09163_ = _09135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03138_;
  assign _09164_ = _09136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03139_;
  assign _09165_ = _09137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03140_;
  assign _09166_ = _09138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03141_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt = _09139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03142_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt = _09140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03143_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt = _09141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03144_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt = _09142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03145_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt = _09143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03146_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt = _09144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03147_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt = _09145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03148_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt = _09146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03149_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt = _09147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03150_;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt = _09148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03151_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt = _09149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03152_;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt = _09150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24283" *) _03153_;
  assign _09167_ = _03154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *) _03157_;
  assign _09168_ = _03155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *) _03158_;
  assign _09169_ = _03156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24298" *) _03159_;
  assign _09170_ = _09167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *) _03160_;
  assign _09171_ = _09168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *) _03161_;
  assign _09172_ = _09169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24299" *) _03162_;
  assign _09173_ = _09170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *) _03163_;
  assign _09174_ = _09171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *) _03164_;
  assign _09175_ = _09172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24300" *) _03165_;
  assign _09176_ = _09173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *) _03166_;
  assign _09177_ = _09174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *) _03167_;
  assign _09178_ = _09175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24301" *) _03168_;
  assign _09179_ = _09176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *) _03169_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt = _09177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *) _03170_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_nl = _09178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24302" *) _03171_;
  assign _09180_ = _03172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03185_;
  assign _09181_ = _03173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03186_;
  assign _09182_ = _03174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03187_;
  assign _09183_ = _03175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03188_;
  assign _09184_ = _03176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03189_;
  assign _09185_ = _03177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03190_;
  assign _09186_ = _03178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03191_;
  assign _09187_ = _03179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03192_;
  assign _09188_ = _03180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03193_;
  assign _09189_ = _03181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03194_;
  assign _09190_ = _03182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03195_;
  assign _09191_ = _03183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03196_;
  assign _09192_ = _03184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24318" *) _03197_;
  assign _09193_ = _09180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03198_;
  assign _09194_ = _09181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03199_;
  assign _09195_ = _09182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03200_;
  assign _09196_ = _09183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03201_;
  assign _09197_ = _09184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03202_;
  assign _09198_ = _09185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03203_;
  assign _09199_ = _09186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03204_;
  assign _09200_ = _09187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03205_;
  assign _09201_ = _09188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03206_;
  assign _09202_ = _09189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03207_;
  assign _09203_ = _09190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03208_;
  assign _09204_ = _09191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03209_;
  assign _09205_ = _09192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24319" *) _03210_;
  assign _09206_ = _09193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03211_;
  assign _09207_ = _09194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03212_;
  assign _09208_ = _09195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03213_;
  assign _09209_ = _09196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03214_;
  assign _09210_ = _09197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03215_;
  assign _09211_ = _09198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03216_;
  assign _09212_ = _09199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03217_;
  assign _09213_ = _09200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03218_;
  assign _09214_ = _09201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03219_;
  assign _09215_ = _09202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03220_;
  assign _09216_ = _09203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03221_;
  assign _09217_ = _09204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03222_;
  assign _09218_ = _09205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24320" *) _03223_;
  assign _09219_ = _09206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03224_;
  assign _09220_ = _09207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03225_;
  assign _09221_ = _09208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03226_;
  assign _09222_ = _09209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03227_;
  assign _09223_ = _09210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03228_;
  assign _09224_ = _09211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03229_;
  assign _09225_ = _09212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03230_;
  assign _09226_ = _09213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03231_;
  assign _09227_ = _09214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03232_;
  assign _09228_ = _09215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03233_;
  assign _09229_ = _09216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03234_;
  assign _09230_ = _09217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03235_;
  assign _09231_ = _09218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24321" *) _03236_;
  assign _09232_ = _09219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03237_;
  assign _09233_ = _09220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03238_;
  assign _09234_ = _09221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03239_;
  assign _09235_ = _09222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03240_;
  assign _09236_ = _09223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03241_;
  assign _09237_ = _09224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03242_;
  assign _09238_ = _09225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03243_;
  assign _09239_ = _09226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03244_;
  assign _09240_ = _09227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03245_;
  assign _09241_ = _09228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03246_;
  assign _09242_ = _09229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03247_;
  assign _09243_ = _09230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03248_;
  assign _09244_ = _09231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24322" *) _03249_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt = _09232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03250_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt = _09233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03251_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt = _09234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03252_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt = _09235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03253_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt = _09236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03254_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt = _09237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03255_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt = _09238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03256_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt = _09239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03257_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt = _09240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03258_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt = _09241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03259_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt = _09242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03260_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt = _09243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03261_;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt = _09244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24323" *) _03262_;
  assign _09245_ = _03263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24335" *) _03264_;
  assign chn_idata_data_mux1h_65_rgt = _09245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24336" *) _03265_;
  assign _09246_ = _03266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03282_;
  assign _09247_ = _03267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03283_;
  assign _09248_ = _03268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03284_;
  assign _09249_ = _03269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03285_;
  assign _09250_ = _03270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03286_;
  assign _09251_ = _03271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03287_;
  assign _09252_ = _03272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03288_;
  assign _09253_ = _03273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03289_;
  assign _09254_ = _03274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03290_;
  assign _09255_ = _03275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03291_;
  assign _09256_ = _03276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03292_;
  assign _09257_ = _03277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03293_;
  assign _09258_ = _03278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03294_;
  assign _09259_ = _03279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03295_;
  assign _09260_ = _03280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03296_;
  assign _09261_ = _03281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24349" *) _03297_;
  assign _09262_ = _09246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03298_;
  assign _09263_ = _09247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03299_;
  assign _09264_ = _09248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03300_;
  assign _09265_ = _09249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03301_;
  assign _09266_ = _09250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03302_;
  assign _09267_ = _09251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03303_;
  assign _09268_ = _09252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03304_;
  assign _09269_ = _09253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03305_;
  assign _09270_ = _09254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03306_;
  assign _09271_ = _09255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03307_;
  assign _09272_ = _09256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03308_;
  assign _09273_ = _09257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03309_;
  assign _09274_ = _09258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03310_;
  assign _09275_ = _09259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03311_;
  assign _09276_ = _09260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03312_;
  assign _09277_ = _09261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24350" *) _03313_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl = _09262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03314_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_1_nl = _09263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03315_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_2_nl = _09264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03316_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_3_nl = _09265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03317_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_4_nl = _09266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03318_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_5_nl = _09267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03319_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_6_nl = _09268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03320_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_7_nl = _09269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03321_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_8_nl = _09270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03322_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_9_nl = _09271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03323_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_10_nl = _09272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03324_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_11_nl = _09273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03325_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_12_nl = _09274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03326_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_13_nl = _09275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03327_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_14_nl = _09276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03328_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_15_nl = _09277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24351" *) _03329_;
  assign _09278_ = _03330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03346_;
  assign _09279_ = _03331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03347_;
  assign _09280_ = _03332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03348_;
  assign _09281_ = _03333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03349_;
  assign _09282_ = _03334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03350_;
  assign _09283_ = _03335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03351_;
  assign _09284_ = _03336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03352_;
  assign _09285_ = _03337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03353_;
  assign _09286_ = _03338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03354_;
  assign _09287_ = _03339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03355_;
  assign _09288_ = _03340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03356_;
  assign _09289_ = _03341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03357_;
  assign _09290_ = _03342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03358_;
  assign _09291_ = _03343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03359_;
  assign _09292_ = _03344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03360_;
  assign _09293_ = _03345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24366" *) _03361_;
  assign _09294_ = _09278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03362_;
  assign _09295_ = _09279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03363_;
  assign _09296_ = _09280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03364_;
  assign _09297_ = _09281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03365_;
  assign _09298_ = _09282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03366_;
  assign _09299_ = _09283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03367_;
  assign _09300_ = _09284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03368_;
  assign _09301_ = _09285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03369_;
  assign _09302_ = _09286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03370_;
  assign _09303_ = _09287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03371_;
  assign _09304_ = _09288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03372_;
  assign _09305_ = _09289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03373_;
  assign _09306_ = _09290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03374_;
  assign _09307_ = _09291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03375_;
  assign _09308_ = _09292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03376_;
  assign _09309_ = _09293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24367" *) _03377_;
  assign _09310_ = _09294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03378_;
  assign _09311_ = _09295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03379_;
  assign _09312_ = _09296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03380_;
  assign _09313_ = _09297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03381_;
  assign _09314_ = _09298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03382_;
  assign _09315_ = _09299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03383_;
  assign _09316_ = _09300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03384_;
  assign _09317_ = _09301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03385_;
  assign _09318_ = _09302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03386_;
  assign _09319_ = _09303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03387_;
  assign _09320_ = _09304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03388_;
  assign _09321_ = _09305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03389_;
  assign _09322_ = _09306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03390_;
  assign _09323_ = _09307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03391_;
  assign _09324_ = _09308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03392_;
  assign _09325_ = _09309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24368" *) _03393_;
  assign _09326_ = _09310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03394_;
  assign _09327_ = _09311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03395_;
  assign _09328_ = _09312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03396_;
  assign _09329_ = _09313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03397_;
  assign _09330_ = _09314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03398_;
  assign _09331_ = _09315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03399_;
  assign _09332_ = _09316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03400_;
  assign _09333_ = _09317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03401_;
  assign _09334_ = _09318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03402_;
  assign _09335_ = _09319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03403_;
  assign _09336_ = _09320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03404_;
  assign _09337_ = _09321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03405_;
  assign _09338_ = _09322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03406_;
  assign _09339_ = _09323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03407_;
  assign _09340_ = _09324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03408_;
  assign _09341_ = _09325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24369" *) _03409_;
  assign _09342_ = _09326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03410_;
  assign _09343_ = _09327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03411_;
  assign _09344_ = _09328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03412_;
  assign _09345_ = _09329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03413_;
  assign _09346_ = _09330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03414_;
  assign _09347_ = _09331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03415_;
  assign _09348_ = _09332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03416_;
  assign _09349_ = _09333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03417_;
  assign _09350_ = _09334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03418_;
  assign _09351_ = _09335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03419_;
  assign _09352_ = _09336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03420_;
  assign _09353_ = _09337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03421_;
  assign _09354_ = _09338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03422_;
  assign _09355_ = _09339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03423_;
  assign _09356_ = _09340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03424_;
  assign _09357_ = _09341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24370" *) _03425_;
  assign _09358_ = _03426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03442_;
  assign _09359_ = _03427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03443_;
  assign _09360_ = _03428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03444_;
  assign _09361_ = _03429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03445_;
  assign _09362_ = _03430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03446_;
  assign _09363_ = _03431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03447_;
  assign _09364_ = _03432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03448_;
  assign _09365_ = _03433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03449_;
  assign _09366_ = _03434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03450_;
  assign _09367_ = _03435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03451_;
  assign _09368_ = _03436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03452_;
  assign _09369_ = _03437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03453_;
  assign _09370_ = _03438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03454_;
  assign _09371_ = _03439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03455_;
  assign _09372_ = _03440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03456_;
  assign _09373_ = _03441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24382" *) _03457_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm = _09358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03458_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm = _09359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03459_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm = _09360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03460_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm = _09361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03461_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm = _09362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03462_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm = _09363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03463_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm = _09364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03464_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm = _09365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03465_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm = _09366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03466_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm = _09367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03467_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm = _09368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03468_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm = _09369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03469_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm = _09370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03470_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm = _09371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03471_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm = _09372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03472_;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm = _09373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24383" *) _03473_;
  assign _09374_ = _03474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03490_;
  assign _09375_ = _03475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03491_;
  assign _09376_ = _03476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03492_;
  assign _09377_ = _03477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03493_;
  assign _09378_ = _03478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03494_;
  assign _09379_ = _03479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03495_;
  assign _09380_ = _03480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03496_;
  assign _09381_ = _03481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03497_;
  assign _09382_ = _03482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03498_;
  assign _09383_ = _03483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03499_;
  assign _09384_ = _03484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03500_;
  assign _09385_ = _03485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03501_;
  assign _09386_ = _03486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03502_;
  assign _09387_ = _03487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03503_;
  assign _09388_ = _03488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03504_;
  assign _03863_ = _03489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24395" *) _03505_;
  assign IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1 = _09374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03506_;
  assign IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1 = _09375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03507_;
  assign IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1 = _09376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03508_;
  assign IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1 = _09377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03509_;
  assign IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1 = _09378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03510_;
  assign IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1 = _09379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03511_;
  assign IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1 = _09380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03512_;
  assign IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1 = _09381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03513_;
  assign IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1 = _09382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03514_;
  assign IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1 = _09383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03515_;
  assign IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1 = _09384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03516_;
  assign IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1 = _09385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03517_;
  assign IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1 = _09386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03518_;
  assign IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1 = _09387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03519_;
  assign IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1 = _09388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) _03520_;
  assign IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1 = _03863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24396" *) { _03846_[6:2], _03521_ };
  assign _09389_ = _03522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24409" *) _03523_;
  assign _09390_ = _09389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24410" *) _03524_;
  assign _09391_ = _09390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24411" *) _03525_;
  assign _09392_ = _03526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03541_;
  assign _09393_ = _03527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03542_;
  assign _09394_ = _03528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03543_;
  assign _09395_ = _03529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03544_;
  assign _09396_ = _03530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03545_;
  assign _09397_ = _03531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03546_;
  assign _09398_ = _03532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03547_;
  assign _09399_ = _03533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03548_;
  assign _09400_ = _03534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03549_;
  assign _09401_ = _03535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03550_;
  assign _09402_ = _03536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03551_;
  assign _09403_ = _03537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03552_;
  assign _09404_ = _03538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03553_;
  assign _09405_ = _03539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03554_;
  assign _09406_ = _03540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24425" *) _03555_;
  assign _09407_ = _09392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03556_;
  assign _09408_ = _09393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03557_;
  assign _09409_ = _09394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03558_;
  assign _09410_ = _09395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03559_;
  assign _09411_ = _09396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03560_;
  assign _09412_ = _09397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03561_;
  assign _09413_ = _09398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03562_;
  assign _09414_ = _09399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03563_;
  assign _09415_ = _09400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03564_;
  assign _09416_ = _09401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03565_;
  assign _09417_ = _09402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03566_;
  assign _09418_ = _09403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03567_;
  assign _09419_ = _09404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03568_;
  assign _09420_ = _09405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03569_;
  assign _09421_ = _09406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24426" *) _03570_;
  assign _09422_ = _09407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03571_;
  assign _09423_ = _09408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03572_;
  assign _09424_ = _09409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03573_;
  assign _09425_ = _09410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03574_;
  assign _09426_ = _09411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03575_;
  assign _09427_ = _09412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03576_;
  assign _09428_ = _09413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03577_;
  assign _09429_ = _09414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03578_;
  assign _09430_ = _09415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03579_;
  assign _09431_ = _09416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03580_;
  assign _09432_ = _09417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03581_;
  assign _09433_ = _09418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03582_;
  assign _09434_ = _09419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03583_;
  assign _09435_ = _09420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03584_;
  assign _09436_ = _09421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24427" *) _03585_;
  assign _09437_ = _09422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03586_;
  assign _09438_ = _09423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03587_;
  assign _09439_ = _09424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03588_;
  assign _09440_ = _09425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03589_;
  assign _09441_ = _09426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03590_;
  assign _09442_ = _09427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03591_;
  assign _09443_ = _09428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03592_;
  assign _09444_ = _09429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03593_;
  assign _09445_ = _09430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03594_;
  assign _09446_ = _09431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03595_;
  assign _09447_ = _09432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03596_;
  assign _09448_ = _09433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03597_;
  assign _09449_ = _09434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03598_;
  assign _09450_ = _09435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03599_;
  assign _09451_ = _09436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24428" *) _03600_;
  assign cvt_or_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8773" *) _03602_;
  assign _09452_ = _07546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8776" *) _04172_;
  assign cvt_or_2_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8779" *) _03605_;
  assign cvt_or_6_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8781" *) _03607_;
  assign cvt_or_10_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8783" *) _03609_;
  assign cvt_or_12_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8785" *) _03611_;
  assign cvt_or_14_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8786" *) _03612_;
  assign cvt_or_18_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8788" *) _03614_;
  assign cvt_or_20_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8790" *) _03616_;
  assign cvt_or_22_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8792" *) _03618_;
  assign cvt_or_24_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8794" *) _03620_;
  assign cvt_or_26_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8796" *) _03622_;
  assign _09453_ = _05300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8799" *) _04566_;
  assign _09454_ = _09453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8799" *) cfg_mode_eql_1_sva_6;
  assign cvt_or_28_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8802" *) _03625_;
  assign cvt_or_30_cse = cvt_asn_319 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8805" *) _03627_;
  assign _09455_ = _03629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8807" *) and_dcpl_98;
  assign _09456_ = _03631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8809" *) and_dcpl_102;
  assign _09457_ = and_550_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8818" *) IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1;
  assign or_306_cse = _05426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8824" *) or_4550_cse;
  assign _09458_ = nor_2040_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8836" *) _04006_;
  assign _09459_ = _09458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8837" *) _04185_;
  assign or_303_cse = _09459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8837" *) or_4550_cse;
  assign _09460_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8861" *) _05317_;
  assign or_419_cse = or_513_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8865" *) or_961_nl;
  assign IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse = and_dcpl_204 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8869" *) and_dcpl_4;
  assign _09461_ = _03634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8872" *) and_dcpl_209;
  assign IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse = and_676_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8878" *) and_685_rgt;
  assign _09462_ = or_961_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8879" *) _04581_;
  assign _09463_ = _03637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8883" *) and_dcpl_217;
  assign _09464_ = _08302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8888" *) _00064_;
  assign _09465_ = _03640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8894" *) and_dcpl_224;
  assign _09466_ = or_961_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8897" *) _04588_;
  assign _09467_ = nor_tmp_636 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8898" *) or_2251_nl;
  assign or_3063_cse = _09467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8898" *) or_dcpl_15;
  assign or_4559_cse = nor_2150_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8912" *) cfg_out_precision_1_sva_st_154[0];
  assign _09468_ = cfg_out_precision_1_sva_st_154[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8913" *) nor_1314_nl;
  assign _09469_ = nor_tmp_636 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8923" *) cfg_out_precision_1_sva_st_154[0];
  assign or_3070_nl = _09469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8923" *) not_tmp_2254;
  assign _09470_ = cfg_proc_precision_1_sva_st_64[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8932" *) nor_2150_cse;
  assign _09471_ = mux_2179_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8947" *) nor_2040_cse;
  assign or_4536_cse = IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8953" *) cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign _09472_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8954" *) _05322_;
  assign or_4535_cse = IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8963" *) cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2;
  assign _09473_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8964" *) _05167_;
  assign _09474_ = or_961_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8966" *) _05323_;
  assign _09475_ = _03654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8977" *) and_dcpl_301;
  assign _09476_ = cfg_proc_precision_1_sva_st_64[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8979" *) _05325_;
  assign _09477_ = cfg_out_precision_1_sva_st_154[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9007" *) _05326_;
  assign _09478_ = mux_2196_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9011" *) nor_2040_cse;
  assign _09479_ = or_961_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9025" *) _05112_;
  assign _09480_ = cfg_out_precision_1_sva_st_154[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9029" *) main_stage_v_2;
  assign or_3170_nl = _09480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9029" *) not_tmp_270;
  assign or_4348_nl = mux_1799_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9037" *) fsm_output[0];
  assign _09481_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9045" *) _05329_;
  assign or_3196_nl = cfg_out_precision_1_sva_st_149[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9051" *) _05330_;
  assign _09482_ = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9061" *) or_2251_nl;
  assign or_3220_nl = _09482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9062" *) or_dcpl_15;
  assign _09483_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9071" *) _05331_;
  assign _09484_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9073" *) _04630_;
  assign _09485_ = and_dcpl_407 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9081" *) and_dcpl_409;
  assign _09486_ = _09485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9081" *) and_dcpl_411;
  assign _09487_ = _05123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9082" *) or_309_cse;
  assign _09488_ = or_300_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9087" *) _00058_;
  assign _09489_ = _09488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9087" *) cfg_mode_eql_1_sva_5;
  assign _09490_ = _05123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9090" *) cfg_out_precision_1_sva_st_149[1];
  assign _09491_ = _09490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9090" *) cfg_proc_precision_1_sva_st_65[0];
  assign _09492_ = _09491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9090" *) nand_219_cse;
  assign or_1176_cse = or_1157_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9093" *) cfg_mode_eql_1_sva_6;
  assign _09493_ = _09488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9096" *) cvt_unequal_tmp_20;
  assign _09494_ = _09493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9096" *) cfg_mode_eql_1_sva_5;
  assign _09495_ = or_1157_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9099" *) _04631_;
  assign _09496_ = _09495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9099" *) cvt_unequal_tmp_21;
  assign _09497_ = _09496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9099" *) cfg_mode_eql_1_sva_6;
  assign IsNaN_5U_10U_aelse_or_cse = _03675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9103" *) and_dcpl_424;
  assign or_4709_cse = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9110" *) nor_2285_cse;
  assign _09498_ = or_dcpl_151 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9128" *) cfg_out_precision_1_sva_st_113[0];
  assign _09499_ = nor_213_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9133" *) cfg_out_precision_1_sva_6[0];
  assign _09500_ = _09499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9133" *) nand_207_cse;
  assign IsNaN_5U_10U_aelse_or_1_cse = and_dcpl_408 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9147" *) and_dcpl_420;
  assign _09501_ = cfg_proc_precision_1_sva_st_65[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9167" *) _05336_;
  assign _09502_ = _04691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9169" *) or_4862_cse;
  assign or_4718_nl = _05337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9170" *) cvt_unequal_tmp_20;
  assign _09503_ = and_2360_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9173" *) cvt_unequal_tmp_20;
  assign _09504_ = _09503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9173" *) _03931_;
  assign _09505_ = nor_1589_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9175" *) nor_183_cse;
  assign _09506_ = _09505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9175" *) nor_213_cse;
  assign _09507_ = _09506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9176" *) cfg_out_precision_1_sva_6[0];
  assign _09508_ = _09507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9176" *) nand_207_cse;
  assign _09509_ = _07450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9178" *) or_1198_cse;
  assign _09510_ = _00070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9191" *) cfg_out_precision_1_sva_st_113[0];
  assign _09511_ = _03693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *) and_2360_cse;
  assign _09512_ = _09511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9204" *) cvt_unequal_tmp_20;
  assign _09513_ = chn_idata_data_sva_2_511_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9227" *) _00058_;
  assign _09514_ = _09513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9228" *) cvt_unequal_tmp_20;
  assign _09515_ = _09514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9228" *) cfg_mode_eql_1_sva_5;
  assign _09516_ = _04631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9229" *) cvt_unequal_tmp_21;
  assign _09517_ = _09516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9229" *) cfg_mode_eql_1_sva_6;
  assign _09518_ = _00058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9231" *) cvt_unequal_tmp_20;
  assign _09519_ = _09518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9231" *) cfg_mode_eql_1_sva_5;
  assign _09520_ = _07450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9234" *) _04947_;
  assign _09521_ = _09520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9234" *) or_1198_cse;
  assign _09522_ = _00070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9246" *) or_dcpl_160;
  assign or_4745_nl = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9257" *) cfg_out_precision_1_sva_st_113[0];
  assign or_4749_cse = _09520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9260" *) cfg_out_precision_1_sva_st_113[0];
  assign or_4755_nl = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9264" *) _05342_;
  assign _09523_ = mux_2232_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9266" *) and_2360_cse;
  assign or_3774_cse = or_dcpl_163 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9267" *) and_1021_cse;
  assign _09524_ = or_3774_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9267" *) cfg_out_precision_1_sva_st_113[0];
  assign _09525_ = nor_183_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9270" *) nor_213_cse;
  assign _09526_ = _09525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9271" *) cfg_out_precision_1_sva_6[0];
  assign _09527_ = _09526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9271" *) nand_207_cse;
  assign _09528_ = nor_151_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9290" *) or_1198_cse;
  assign _09529_ = nor_2219_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *) cfg_out_precision_1_sva_st_113[0];
  assign _09530_ = _03712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *) and_2360_cse;
  assign _09531_ = _09530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9294" *) cvt_unequal_tmp_20;
  assign _09532_ = cvt_unequal_tmp_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9310" *) mux_1888_nl;
  assign _09533_ = cvt_unequal_tmp_21 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9312" *) mux_1832_nl;
  assign _09534_ = _00069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9353" *) or_dcpl_160;
  assign _09535_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9364" *) nor_2219_cse;
  assign or_4788_cse = cfg_out_precision_1_sva_st_113[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9367" *) _05353_;
  assign _09536_ = or_3817_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9402" *) cfg_out_precision_1_sva_st_113[0];
  assign _09537_ = or_dcpl_178 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9481" *) _04631_;
  assign _09538_ = or_dcpl_195 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9484" *) _04631_;
  assign _09539_ = cfg_proc_precision_1_sva_st_108[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9489" *) _04634_;
  assign _09540_ = _04634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *) and_1059_cse;
  assign _09541_ = _09540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9494" *) _04631_;
  assign _09542_ = or_dcpl_197 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9495" *) _04631_;
  assign _09543_ = _08470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9497" *) _04582_;
  assign _09544_ = _09543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9497" *) cfg_mode_eql_1_sva_5;
  assign _09545_ = or_1431_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9501" *) _04631_;
  assign _09546_ = _09545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9501" *) _04566_;
  assign _09547_ = _09546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9501" *) cfg_mode_eql_1_sva_6;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_15_nl = _03750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9513" *) _03752_;
  assign _09548_ = _04582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9522" *) or_1198_cse;
  assign or_1587_cse = _09548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9522" *) cfg_mode_eql_1_sva_5;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_14_nl = _03755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9533" *) _03756_;
  assign _09549_ = nor_213_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9540" *) nor_1672_cse;
  assign _09550_ = _09549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9540" *) _04631_;
  assign _09551_ = _09550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *) _04566_;
  assign _09552_ = _09551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *) cfg_mode_eql_1_sva_6;
  assign _09553_ = _09552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *) _04150_;
  assign _09554_ = _09553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9541" *) _04173_;
  assign _09555_ = _07441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9543" *) _04582_;
  assign _09556_ = _09555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9543" *) cfg_mode_eql_1_sva_5;
  assign _09557_ = _09556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9544" *) or_1198_cse;
  assign _09558_ = _09557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9544" *) nor_50_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_13_nl = _03757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9554" *) _03758_;
  assign _09559_ = _08566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9562" *) _04632_;
  assign _09560_ = _08568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9564" *) _04632_;
  assign _09561_ = or_dcpl_353 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9568" *) _00058_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_12_nl = _03763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9582" *) _03765_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_11_nl = _03766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9595" *) _03767_;
  assign FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse = _03771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9605" *) and_1104_rgt;
  assign _09562_ = main_stage_v_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9606" *) _05373_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_10_nl = _03772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9614" *) _03773_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_9_nl = _03774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9627" *) _03775_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_8_nl = _03776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9640" *) _03777_;
  assign _09563_ = cfg_proc_precision_1_sva_st_65[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9647" *) nor_2219_cse;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_7_nl = _03779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9657" *) _03781_;
  assign FpIntToFloat_17U_5U_10U_is_inf_or_cse = _03782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9665" *) and_dcpl_617;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_6_nl = _03783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9672" *) _03784_;
  assign _09564_ = cfg_proc_precision_1_sva_st_101[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9679" *) _00069_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_5_nl = _03786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9689" *) _03788_;
  assign or_1919_cse = cfg_mode_eql_1_sva_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9696" *) cfg_out_precision_1_sva_6[0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_4_nl = _03790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9705" *) _03792_;
  assign _09565_ = _03793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9714" *) and_dcpl_631;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_3_nl = _03795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9722" *) _03797_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_2_nl = _03798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9735" *) _03799_;
  assign _09566_ = _03800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9749" *) and_dcpl_648;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_1_nl = _03801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9755" *) _03802_;
  assign FpIntToFloat_17U_5U_10U_o_expo_or_nl = _03804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9770" *) _03806_;
  assign or_3597_nl = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9811" *) mux_2011_nl;
  assign or_3600_nl = cfg_out_precision_1_sva_6[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9813" *) cfg_mode_eql_1_sva_6;
  assign or_3606_nl = cfg_mode_eql_1_sva_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9818" *) mux_2017_nl;
  assign or_3607_nl = _07616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9819" *) cfg_mode_eql_1_sva_6;
  assign or_3609_nl = nor_1629_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9820" *) cfg_mode_eql_1_sva_6;
  assign FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse = _03816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9832" *) and_1249_cse;
  assign _09567_ = _07438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9852" *) _04186_;
  assign _09568_ = _09567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9852" *) cfg_mode_eql_1_sva_4;
  assign _09569_ = or_1587_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9854" *) _00058_;
  assign _09570_ = cfg_proc_precision_1_sva_st_89[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9858" *) _04629_;
  assign _09571_ = or_2140_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9861" *) _05386_;
  assign _09572_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9864" *) _05387_;
  assign _09573_ = or_3623_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9869" *) _05388_;
  assign _09574_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9875" *) _04185_;
  assign _09575_ = or_2140_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9879" *) _05389_;
  assign _09576_ = reg_cfg_proc_precision_1_sva_st_40_cse[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9881" *) _04600_;
  assign _09577_ = or_3623_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9884" *) _05390_;
  assign _09578_ = _07568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9891" *) cfg_out_precision_1_sva_st_154[0];
  assign _09579_ = _09578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9891" *) nand_171_cse;
  assign or_3696_cse = or_dcpl_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9896" *) or_2251_nl;
  assign _09580_ = cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9966" *) cvt_16_IntSaturation_17U_16U_if_acc_4_nl[2];
  assign _09581_ = _09580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9966" *) and_dcpl_93;
  assign _09582_ = cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9972" *) cvt_15_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _09583_ = _09582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9972" *) and_dcpl_93;
  assign _09584_ = cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9978" *) cvt_14_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _09585_ = _09584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9978" *) and_dcpl_93;
  assign _09586_ = cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9984" *) cvt_13_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _09587_ = _09586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9984" *) and_dcpl_93;
  assign _09588_ = cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9990" *) cvt_12_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign _09589_ = _09588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9990" *) and_dcpl_93;
  assign _09590_ = cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9996" *) cvt_11_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign _09591_ = _09590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:9996" *) and_dcpl_93;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs <= 1'b0;
    else
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs <= _00987_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs <= _00974_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs <= _00960_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs <= _00947_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs <= _00934_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs <= _00921_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs <= _00908_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs <= _01115_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs <= _01101_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs <= _01087_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs <= _01073_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs <= _01058_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs <= _01043_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs <= _01028_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs <= _01014_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpMantRNE_24U_11U_else_and_svs <= 1'b0;
    else
      cvt_1_FpMantRNE_24U_11U_else_and_svs <= _00999_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs <= 1'b0;
    else
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs <= _00983_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    else
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= _00970_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    else
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= _00956_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    else
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= _00930_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    else
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= _00904_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    else
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= _00917_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    else
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= _01097_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    else
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= _01069_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    else
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= _01083_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva <= _00625_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs <= 1'b0;
    else
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs <= _01053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    else
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= _01039_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    else
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= _00943_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva <= _00617_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 <= _00311_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3 <= _00320_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 <= _00323_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3 <= _00325_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 <= _00305_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 <= _00307_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_15 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_15 <= _00295_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpMantRNE_17U_11U_else_and_4_svs <= 1'b0;
    else
      cvt_16_FpMantRNE_17U_11U_else_and_4_svs <= _00986_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_14 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_14 <= _00294_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_15_FpMantRNE_17U_11U_else_and_3_svs <= _00973_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_13 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_13 <= _00293_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_14_FpMantRNE_17U_11U_else_and_3_svs <= _00959_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_12 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_12 <= _00292_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_13_FpMantRNE_17U_11U_else_and_2_svs <= _00946_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_11 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_11 <= _00291_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_12_FpMantRNE_17U_11U_else_and_3_svs <= _00933_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_10 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_10 <= _00290_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_11_FpMantRNE_17U_11U_else_and_2_svs <= _00920_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_9 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_9 <= _00304_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_10_FpMantRNE_17U_11U_else_and_2_svs <= _00907_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_8 <= _00303_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_9_FpMantRNE_17U_11U_else_and_1_svs <= _01114_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_7 <= _00302_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    else
      cvt_8_FpMantRNE_17U_11U_else_and_3_svs <= _01100_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_6 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_6 <= _00301_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_7_FpMantRNE_17U_11U_else_and_2_svs <= _01086_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_5 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_5 <= _00300_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_6_FpMantRNE_17U_11U_else_and_2_svs <= _01072_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_4 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_4 <= _00299_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_5_FpMantRNE_17U_11U_else_and_1_svs <= _01057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_3 <= _00298_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    else
      cvt_4_FpMantRNE_17U_11U_else_and_2_svs <= _01042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_2 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_2 <= _00297_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_3_FpMantRNE_17U_11U_else_and_1_svs <= _01027_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_1 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_1 <= _00296_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    else
      cvt_2_FpMantRNE_17U_11U_else_and_1_svs <= _01013_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_unequal_tmp <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_unequal_tmp <= _00289_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpMantRNE_17U_11U_else_and_svs <= 1'b0;
    else
      cvt_1_FpMantRNE_17U_11U_else_and_svs <= _00998_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm <= _00566_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm <= _00559_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm <= _00565_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm <= _00574_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm <= _00563_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm <= _00564_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm <= _00562_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm <= _00560_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm <= _00561_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm <= _00570_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm <= _00573_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm <= _00571_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm <= _00572_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm <= _00569_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm <= _00567_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm <= _00568_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2 <= 1'b0;
    else
      IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2 <= _00681_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_nor_14_itm_2 <= 1'b0;
    else
      IsNaN_5U_10U_nor_14_itm_2 <= _00713_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 <= 1'b0;
    else
      IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 <= _00682_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_nor_1_itm_2 <= 1'b0;
    else
      IsNaN_5U_10U_nor_1_itm_2 <= _00714_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2 <= 1'b0;
    else
      IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2 <= _00683_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_nor_itm_2 <= 1'b0;
    else
      IsNaN_5U_10U_nor_itm_2 <= _00715_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_15_0_1 <= 16'b0000000000000000;
    else
      chn_idata_data_sva_2_15_0_1 <= _00771_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2 <= _00515_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2 <= _00514_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2 <= _00510_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2 <= _00509_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2 <= _00508_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2 <= _00525_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2 <= _00524_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2 <= _00523_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2 <= _00522_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2 <= _00521_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2 <= _00520_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2 <= _00519_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2 <= _00518_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2 <= _00516_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2 <= _00526_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5 <= _00533_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6 <= _00534_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6 <= _00535_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7 <= _00536_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6 <= _00537_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7 <= _00538_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7 <= _00539_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8 <= _00540_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6 <= _00541_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7 <= _00527_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7 <= _00528_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8 <= _00529_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7 <= _00530_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8 <= _00531_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8 <= _00532_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9 <= 15'b000000000000000;
    else
      IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9 <= _00542_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpMantRNE_24U_11U_else_and_svs_2 <= 1'b0;
    else
      cvt_1_FpMantRNE_24U_11U_else_and_svs_2 <= _01000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9 <= _00448_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    else
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2 <= _01015_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9 <= _00451_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    else
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2 <= _01029_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9 <= _00454_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    else
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2 <= _01044_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9 <= _00457_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    else
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2 <= _01059_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9 <= _00460_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    else
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2 <= _01074_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9 <= _00463_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    else
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 <= _01088_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9 <= _00466_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    else
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2 <= _01102_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9 <= _00469_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    else
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2 <= _01116_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9 <= _00472_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    else
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2 <= _00909_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9 <= _00430_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    else
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2 <= _00922_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9 <= _00433_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    else
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2 <= _00935_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9 <= _00436_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    else
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2 <= _00948_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9 <= _00439_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    else
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2 <= _00961_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9 <= _00442_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    else
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2 <= _00975_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9 <= _00445_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2 <= 1'b0;
    else
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2 <= _00988_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9 <= 5'b00000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9 <= _00475_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_sva_2 <= _00363_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 <= _00347_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_15_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_15_sva_2 <= _00353_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 <= _00337_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_14_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_14_sva_2 <= _00352_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 <= _00336_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_13_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_13_sva_2 <= _00351_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 <= _00335_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_12_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_12_sva_2 <= _00350_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 <= _00334_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_11_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_11_sva_2 <= _00349_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 <= _00333_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_10_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_10_sva_2 <= _00348_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 <= _00332_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_9_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_9_sva_2 <= _00362_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2 <= _00346_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_8_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_8_sva_2 <= _00361_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2 <= _00345_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_7_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_7_sva_2 <= _00360_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 <= _00344_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_6_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_6_sva_2 <= _00359_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 <= _00343_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_5_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_5_sva_2 <= _00358_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 <= _00342_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_4_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_4_sva_2 <= _00357_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 <= _00341_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_3_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_3_sva_2 <= _00356_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 <= _00340_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_2_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_2_sva_2 <= _00355_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 <= _00339_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_24U_11U_else_carry_1_sva_2 <= 1'b0;
    else
      FpMantRNE_24U_11U_else_carry_1_sva_2 <= _00354_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 <= 5'b00000;
    else
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 <= _00338_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_511_1 <= 1'b0;
    else
      chn_idata_data_sva_1_511_1 <= _00766_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_sva <= _00635_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_sva <= _00678_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva <= _00615_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_15_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_15_sva <= _00652_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva <= _00623_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_4_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_4_sva <= _00662_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva <= _00611_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_13_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_13_sva <= _00646_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva <= _00613_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_14_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_14_sva <= _00649_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm <= _00511_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva <= _00609_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_12_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_12_sva <= _00643_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva <= _00619_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_2_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_2_sva <= _00657_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva <= _00621_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva <= _00633_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva <= _00605_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_10_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_10_sva <= _00637_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva <= _00607_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_11_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_11_sva <= _00640_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva <= _00631_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_8_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_8_sva <= _00673_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva <= _00627_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_6_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_6_sva <= _00667_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva <= _00629_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_7_sva <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_7_sva <= _00670_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
    else
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= _00957_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
    else
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= _00944_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
    else
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= _00971_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2 <= 1'b0;
    else
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2 <= _00984_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
    else
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= _01098_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
    else
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= _00931_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
    else
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= _01054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
    else
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= _01040_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
    else
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= _01070_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
    else
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= _01084_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
    else
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= _00905_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
    else
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= _00918_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
    else
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= _01010_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
    else
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= _01024_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
    else
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= _01111_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 <= _00315_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 <= _00330_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 <= _00313_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3 <= _00327_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3 <= _00309_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_idata_data_sva_3_15_0_2_reg <= 10'b0000000000;
    else
      reg_chn_idata_data_sva_3_15_0_2_reg <= _01229_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_idata_data_sva_3_15_0_1_reg <= 5'b00000;
    else
      reg_chn_idata_data_sva_3_15_0_1_reg <= _01228_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_idata_data_sva_3_15_0_reg <= 1'b0;
    else
      reg_chn_idata_data_sva_3_15_0_reg <= _01230_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_out_precision_1_sva_st_136 <= 2'b00;
    else
      cfg_out_precision_1_sva_st_136 <= _00738_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_90 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_90 <= _00750_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_out_precision_1_sva_st_144 <= 2'b00;
    else
      cfg_out_precision_1_sva_st_144 <= _00739_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_102 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_102 <= _00744_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_108 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_108 <= _00745_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_out_precision_1_sva_st_156 <= 2'b00;
    else
      cfg_out_precision_1_sva_st_156 <= _00742_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm <= _01223_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm <= _01224_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm <= _01203_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm <= _01204_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8 <= _00316_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9 <= _00331_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg <= 10'b0000000000;
    else
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg <= _01226_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg <= 5'b00000;
    else
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg <= _01225_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm <= _01201_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm <= _01202_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4 <= _00513_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_4 <= _00583_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm <= _01199_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm <= _01200_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 <= _00312_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 <= _00314_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm <= _01197_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm <= _01198_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8 <= _00310_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm <= _01195_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm <= _01196_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7 <= _00308_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm <= _01193_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm <= _01194_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 <= _00306_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2 <= 1'b0;
    else
      cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2 <= _01120_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm <= _01221_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm <= _01222_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7 <= _00329_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm <= _01219_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm <= _01220_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8 <= _00328_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm <= _01217_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm <= _01218_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7 <= _00326_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm <= _01215_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm <= _01216_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 <= _00324_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2 <= 1'b0;
    else
      cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2 <= _01063_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm <= _01213_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm <= _01214_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm <= _01211_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm <= _01212_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 <= _00321_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2 <= 1'b0;
    else
      cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2 <= _01033_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm <= _01209_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm <= _01210_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7 <= _00319_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7 <= _00322_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm <= _01207_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm <= _01208_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6 <= _00318_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2 <= 1'b0;
    else
      cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2 <= _01004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm <= 4'b0000;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm <= _01205_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm <= 1'b0;
    else
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm <= _01206_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6 <= _00317_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_4 <= _00602_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_4 <= _00594_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_4 <= _00590_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_4 <= _00677_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_odata_data_13_0_lpi_1_dfm_1 <= 1'b0;
    else
      chn_odata_data_13_0_lpi_1_dfm_1 <= _00803_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_45 <= 1'b0;
    else
      cvt_else_equal_tmp_45 <= _01127_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_46 <= 1'b0;
    else
      cvt_else_equal_tmp_46 <= _01128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_nor_dfs_15 <= 1'b0;
    else
      cvt_else_nor_dfs_15 <= _01133_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_nor_dfs_10 <= 1'b0;
    else
      cvt_else_nor_dfs_10 <= _01131_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_33 <= 1'b0;
    else
      cvt_else_equal_tmp_33 <= _01125_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_34 <= 1'b0;
    else
      cvt_else_equal_tmp_34 <= _01126_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_nor_dfs_11 <= 1'b0;
    else
      cvt_else_nor_dfs_11 <= _01132_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_28 <= 1'b0;
    else
      cvt_else_equal_tmp_28 <= _01124_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cvt_else_nor_dfs_9_cse <= 1'b0;
    else
      reg_cvt_else_nor_dfs_9_cse <= _01232_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_4 <= _00666_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_16 <= 1'b0;
    else
      cvt_else_equal_tmp_16 <= _01123_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_4 <= _00661_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_9 <= 1'b0;
    else
      cvt_else_equal_tmp_9 <= _01130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_equal_tmp_5 <= 1'b0;
    else
      cvt_else_equal_tmp_5 <= _01129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_else_nor_dfs_2 <= 1'b0;
    else
      cvt_else_nor_dfs_2 <= _01134_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_3 <= _00598_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_3 <= _00577_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_3 <= _00581_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_3 <= _00585_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_sva_3 <= _00604_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1 <= 1'b0;
    else
      cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1 <= _00965_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_3 <= _00579_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_3 <= _00600_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_3 <= _00596_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_3 <= _00592_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_3 <= _00588_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_3 <= _00659_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_3 <= _00664_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_3 <= _00669_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_3 <= _00672_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_3 <= _00675_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_3 <= _00639_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_3 <= _00642_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_3 <= _00645_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_3 <= _00648_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_3 <= _00651_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_3 <= _00654_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_sva_3 <= _00680_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_4 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_4 <= _00656_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_out_precision_1_sva_6 <= 2'b00;
    else
      cfg_out_precision_1_sva_6 <= _00736_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_mode_eql_1_sva_6 <= 1'b0;
    else
      cfg_mode_eql_1_sva_6 <= _00735_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_unequal_tmp_21 <= 1'b0;
    else
      cvt_unequal_tmp_21 <= _01137_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _00992_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _00979_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _00966_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _00952_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _00939_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _00926_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _00913_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01121_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01106_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01092_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01078_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01064_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01019_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= 1'b0;
    else
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2 <= _01005_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_66 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_66 <= _00748_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= 1'b0;
    else
      cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= _00914_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= 1'b0;
    else
      cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= _00901_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_335_319_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_335_319_1 <= _00793_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 <= 1'b0;
    else
      cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 <= _00927_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_303_287_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_303_287_1 <= _00792_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 <= 1'b0;
    else
      cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 <= _01108_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_367_351_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_367_351_1 <= _00794_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= 1'b0;
    else
      cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= _00940_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_271_255_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_271_255_1 <= _00791_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 <= 1'b0;
    else
      cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 <= _01094_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_399_383_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_399_383_1 <= _00795_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg <= _01147_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg <= _01148_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_14_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_5U_10U_land_14_lpi_1_dfm_6 <= _00693_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 <= 1'b0;
    else
      cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 <= _00953_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_7_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_5U_10U_land_7_lpi_1_dfm_6 <= _00706_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_239_223_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_239_223_1 <= _00790_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2 <= 1'b0;
    else
      cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2 <= _01080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_431_415_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_431_415_1 <= _00796_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg <= _01149_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg <= _01150_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 <= 1'b0;
    else
      cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 <= _00967_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg <= _01159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg <= _01161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg <= _01143_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg <= _01141_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg <= _01160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg <= _01162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg <= _01164_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_207_191_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_207_191_1 <= _00789_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= 1'b0;
    else
      cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= _01066_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_463_447_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_463_447_1 <= _00797_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg <= _01151_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg <= _01145_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg <= _01152_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg <= _01146_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1 <= 1'b0;
    else
      cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1 <= _00980_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_sva_3 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_sva_3 <= _00266_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_175_159_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_175_159_1 <= _00788_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2 <= 1'b0;
    else
      cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2 <= _01050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_495_479_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_495_479_1 <= _00799_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg <= _01167_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg <= _01163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg <= _01168_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg <= _01144_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg <= _01142_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5 <= 15'b000000000000000;
    else
      FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5 <= _00267_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_143_127_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_143_127_1 <= _00787_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= 1'b0;
    else
      cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 <= _01036_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg <= _01155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg <= _01157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg <= _01165_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg <= _01156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg <= _01158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg <= _01166_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_4_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_4_lpi_1_dfm_5 <= _00700_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_8_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_8_lpi_1_dfm_5 <= _00708_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_11_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_11_lpi_1_dfm_5 <= _00687_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_13_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_13_lpi_1_dfm_5 <= _00691_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_lpi_1_dfm_5 <= _00712_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_12_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_12_lpi_1_dfm_5 <= _00689_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_10_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_10_lpi_1_dfm_5 <= _00685_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_9_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_9_lpi_1_dfm_5 <= _00710_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_6_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_6_lpi_1_dfm_5 <= _00704_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_5_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_5_lpi_1_dfm_5 <= _00702_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_3_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_3_lpi_1_dfm_5 <= _00698_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1 <= 10'b0000000000;
    else
      FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1 <= _00268_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3 <= _00517_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_111_95_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_111_95_1 <= _00786_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 <= 1'b0;
    else
      cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 <= _01021_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg <= _01153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg <= _01154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_2_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_2_lpi_1_dfm_4 <= _00696_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_79_63_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_79_63_1 <= _00800_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 <= 1'b0;
    else
      cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 <= _01007_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_1_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_5U_10U_land_1_lpi_1_dfm_3 <= _00695_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_15_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_5U_10U_land_15_lpi_1_dfm_3 <= _00694_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2 <= 1'b0;
    else
      cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2 <= _00994_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= 1'b0;
    else
      cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= _01008_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= 1'b0;
    else
      cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= _01037_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= 1'b0;
    else
      cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= _01081_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= 1'b0;
    else
      cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= _01095_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= 1'b0;
    else
      cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= _00915_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= 1'b0;
    else
      cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= _00941_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= 1'b0;
    else
      cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= _00954_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2 <= 1'b0;
    else
      cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2 <= _00981_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= 1'b0;
    else
      cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= _00968_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= 1'b0;
    else
      cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 <= _00928_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= 1'b0;
    else
      cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= _00902_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= 1'b0;
    else
      cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= _01109_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= 1'b0;
    else
      cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 <= _01067_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= 1'b0;
    else
      cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= _01051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= 1'b0;
    else
      cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 <= _01022_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_3_47_31_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_3_47_31_1 <= _00798_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2 <= 1'b0;
    else
      cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2 <= _00993_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2 <= _00256_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2 <= _00255_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2 <= _00254_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2 <= _00253_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2 <= _00252_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2 <= _00251_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2 <= _00265_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2 <= _00264_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2 <= _00263_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2 <= _00262_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2 <= _00261_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2 <= _00260_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2 <= _00259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2 <= _00258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2 <= 1'b0;
    else
      FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2 <= _00257_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_3 <= 1'b0;
    else
      main_stage_v_3 <= _01140_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2 <= 1'b0;
    else
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2 <= _01006_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_89 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_89 <= _00749_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2 <= 1'b0;
    else
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2 <= _01122_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_101 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_101 <= _00743_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_out_precision_1_sva_st_149 <= 2'b00;
    else
      cfg_out_precision_1_sva_st_149 <= _00740_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2 <= 1'b0;
    else
      cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2 <= _00985_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 <= _00284_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg <= _01191_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_sva_2 <= _00636_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_sva_2 <= _00679_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_sva_2 <= _00558_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= 1'b0;
    else
      cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= _00972_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 <= _00274_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg <= _01179_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2 <= _00616_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_2 <= _00653_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_15_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_15_sva_2 <= _00548_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= 1'b0;
    else
      cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= _00958_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 <= _00273_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg <= _01177_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg <= _01178_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2 <= _00614_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_2 <= _00650_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3 <= 1'b0;
    else
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3 <= _00512_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_14_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_14_sva_2 <= _00547_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= 1'b0;
    else
      cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= _00945_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 <= _00272_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2 <= _00612_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_2 <= _00647_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_13_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_13_sva_2 <= _00546_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= 1'b0;
    else
      cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= _00932_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 <= _00271_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg <= _01173_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg <= _01175_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2 <= _00610_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_2 <= _00644_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_12_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_12_sva_2 <= _00545_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= 1'b0;
    else
      cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= _00919_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 <= _00270_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2 <= _00608_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_2 <= _00641_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_11_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_11_sva_2 <= _00544_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= 1'b0;
    else
      cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= _00906_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 <= _00269_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2 <= _00606_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_2 <= _00638_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_10_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_10_sva_2 <= _00543_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= 1'b0;
    else
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= _01112_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= 1'b0;
    else
      cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= _01113_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6 <= 15'b000000000000000;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6 <= _00288_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 <= _00283_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2 <= _00634_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_9_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_9_sva_2 <= _00557_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 <= 1'b0;
    else
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 <= _01065_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2 <= 1'b0;
    else
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2 <= _01107_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= 1'b0;
    else
      cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2 <= _01099_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 <= _00282_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg <= _01189_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2 <= _00632_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_2 <= _00674_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_8_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_8_sva_2 <= _00556_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= 1'b0;
    else
      cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= _01085_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 <= _00281_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2 <= _00630_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_2 <= _00671_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_7_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_7_sva_2 <= _00555_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2 <= 1'b0;
    else
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2 <= _01079_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2 <= 1'b0;
    else
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2 <= _01093_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= 1'b0;
    else
      cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= _01071_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 <= _00280_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg <= _01185_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg <= _01187_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2 <= _00628_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_2 <= _00668_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_6_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_6_sva_2 <= _00554_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= 1'b0;
    else
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= _01055_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= 1'b0;
    else
      cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= _01056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 <= _00279_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg <= _01183_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2 <= _00626_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_5_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_5_sva_2 <= _00553_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2 <= 1'b0;
    else
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2 <= _01049_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= 1'b0;
    else
      cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2 <= _01041_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 <= _00278_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg <= _01181_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg <= _01169_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg <= 10'b0000000000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg <= _01171_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg <= _01182_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg <= _01184_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg <= _01186_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg <= _01188_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg <= _01190_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg <= _01170_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg <= _01172_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg <= _01174_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg <= _01176_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg <= _01180_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg <= 5'b00000;
    else
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg <= _01192_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2 <= _00624_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_2 <= _00663_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_4_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_4_sva_2 <= _00552_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= 1'b0;
    else
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= _01025_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= 1'b0;
    else
      cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= _01026_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6 <= 15'b000000000000000;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6 <= _00287_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 <= _00277_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2 <= _00622_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_3_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_3_sva_2 <= _00551_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 <= 1'b0;
    else
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 <= _01020_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 <= 1'b0;
    else
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 <= _01035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= 1'b0;
    else
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <= _01011_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= 1'b0;
    else
      cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2 <= _01012_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6 <= 15'b000000000000000;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6 <= _00286_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 <= _00276_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2 <= _00620_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_2 <= _00658_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_2_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_2_sva_2 <= _00550_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2 <= 1'b0;
    else
      cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2 <= _00996_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2 <= 1'b0;
    else
      cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2 <= _00997_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5 <= 15'b000000000000000;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5 <= _00285_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 <= 1'b0;
    else
      FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 <= _00275_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2 <= 15'b000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2 <= _00618_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_i_1_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntShiftRightSat_49U_6U_17U_i_1_sva_2 <= _00549_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2 <= 5'b00000;
    else
      cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2 <= _00982_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9 <= _00491_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_511_1 <= 1'b0;
    else
      chn_idata_data_sva_2_511_1 <= _00784_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8 <= _00481_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8 <= _00480_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8 <= _00479_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8 <= _00478_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8 <= _00477_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8 <= _00476_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b00000;
    else
      cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= _01110_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b00000;
    else
      cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= _00929_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b00000;
    else
      cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= _00955_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8 <= _00490_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8 <= _00489_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8 <= _00488_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b00000;
    else
      cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= _01068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b00000;
    else
      cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= _01082_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b00000;
    else
      cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= _01096_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b00000;
    else
      cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= _00903_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b00000;
    else
      cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= _00916_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b00000;
    else
      cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= _00942_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b00000;
    else
      cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= _00969_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8 <= _00487_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b00000;
    else
      cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= _01052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8 <= _00486_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8 <= _00485_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8 <= _00484_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b00000;
    else
      cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= _01009_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b00000;
    else
      cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= _01023_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b00000;
    else
      cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= _01038_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8 <= _00483_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2 <= 5'b00000;
    else
      cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2 <= _00995_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8 <= 10'b0000000000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8 <= _00482_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_1_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_1_sva_2 <= _00586_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_4_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_4_lpi_1_dfm_4 <= _00699_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_7_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_7_lpi_1_dfm_5 <= _00705_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_2 <= _00597_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_8_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_8_lpi_1_dfm_4 <= _00707_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_11_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_11_lpi_1_dfm_4 <= _00686_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_2 <= _00576_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_13_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_13_lpi_1_dfm_4 <= _00690_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_2 <= _00580_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_14_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_5U_10U_land_14_lpi_1_dfm_5 <= _00692_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_lpi_1_dfm_4 <= _00711_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_2 <= _00584_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_12_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_12_lpi_1_dfm_4 <= _00688_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_10_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_10_lpi_1_dfm_4 <= _00684_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_9_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_9_lpi_1_dfm_4 <= _00709_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_3 <= _00601_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_6_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_6_lpi_1_dfm_4 <= _00703_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_5_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_5_lpi_1_dfm_4 <= _00701_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_3 <= _00593_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_5U_10U_land_3_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_5U_10U_land_3_lpi_1_dfm_4 <= _00697_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_3 <= _00589_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_3 <= _00655_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_3 <= _00676_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_3 <= _00665_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_3 <= _00660_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_sva_2 <= _00603_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_3 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_3 <= _00582_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_2 <= _00578_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_10_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_10_sva_2 <= _00575_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_2 <= _00599_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_2 <= _00595_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_2 <= _00591_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_2 <= 1'b0;
    else
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_2 <= _00587_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_mode_eql_1_sva_5 <= 1'b0;
    else
      cfg_mode_eql_1_sva_5 <= _00734_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_unequal_tmp_20 <= 1'b0;
    else
      cvt_unequal_tmp_20 <= _01136_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_65 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_65 <= _00747_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_out_precision_1_sva_st_113 <= 2'b00;
    else
      cfg_out_precision_1_sva_st_113 <= _00737_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1 <= _00447_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1 <= _00446_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1 <= _00450_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1 <= _00449_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1 <= _00453_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1 <= _00452_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1 <= _00456_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1 <= _00455_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1 <= _00459_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1 <= _00458_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1 <= _00462_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1 <= _00461_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1 <= _00465_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1 <= _00464_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1 <= _00468_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1 <= _00467_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1 <= _00471_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1 <= _00470_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1 <= _00429_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1 <= _00428_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1 <= _00432_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1 <= _00431_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1 <= _00435_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1 <= _00434_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1 <= _00438_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1 <= _00437_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1 <= _00441_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1 <= _00440_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1 <= _00444_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1 <= _00443_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1 <= _00474_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1 <= 4'b0000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1 <= _00473_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_495_479_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_495_479_1 <= _00783_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_463_447_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_463_447_1 <= _00781_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_431_415_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_431_415_1 <= _00780_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_399_383_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_399_383_1 <= _00779_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_367_351_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_367_351_1 <= _00778_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_335_319_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_335_319_1 <= _00777_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_303_287_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_303_287_1 <= _00776_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_271_255_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_271_255_1 <= _00775_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_239_223_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_239_223_1 <= _00774_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_207_191_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_207_191_1 <= _00773_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_175_159_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_175_159_1 <= _00772_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_143_127_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_143_127_1 <= _00770_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_111_95_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_111_95_1 <= _00769_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_79_63_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_79_63_1 <= _00785_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_2_47_31_1 <= 17'b00000000000000000;
    else
      chn_idata_data_sva_2_47_31_1 <= _00782_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_2 <= 1'b0;
    else
      main_stage_v_2 <= _01139_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_1_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_1_sva_2 <= _00498_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_proc_precision_1_sva_st_40_cse <= 2'b00;
    else
      reg_cfg_proc_precision_1_sva_st_40_cse <= _01227_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_out_precision_1_sva_st_154 <= 2'b00;
    else
      cfg_out_precision_1_sva_st_154 <= _00741_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_5_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_5_sva_2 <= _00502_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_6_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_6_sva_1 <= _00503_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_7_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_7_sva_1 <= _00504_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_8_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_8_sva_1 <= _00505_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_10_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_10_sva_1 <= _00492_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_11_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_11_sva_1 <= _00493_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_12_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_12_sva_1 <= _00494_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_13_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_13_sva_1 <= _00495_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_14_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_14_sva_1 <= _00496_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_15_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_15_sva_1 <= _00497_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_sva_1 <= _00507_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_4_sva_1 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_4_sva_1 <= _00501_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_2_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_2_sva_2 <= _00499_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_3_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_3_sva_2 <= _00500_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntMulExt_33U_16U_49U_return_9_sva_2 <= 49'b0000000000000000000000000000000000000000000000000;
    else
      IntMulExt_33U_16U_49U_return_9_sva_2 <= _00506_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2 <= 1'b0;
    else
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2 <= _00989_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2 <= _00410_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= 1'b0;
    else
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= _00976_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2 <= _00390_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= 1'b0;
    else
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= _00962_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2 <= _00388_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= 1'b0;
    else
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= _00949_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2 <= _00386_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= 1'b0;
    else
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= _00936_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2 <= _00384_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= 1'b0;
    else
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= _00923_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2 <= _00382_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= 1'b0;
    else
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= _00910_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2 <= _00380_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= 1'b0;
    else
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= _01117_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2 <= _00408_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= 1'b0;
    else
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 <= _01103_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2 <= _00406_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= 1'b0;
    else
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= _01089_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2 <= _00404_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= 1'b0;
    else
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= _01075_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2 <= _00402_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= 1'b0;
    else
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= _01060_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2 <= _00400_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= 1'b0;
    else
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 <= _01045_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2 <= _00398_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= 1'b0;
    else
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= _01030_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2 <= _00396_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= 1'b0;
    else
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 <= _01016_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2 <= _00394_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2 <= 1'b0;
    else
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2 <= _01001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2 <= _00392_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_3 <= _00723_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_3 <= _00724_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_3 <= _00725_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_4_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_4_lpi_1_dfm_3 <= _00726_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_6_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_6_lpi_1_dfm_3 <= _00727_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_7_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_7_lpi_1_dfm_3 <= _00728_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_8_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_8_lpi_1_dfm_3 <= _00729_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_9_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_9_lpi_1_dfm_3 <= _00730_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_10_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_10_lpi_1_dfm_3 <= _00717_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_11_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_11_lpi_1_dfm_3 <= _00718_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_12_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_12_lpi_1_dfm_3 <= _00719_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_13_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_13_lpi_1_dfm_3 <= _00720_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_14_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_14_lpi_1_dfm_3 <= _00721_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_15_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_15_lpi_1_dfm_3 <= _00722_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_3 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_3 <= _00731_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2 <= _00427_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2 <= _00418_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2 <= _00419_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2 <= _00420_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2 <= _00421_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_nor_4_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_nor_4_itm_2 <= _00732_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2 <= _00716_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2 <= _00422_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2 <= _00423_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2 <= _00424_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2 <= _00425_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2 <= _00426_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2 <= _00412_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2 <= _00413_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2 <= _00414_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2 <= _00415_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2 <= _00416_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2 <= _00417_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2 <= 1'b0;
    else
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2 <= _01003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= _01018_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= _01032_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= _01047_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= _01062_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= _01077_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= _01091_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= _01105_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 <= _01119_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= _00912_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= _00925_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= _00938_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 <= _00951_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= _00964_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 <= _00978_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2 <= 1'b0;
    else
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2 <= _00991_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2 <= _00411_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2 <= 1'b0;
    else
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2 <= _00990_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2 <= _00371_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2 <= _00391_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= _00977_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2 <= _00370_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2 <= _00389_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= _00963_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2 <= _00369_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2 <= _00387_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= _00950_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2 <= _00368_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2 <= _00385_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= _00937_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2 <= _00367_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2 <= _00383_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= _00924_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2 <= _00366_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2 <= _00381_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= _00911_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2 <= _00365_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2 <= _00409_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= _01118_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2 <= _00364_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2 <= _00407_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= 1'b0;
    else
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2 <= _01104_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2 <= _00379_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2 <= _00405_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= _01090_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2 <= _00378_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2 <= _00403_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= _01076_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2 <= _00377_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2 <= _00401_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= _01061_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2 <= _00376_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2 <= _00399_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= 1'b0;
    else
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 <= _01046_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2 <= _00375_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2 <= _00397_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= _01031_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2 <= _00374_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2 <= _00395_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= 1'b0;
    else
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2 <= _01017_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_truncate_1_sva_2 <= 6'b000000;
    else
      cfg_truncate_1_sva_2 <= _00751_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_mode_eql_1_sva_4 <= 1'b0;
    else
      cfg_mode_eql_1_sva_4 <= _00733_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_unequal_tmp_19 <= 1'b0;
    else
      cvt_unequal_tmp_19 <= _01135_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_proc_precision_1_sva_st_64 <= 2'b00;
    else
      cfg_proc_precision_1_sva_st_64 <= _00746_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_507_479_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_507_479_1 <= _00765_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_475_447_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_475_447_1 <= _00764_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_443_415_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_443_415_1 <= _00763_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_411_383_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_411_383_1 <= _00762_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_379_351_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_379_351_1 <= _00761_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_347_319_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_347_319_1 <= _00760_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_315_287_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_315_287_1 <= _00759_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_283_255_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_283_255_1 <= _00758_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_251_223_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_251_223_1 <= _00756_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_219_191_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_219_191_1 <= _00755_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_187_159_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_187_159_1 <= _00754_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_155_127_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_155_127_1 <= _00753_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_123_95_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_123_95_1 <= _00752_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_91_63_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_91_63_1 <= _00768_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_59_31_1 <= 29'b00000000000000000000000000000;
    else
      chn_idata_data_sva_1_59_31_1 <= _00767_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2 <= _00373_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2 <= 1'b0;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2 <= _00393_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2 <= 1'b0;
    else
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2 <= _01002_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_idata_data_sva_1_27_0_1 <= 28'b0000000000000000000000000000;
    else
      chn_idata_data_sva_1_27_0_1 <= _00757_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2 <= 3'b000;
    else
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2 <= _00372_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_1 <= 1'b0;
    else
      main_stage_v_1 <= _01138_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_out_rsci_ld_core_psct_cse <= 1'b0;
    else
      reg_chn_out_rsci_ld_core_psct_cse <= _01231_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_255 <= 1'b0;
    else
      chn_out_rsci_d_255 <= _00857_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_240 <= 1'b0;
    else
      chn_out_rsci_d_240 <= _00853_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_127 <= 1'b0;
    else
      chn_out_rsci_d_127 <= _00813_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_96 <= 1'b0;
    else
      chn_out_rsci_d_96 <= _00898_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_95 <= 1'b0;
    else
      chn_out_rsci_d_95 <= _00897_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_64 <= 1'b0;
    else
      chn_out_rsci_d_64 <= _00888_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_63 <= 1'b0;
    else
      chn_out_rsci_d_63 <= _00887_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_32 <= 1'b0;
    else
      chn_out_rsci_d_32 <= _00878_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_31 <= 1'b0;
    else
      chn_out_rsci_d_31 <= _00877_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_0 <= 1'b0;
    else
      chn_out_rsci_d_0 <= _00804_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_239 <= 1'b0;
    else
      chn_out_rsci_d_239 <= _00852_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_224 <= 1'b0;
    else
      chn_out_rsci_d_224 <= _00848_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_223 <= 1'b0;
    else
      chn_out_rsci_d_223 <= _00847_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_208 <= 1'b0;
    else
      chn_out_rsci_d_208 <= _00843_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_207 <= 1'b0;
    else
      chn_out_rsci_d_207 <= _00842_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_192 <= 1'b0;
    else
      chn_out_rsci_d_192 <= _00838_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_191 <= 1'b0;
    else
      chn_out_rsci_d_191 <= _00837_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_176 <= 1'b0;
    else
      chn_out_rsci_d_176 <= _00833_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_175 <= 1'b0;
    else
      chn_out_rsci_d_175 <= _00832_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_160 <= 1'b0;
    else
      chn_out_rsci_d_160 <= _00827_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_159 <= 1'b0;
    else
      chn_out_rsci_d_159 <= _00825_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_144 <= 1'b0;
    else
      chn_out_rsci_d_144 <= _00820_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_143 <= 1'b0;
    else
      chn_out_rsci_d_143 <= _00819_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_128 <= 1'b0;
    else
      chn_out_rsci_d_128 <= _00814_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_112 <= 1'b0;
    else
      chn_out_rsci_d_112 <= _00809_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_111 <= 1'b0;
    else
      chn_out_rsci_d_111 <= _00808_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_80 <= 1'b0;
    else
      chn_out_rsci_d_80 <= _00893_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_79 <= 1'b0;
    else
      chn_out_rsci_d_79 <= _00892_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_48 <= 1'b0;
    else
      chn_out_rsci_d_48 <= _00883_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_47 <= 1'b0;
    else
      chn_out_rsci_d_47 <= _00882_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_16 <= 1'b0;
    else
      chn_out_rsci_d_16 <= _00829_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_15 <= 1'b0;
    else
      chn_out_rsci_d_15 <= _00826_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_237_234 <= 4'b0000;
    else
      chn_out_rsci_d_237_234 <= _00850_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_253_250 <= 4'b0000;
    else
      chn_out_rsci_d_253_250 <= _00855_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_221_218 <= 4'b0000;
    else
      chn_out_rsci_d_221_218 <= _00845_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_205_202 <= 4'b0000;
    else
      chn_out_rsci_d_205_202 <= _00840_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_189_186 <= 4'b0000;
    else
      chn_out_rsci_d_189_186 <= _00835_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_173_170 <= 4'b0000;
    else
      chn_out_rsci_d_173_170 <= _00830_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_157_154 <= 4'b0000;
    else
      chn_out_rsci_d_157_154 <= _00823_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_125_122 <= 4'b0000;
    else
      chn_out_rsci_d_125_122 <= _00811_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_109_106 <= 4'b0000;
    else
      chn_out_rsci_d_109_106 <= _00806_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_93_90 <= 4'b0000;
    else
      chn_out_rsci_d_93_90 <= _00895_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_61_58 <= 4'b0000;
    else
      chn_out_rsci_d_61_58 <= _00885_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_29_26 <= 4'b0000;
    else
      chn_out_rsci_d_29_26 <= _00875_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_105_97 <= 9'b000000000;
    else
      chn_out_rsci_d_105_97 <= _00805_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_73_65 <= 9'b000000000;
    else
      chn_out_rsci_d_73_65 <= _00889_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_41_33 <= 9'b000000000;
    else
      chn_out_rsci_d_41_33 <= _00879_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_9_1 <= 9'b000000000;
    else
      chn_out_rsci_d_9_1 <= _00899_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_271 <= 1'b0;
    else
      chn_out_rsci_d_271 <= _00874_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_270 <= 1'b0;
    else
      chn_out_rsci_d_270 <= _00873_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_269 <= 1'b0;
    else
      chn_out_rsci_d_269 <= _00872_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_268 <= 1'b0;
    else
      chn_out_rsci_d_268 <= _00871_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_267 <= 1'b0;
    else
      chn_out_rsci_d_267 <= _00870_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_266 <= 1'b0;
    else
      chn_out_rsci_d_266 <= _00869_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_265 <= 1'b0;
    else
      chn_out_rsci_d_265 <= _00868_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_264 <= 1'b0;
    else
      chn_out_rsci_d_264 <= _00867_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_263 <= 1'b0;
    else
      chn_out_rsci_d_263 <= _00866_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_262 <= 1'b0;
    else
      chn_out_rsci_d_262 <= _00865_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_261 <= 1'b0;
    else
      chn_out_rsci_d_261 <= _00864_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_260 <= 1'b0;
    else
      chn_out_rsci_d_260 <= _00863_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_259 <= 1'b0;
    else
      chn_out_rsci_d_259 <= _00861_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_258 <= 1'b0;
    else
      chn_out_rsci_d_258 <= _00860_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_257 <= 1'b0;
    else
      chn_out_rsci_d_257 <= _00859_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_256 <= 1'b0;
    else
      chn_out_rsci_d_256 <= _00858_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_249_241 <= 9'b000000000;
    else
      chn_out_rsci_d_249_241 <= _00854_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_233_225 <= 9'b000000000;
    else
      chn_out_rsci_d_233_225 <= _00849_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_217_209 <= 9'b000000000;
    else
      chn_out_rsci_d_217_209 <= _00844_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_201_193 <= 9'b000000000;
    else
      chn_out_rsci_d_201_193 <= _00839_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_185_177 <= 9'b000000000;
    else
      chn_out_rsci_d_185_177 <= _00834_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_169_161 <= 9'b000000000;
    else
      chn_out_rsci_d_169_161 <= _00828_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_153_145 <= 9'b000000000;
    else
      chn_out_rsci_d_153_145 <= _00822_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_137_129 <= 9'b000000000;
    else
      chn_out_rsci_d_137_129 <= _00815_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_121_113 <= 9'b000000000;
    else
      chn_out_rsci_d_121_113 <= _00810_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_89_81 <= 9'b000000000;
    else
      chn_out_rsci_d_89_81 <= _00894_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_57_49 <= 9'b000000000;
    else
      chn_out_rsci_d_57_49 <= _00884_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_25_17 <= 9'b000000000;
    else
      chn_out_rsci_d_25_17 <= _00862_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_254 <= 1'b0;
    else
      chn_out_rsci_d_254 <= _00856_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_238 <= 1'b0;
    else
      chn_out_rsci_d_238 <= _00851_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_222 <= 1'b0;
    else
      chn_out_rsci_d_222 <= _00846_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_206 <= 1'b0;
    else
      chn_out_rsci_d_206 <= _00841_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_190 <= 1'b0;
    else
      chn_out_rsci_d_190 <= _00836_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_174 <= 1'b0;
    else
      chn_out_rsci_d_174 <= _00831_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_158 <= 1'b0;
    else
      chn_out_rsci_d_158 <= _00824_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_142 <= 1'b0;
    else
      chn_out_rsci_d_142 <= _00818_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_126 <= 1'b0;
    else
      chn_out_rsci_d_126 <= _00812_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_110 <= 1'b0;
    else
      chn_out_rsci_d_110 <= _00807_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_94 <= 1'b0;
    else
      chn_out_rsci_d_94 <= _00896_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_78 <= 1'b0;
    else
      chn_out_rsci_d_78 <= _00891_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_62 <= 1'b0;
    else
      chn_out_rsci_d_62 <= _00886_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_46 <= 1'b0;
    else
      chn_out_rsci_d_46 <= _00881_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_30 <= 1'b0;
    else
      chn_out_rsci_d_30 <= _00876_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_14 <= 1'b0;
    else
      chn_out_rsci_d_14 <= _00821_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_141_138 <= 4'b0000;
    else
      chn_out_rsci_d_141_138 <= _00817_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_77_74 <= 4'b0000;
    else
      chn_out_rsci_d_77_74 <= _00890_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_45_42 <= 4'b0000;
    else
      chn_out_rsci_d_45_42 <= _00880_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_d_13_10 <= 4'b0000;
    else
      chn_out_rsci_d_13_10 <= _00816_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_in_rsci_ld_core_psct <= 1'b0;
    else
      chn_in_rsci_ld_core_psct <= _00802_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_out_rsci_iswt0 <= 1'b0;
    else
      chn_out_rsci_iswt0 <= _00900_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_in_rsci_iswt0 <= 1'b0;
    else
      chn_in_rsci_iswt0 <= _00801_;
  assign mux_153_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_275_nl;
  assign mux_150_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_270_nl;
  assign mux_143_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_263_nl;
  assign mux_131_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_236_nl;
  assign mux_121_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_tmp_218;
  assign mux_1415_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1414_nl : mux_tmp_1409;
  assign mux_1414_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1413_nl : mux_tmp_1409;
  assign mux_1413_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1409 : mux_1412_nl;
  assign mux_1412_nl = cfg_out_precision_1_sva_st_154[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00067_ : mux_tmp_1409;
  assign mux_1743_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2823_nl : or_2830_nl;
  assign mux_1734_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2809_nl : or_2815_nl;
  assign mux_1727_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2796_nl : or_2802_nl;
  assign mux_1720_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2784_nl : or_2789_nl;
  assign mux_1715_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2774_nl : or_2778_nl;
  assign mux_1711_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2764_nl : or_2768_nl;
  assign mux_1707_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2754_nl : or_2758_nl;
  assign mux_1704_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2744_nl : or_2749_nl;
  assign mux_1700_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2733_nl : or_2737_nl;
  assign mux_1697_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2723_nl : or_2727_nl;
  assign mux_1694_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2714_nl : or_2717_nl;
  assign mux_1692_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2705_nl : or_2709_nl;
  assign mux_1689_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2696_nl : or_2699_nl;
  assign mux_1687_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2688_nl : or_2691_nl;
  assign mux_803_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_801_nl : mux_802_nl;
  assign mux_802_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_208_nl : _00066_;
  assign mux_208_nl = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_389 : mux_207_nl;
  assign mux_207_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_50_cse : or_tmp_389;
  assign mux_801_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_92_nl : _00065_;
  assign mux_92_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_186_cse : and_dcpl_3;
  assign mux_799_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : mux_798_nl;
  assign mux_798_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1145_nl : _00064_;
  assign mux_789_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : or_1134_nl;
  assign mux_770_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : or_1118_nl;
  assign mux_454_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : or_733_nl;
  assign mux_449_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : or_724_nl;
  assign mux_1685_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1654_cse : mux_1684_nl;
  assign mux_1684_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_201_cse : mux_1683_nl;
  assign mux_1683_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1186_cse : mux_201_cse;
  assign mux_1674_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1654_cse : mux_1673_nl;
  assign mux_1673_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_786_cse_1 : mux_1672_nl;
  assign mux_1672_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1186_cse : mux_786_cse_1;
  assign mux_1663_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1661_nl : mux_1662_nl;
  assign mux_1662_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1310_cse : nor_1186_cse;
  assign mux_1661_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1309_cse : nor_1185_cse;
  assign mux_1660_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1654_cse : mux_1659_nl;
  assign mux_1659_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_660_cse : mux_1658_nl;
  assign mux_1658_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1186_cse : mux_660_cse;
  assign mux_1649_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1644_nl : mux_1648_nl;
  assign mux_1648_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1463_cse : mux_1647_nl;
  assign mux_1647_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1186_cse : mux_1463_cse;
  assign mux_1644_nl = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1460_cse : mux_1643_nl;
  assign mux_1643_nl = cfg_proc_precision_1_sva_st_64[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1185_cse : mux_1460_cse;
  assign mux_1640_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1633_nl : mux_1639_nl;
  assign mux_1639_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_767_cse : mux_1638_nl;
  assign mux_1638_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1186_cse : mux_767_cse;
  assign mux_1633_nl = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_719 : mux_1632_nl;
  assign mux_1632_nl = cfg_proc_precision_1_sva_st_64[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1185_cse : mux_tmp_719;
  assign mux_1627_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2239_cse : and_2160_nl;
  assign mux_1625_nl = _08964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1624_nl : mux_1623_nl;
  assign mux_1624_nl = cvt_1_FpMantRNE_24U_11U_else_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1622 : or_tmp_2612;
  assign mux_1623_nl = cvt_1_FpMantRNE_24U_11U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1622 : or_tmp_2612;
  assign mux_1621_nl = _08963_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1620_nl : mux_1619_nl;
  assign mux_1620_nl = cvt_2_FpMantRNE_24U_11U_else_and_1_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1618 : or_tmp_2610;
  assign mux_1619_nl = cvt_2_FpMantRNE_24U_11U_else_and_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1618 : or_tmp_2610;
  assign mux_1617_nl = _08961_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1616_nl : mux_1615_nl;
  assign mux_1616_nl = cvt_3_FpMantRNE_24U_11U_else_and_1_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1614 : or_tmp_2608;
  assign mux_1615_nl = cvt_3_FpMantRNE_24U_11U_else_and_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1614 : or_tmp_2608;
  assign mux_1613_nl = _08959_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1612_nl : mux_1611_nl;
  assign mux_1612_nl = cvt_4_FpMantRNE_24U_11U_else_and_2_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1610 : or_tmp_2606;
  assign mux_1611_nl = cvt_4_FpMantRNE_24U_11U_else_and_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1610 : or_tmp_2606;
  assign mux_1609_nl = _08957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1608_nl : mux_1607_nl;
  assign mux_1608_nl = cvt_5_FpMantRNE_24U_11U_else_and_1_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1606 : or_tmp_2604;
  assign mux_1607_nl = cvt_5_FpMantRNE_24U_11U_else_and_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1606 : or_tmp_2604;
  assign mux_1605_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1604_nl : nor_1198_nl;
  assign mux_1604_nl = _08954_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2161_nl : and_nl;
  assign mux_1603_nl = _08952_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1602_nl : mux_1601_nl;
  assign mux_1602_nl = cvt_7_FpMantRNE_24U_11U_else_and_2_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1600 : or_tmp_2595;
  assign mux_1601_nl = cvt_7_FpMantRNE_24U_11U_else_and_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1600 : or_tmp_2595;
  assign mux_1599_nl = _08950_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1598_nl : mux_1597_nl;
  assign mux_1598_nl = cvt_8_FpMantRNE_24U_11U_else_and_3_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1596 : or_tmp_2590;
  assign mux_1597_nl = cvt_8_FpMantRNE_24U_11U_else_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1596 : or_tmp_2590;
  assign mux_1595_nl = _08948_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1594_nl : mux_1593_nl;
  assign mux_1594_nl = cvt_9_FpMantRNE_24U_11U_else_and_1_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1592 : or_tmp_2588;
  assign mux_1593_nl = cvt_9_FpMantRNE_24U_11U_else_and_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1592 : or_tmp_2588;
  assign mux_1591_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1590_nl : nor_1200_nl;
  assign mux_1590_nl = _08944_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2162_nl : and_2243_nl;
  assign mux_1589_nl = _08942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1588_nl : mux_1587_nl;
  assign mux_1588_nl = cvt_11_FpMantRNE_24U_11U_else_and_2_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1586 : or_tmp_2579;
  assign mux_1587_nl = cvt_11_FpMantRNE_24U_11U_else_and_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1586 : or_tmp_2579;
  assign mux_1585_nl = _08940_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1584_nl : mux_1583_nl;
  assign mux_1584_nl = cvt_12_FpMantRNE_24U_11U_else_and_3_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1582 : or_tmp_2577;
  assign mux_1583_nl = cvt_12_FpMantRNE_24U_11U_else_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1582 : or_tmp_2577;
  assign mux_1581_nl = _08938_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1580_nl : mux_1579_nl;
  assign mux_1580_nl = cvt_13_FpMantRNE_24U_11U_else_and_2_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1578 : or_tmp_2575;
  assign mux_1579_nl = cvt_13_FpMantRNE_24U_11U_else_and_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1578 : or_tmp_2575;
  assign mux_1577_nl = _08936_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1576_nl : mux_1575_nl;
  assign mux_1576_nl = cvt_14_FpMantRNE_24U_11U_else_and_3_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1574 : or_tmp_2573;
  assign mux_1575_nl = cvt_14_FpMantRNE_24U_11U_else_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1574 : or_tmp_2573;
  assign mux_1573_nl = _08934_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1572_nl : mux_1571_nl;
  assign mux_1572_nl = cvt_15_FpMantRNE_24U_11U_else_and_3_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1570 : or_tmp_2571;
  assign mux_1571_nl = cvt_15_FpMantRNE_24U_11U_else_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1570 : or_tmp_2571;
  assign mux_1569_nl = _08932_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1568_nl : mux_1567_nl;
  assign mux_1568_nl = cvt_16_FpMantRNE_24U_11U_else_and_4_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1566 : or_tmp_2569;
  assign mux_1567_nl = cvt_16_FpMantRNE_24U_11U_else_and_4_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1566 : or_tmp_2569;
  assign mux_1565_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1201_nl : nor_1202_nl;
  assign mux_1564_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1203_nl : nor_1204_nl;
  assign mux_1563_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1205_nl : nor_1206_nl;
  assign mux_1562_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1207_nl : nor_1208_nl;
  assign mux_1561_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1209_nl : nor_1210_nl;
  assign mux_1560_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1211_nl : nor_1212_nl;
  assign mux_1559_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1213_nl : nor_1214_nl;
  assign mux_1558_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1215_nl : nor_1216_nl;
  assign mux_1557_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1217_nl : nor_1218_nl;
  assign mux_1556_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1219_nl : nor_1220_nl;
  assign mux_1555_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1221_nl : nor_1222_nl;
  assign mux_1554_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1223_nl : nor_1224_nl;
  assign mux_1553_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1225_nl : nor_1226_nl;
  assign mux_1552_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1227_nl : nor_1228_nl;
  assign mux_1551_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1229_nl : nor_1230_nl;
  assign mux_1550_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1231_nl : nor_1232_nl;
  assign mux_1549_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1233_nl : nor_1234_nl;
  assign mux_1548_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1235_nl : nor_1236_nl;
  assign mux_1547_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1237_nl : nor_1238_nl;
  assign mux_1546_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1239_nl : nor_1240_nl;
  assign mux_1545_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1241_nl : nor_1242_nl;
  assign mux_1544_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1243_nl : nor_1244_nl;
  assign mux_1543_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1245_nl : nor_1246_nl;
  assign mux_1542_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1247_nl : nor_1248_nl;
  assign mux_1541_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1249_nl : nor_1250_nl;
  assign mux_1540_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1251_nl : nor_1252_nl;
  assign mux_1539_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1253_nl : nor_1254_nl;
  assign mux_1538_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1255_nl : nor_1256_nl;
  assign mux_1537_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1257_nl : nor_1258_nl;
  assign mux_1536_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1259_nl : nor_1260_nl;
  assign mux_1535_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1261_nl : nor_1262_nl;
  assign mux_1534_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1263_nl : nor_1264_nl;
  assign mux_1533_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1532_nl : mux_tmp_189;
  assign mux_1532_nl = or_2433_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2432 : mux_1531_nl;
  assign mux_1531_nl = cfg_proc_precision_rsci_d[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00063_ : or_tmp_2432;
  assign mux_1472_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1467_nl : mux_1471_nl;
  assign mux_1471_nl = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1302_nl : main_stage_v_2;
  assign mux_1470_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1469 : nor_1303_nl;
  assign mux_1467_nl = or_2289_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2113_nl : main_stage_v_1;
  assign mux_1429_nl = or_2242_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_tmp_48 : mux_1428_nl;
  assign mux_1428_nl = chn_in_rsci_bawt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1427_nl : nand_tmp_48;
  assign mux_1427_nl = or_4524_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00062_ : nand_tmp_48;
  assign mux_1426_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1425_nl : or_5189_cse;
  assign mux_1425_nl = or_2251_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1424_nl : not_tmp_1709;
  assign mux_1424_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1423_nl : or_5189_cse;
  assign mux_1423_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1421_nl : or_5189_cse;
  assign mux_1421_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5189_cse : mux_1420_nl;
  assign mux_1420_nl = cfg_out_precision_1_sva_st_154[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00061_ : or_5189_cse;
  assign mux_2249_nl = cfg_out_precision_1_sva_st_113[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2248_nl : nor_2252_nl;
  assign mux_2248_nl = or_4857_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_out_precision_1_sva_st_113[1] : nor_2251_nl;
  assign mux_1266_nl = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1264 : mux_1265_nl;
  assign mux_1265_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1338_nl : mux_tmp_1264;
  assign mux_1262_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_223_nl : mux_1252_nl;
  assign mux_1252_nl = cfg_proc_precision_1_sva_st_108[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1227 : nor_1351_nl;
  assign mux_2281_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2396_nl : nor_2099_cse;
  assign mux_2280_nl = cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5086_cse : and_2780_nl;
  assign mux_2279_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2401_nl : nor_2099_cse;
  assign mux_2278_nl = cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5069_cse : and_2782_nl;
  assign mux_2277_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2406_nl : nor_2099_cse;
  assign mux_2276_nl = cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5053_cse : and_2784_nl;
  assign mux_1213_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_46_nl : mux_1212_nl;
  assign mux_1212_nl = cfg_proc_precision_1_sva_st_108[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_1992 : mux_1211_nl;
  assign mux_1211_nl = cfg_proc_precision_1_sva_st_108[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_199_nl : or_tmp_1992;
  assign mux_1204_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_45_nl : mux_1203_nl;
  assign mux_1203_nl = cfg_proc_precision_1_sva_st_108[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_1981 : mux_1202_nl;
  assign mux_1202_nl = cfg_proc_precision_1_sva_st_108[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_201_nl : or_tmp_1981;
  assign mux_2275_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2411_nl : nor_2099_cse;
  assign mux_2274_nl = cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5038_cse : and_2786_nl;
  assign mux_2273_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_3373_nl : nor_2099_cse;
  assign mux_2272_nl = cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1925_cse_1 : and_2788_nl;
  assign mux_1179_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1174_nl : mux_1178_nl;
  assign mux_1178_nl = or_1918_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_994 : mux_1177_nl;
  assign mux_1177_nl = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1176_nl : mux_989_cse;
  assign mux_1176_nl = or_1919_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_987 : mux_1175_nl;
  assign mux_1175_nl = cfg_out_precision_1_sva_6[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1403_nl : mux_tmp_987;
  assign mux_1174_nl = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_992 : mux_1173_nl;
  assign mux_1173_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1172_nl : mux_tmp_944;
  assign mux_1172_nl = cfg_out_precision_1_sva_st_149[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1142_cse : and_3372_nl;
  assign mux_2271_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2789_nl : nor_2099_cse;
  assign mux_2270_nl = cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1892_cse_1 : and_2791_nl;
  assign mux_1163_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1154_nl : mux_1053_cse;
  assign mux_1154_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1152 : mux_1153_nl;
  assign mux_1153_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00040_ : mux_tmp_1152;
  assign mux_2269_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2425_nl : nor_2099_cse;
  assign mux_2268_nl = cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1851_cse_1 : and_2793_nl;
  assign mux_1134_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1488_cse : mux_1133_nl;
  assign mux_1133_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_94 : nor_1489_cse;
  assign mux_2267_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2429_nl : nor_2099_cse;
  assign mux_2266_nl = cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1829_cse : and_2795_nl;
  assign mux_1127_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1433_nl : nor_1500_cse;
  assign FpIntToFloat_17U_5U_10U_else_mux_25_nl = cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_8 : or_1829_cse;
  assign FpMantRNE_17U_11U_else_mux_17_nl = or_3920_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_9_FpMantRNE_17U_11U_else_and_1_svs : cvt_9_FpMantRNE_17U_11U_else_and_1_tmp;
  assign mux_2265_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2433_nl : nor_2099_cse;
  assign mux_2264_nl = cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1789_cse_1 : and_2797_nl;
  assign mux_1116_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1107_nl : mux_1115_nl;
  assign mux_1115_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1113_nl : mux_1114_nl;
  assign mux_1114_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_tmp_175;
  assign mux_1113_nl = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1111 : mux_1112_nl;
  assign mux_1112_nl = cfg_proc_precision_1_sva_st_64[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00041_ : mux_tmp_1111;
  assign mux_1107_nl = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1105 : mux_1106_nl;
  assign mux_1106_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00041_ : mux_tmp_1105;
  assign mux_2263_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2437_nl : nor_2099_cse;
  assign mux_2262_nl = cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1752_cse_1 : and_2799_nl;
  assign mux_1091_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1090_nl : mux_1089_nl;
  assign mux_1090_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_961 : mux_tmp_1088;
  assign mux_1089_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1071_cse : mux_tmp_1088;
  assign mux_2261_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2441_nl : nor_2099_cse;
  assign mux_2260_nl = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1720_cse_1 : and_2801_nl;
  assign mux_1077_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1076_nl : mux_1075_nl;
  assign mux_1076_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_961 : mux_tmp_1074;
  assign mux_1075_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1071_cse : mux_tmp_1074;
  assign mux_1070_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1465_nl : mux_1069_nl;
  assign mux_1069_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2230_cse : nor_1466_nl;
  assign mux_2259_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2445_nl : nor_2099_cse;
  assign mux_2258_nl = cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1693_cse : and_2803_nl;
  assign mux_2257_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2449_nl : nor_2099_cse;
  assign mux_2256_nl = cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1659_cse_1 : and_2805_nl;
  assign mux_1054_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1045_nl : mux_1053_cse;
  assign mux_1045_nl = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1043 : mux_1044_nl;
  assign mux_1044_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00040_ : mux_tmp_1043;
  assign mux_1035_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1488_cse : mux_1034_nl;
  assign mux_1034_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_1078_cse : nor_1489_cse;
  assign mux_2255_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2453_nl : nor_2099_cse;
  assign mux_2254_nl = cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1625_cse : and_2807_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_13_nl = cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_4 : or_1693_cse;
  assign FpMantRNE_17U_11U_else_mux_9_nl = or_3879_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_FpMantRNE_17U_11U_else_and_1_svs : cvt_5_FpMantRNE_17U_11U_else_and_1_tmp;
  assign FpIntToFloat_17U_5U_10U_else_mux_7_nl = cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_2 : or_1625_cse;
  assign FpMantRNE_17U_11U_else_mux_5_nl = or_3860_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_3_FpMantRNE_17U_11U_else_and_1_svs : cvt_3_FpMantRNE_17U_11U_else_and_1_tmp;
  assign mux_2253_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2457_nl : nor_2099_cse;
  assign mux_2252_nl = cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1596_cse : and_2809_nl;
  assign mux_1018_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1017_nl : mux_1016_nl;
  assign mux_1017_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_945 : mux_tmp_1015;
  assign mux_1016_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1012_nl : mux_tmp_1015;
  assign mux_1012_nl = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_945 : nor_1508_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_4_nl = cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_1 : or_1596_cse;
  assign FpMantRNE_17U_11U_else_mux_3_nl = or_3850_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_2_FpMantRNE_17U_11U_else_and_1_svs : cvt_2_FpMantRNE_17U_11U_else_and_1_tmp;
  assign mux_1011_nl = or_425_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1510_nl : mux_1010_nl;
  assign mux_1010_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2237_cse : nor_1511_nl;
  assign mux_2251_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2461_nl : nor_2099_cse;
  assign mux_2250_nl = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1202_cse : and_2811_nl;
  assign mux_1004_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1519_nl : nor_1521_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_1_nl = cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp : or_1202_cse;
  assign FpMantRNE_17U_11U_else_mux_1_nl = or_3841_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_1_FpMantRNE_17U_11U_else_and_svs : cvt_1_FpMantRNE_17U_11U_else_and_tmp;
  assign mux_1000_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1526_nl : nor_1527_nl;
  assign mux_995_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_992 : mux_tmp_994;
  assign mux_982_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1537_nl : nor_1538_nl;
  assign mux_964_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_961 : mux_tmp_963;
  assign mux_959_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1547_nl : nor_1548_nl;
  assign mux_954_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_950_nl : mux_953_nl;
  assign mux_953_nl = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_951_nl : mux_952_nl;
  assign mux_952_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_321 : and_tmp_16;
  assign mux_951_nl = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_166 : nor_1555_nl;
  assign mux_950_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_321 : mux_949_nl;
  assign mux_949_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_117 : and_2186_cse;
  assign mux_943_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_940_nl : nor_1558_nl;
  assign mux_940_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1557_nl : nor_1556_cse;
  assign mux_939_nl = cfg_out_precision_1_sva_st_113[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1483_nl : or_1484_nl;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_32_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0 : IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_2_nl = _01589_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0 : IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_6_nl = and_tmp_50 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0 : IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_4_nl = or_dcpl_353 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_14_nl = or_dcpl_163 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_8_nl = or_3774_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_12_nl = or_3774_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_10_nl = or_3774_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_30_nl = mux_tmp_455 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0 : IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_16_nl = or_3817_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_20_nl = or_3817_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_18_nl = mux_1142_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0 : IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_28_nl = or_3817_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_22_nl = or_3817_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_26_nl = or_3817_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm : IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0;
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_24_nl = and_tmp_225 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0 : IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm;
  assign mux_937_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_261_nl : and_262_nl;
  assign mux_936_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_26_nl;
  assign mux_934_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1563_nl;
  assign mux_933_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_259_nl : and_260_nl;
  assign mux_932_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_25_nl;
  assign mux_930_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1566_nl;
  assign mux_929_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_257_nl : and_258_nl;
  assign mux_928_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_24_nl;
  assign mux_926_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1569_nl;
  assign mux_925_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_255_nl : and_256_nl;
  assign mux_924_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_23_nl;
  assign mux_922_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1572_nl;
  assign mux_921_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_917_nl : nor_1579_nl;
  assign mux_920_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_918_nl : nand_22_nl;
  assign mux_1832_nl = or_1157_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nor_1672_cse;
  assign mux_918_nl = or_1431_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nor_1672_cse;
  assign mux_917_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_916_nl : mux_915_nl;
  assign mux_916_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1577_nl : nor_1578_nl;
  assign mux_915_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1666_cse : mux_914_nl;
  assign mux_914_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1574_nl : nor_1575_nl;
  assign mux_913_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_252_nl : and_253_nl;
  assign mux_912_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_21_nl;
  assign mux_910_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1583_nl;
  assign mux_2239_nl = cfg_out_precision_1_sva_st_113[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4793_nl : and_2422_cse;
  assign mux_2237_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2422_cse : mux_2230_cse;
  assign mux_909_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2189_nl : nor_1588_nl;
  assign mux_908_nl = or_1159_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1409_nl : or_1402_nl;
  assign mux_906_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1585_nl : nor_1584_nl;
  assign mux_904_nl = FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_902_nl : mux_903_nl;
  assign mux_903_nl = or_1396_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1399_nl : or_tmp_1393;
  assign mux_902_nl = FpIntToFloat_17U_5U_10U_else_unequal_tmp_14 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1393_nl : or_tmp_1393;
  assign mux_899_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1375_nl : mux_898_nl;
  assign mux_898_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1379_nl : mux_897_nl;
  assign mux_897_nl = or_1157_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_1375 : or_1383_nl;
  assign mux_895_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_894_nl : or_1196_cse;
  assign mux_894_nl = and_2190_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_16_nl : mux_892_nl;
  assign mux_892_nl = FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_17_nl : or_1374_nl;
  assign mux_891_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_250_nl : and_251_nl;
  assign mux_890_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_15_nl;
  assign mux_888_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1596_nl;
  assign mux_887_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_883_nl : nor_1603_nl;
  assign mux_886_nl = or_1157_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_884_nl : mux_885_nl;
  assign mux_885_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1672_cse : or_4526_nl;
  assign mux_884_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nand_204_nl;
  assign mux_883_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_882_nl : mux_881_nl;
  assign mux_882_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1669_cse : nor_1602_nl;
  assign mux_881_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1666_cse : mux_880_nl;
  assign mux_880_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1598_nl : nor_1599_nl;
  assign mux_879_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_247_nl : and_248_nl;
  assign mux_878_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_13_nl;
  assign mux_876_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1608_nl;
  assign mux_875_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_871_nl : nor_1615_nl;
  assign mux_874_nl = or_1157_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_872_nl : mux_873_nl;
  assign mux_873_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1672_cse : or_4528_nl;
  assign mux_872_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nand_205_nl;
  assign mux_871_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_870_nl : mux_869_nl;
  assign mux_870_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1669_cse : nor_1614_nl;
  assign mux_869_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1666_cse : mux_868_nl;
  assign mux_868_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1610_nl : nor_1611_nl;
  assign mux_867_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_244_nl : and_245_nl;
  assign mux_866_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_11_nl;
  assign mux_864_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1620_nl;
  assign mux_863_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_242_nl : and_243_nl;
  assign mux_862_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_10_nl;
  assign mux_860_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1623_nl;
  assign mux_859_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_856_nl : mux_858_nl;
  assign mux_858_nl = or_1280_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_857_nl : nor_1630_cse;
  assign mux_857_nl = or_1159_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1630_cse : nor_1628_nl;
  assign mux_856_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1624_cse : mux_855_nl;
  assign mux_855_nl = or_300_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1626_cse : mux_854_nl;
  assign mux_854_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1624_cse : nor_1625_nl;
  assign mux_853_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_240_nl : and_241_nl;
  assign mux_852_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_9_nl;
  assign mux_850_nl = or_300_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1634_nl;
  assign mux_849_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_845_nl : nor_1641_nl;
  assign mux_848_nl = or_1157_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_846_nl : mux_847_nl;
  assign mux_847_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1672_cse : or_4530_nl;
  assign mux_846_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nand_206_nl;
  assign mux_845_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_844_nl : mux_843_nl;
  assign mux_844_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1669_cse : nor_1640_nl;
  assign mux_843_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1666_cse : mux_842_nl;
  assign mux_842_nl = or_300_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1636_nl : nor_1637_nl;
  assign mux_841_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_237_nl : and_238_nl;
  assign mux_840_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_7_nl;
  assign mux_838_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1646_nl;
  assign mux_837_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_235_nl : and_236_nl;
  assign mux_836_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_6_nl;
  assign mux_834_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1649_nl;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_nl = cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_3_FpMantRNE_17U_11U_else_acc_1_nl;
  assign mux_833_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_233_nl : and_234_nl;
  assign mux_832_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_5_nl;
  assign mux_830_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1652_nl;
  assign mux_2224_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2357_nl : or_4709_cse;
  assign mux_829_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1653_nl : nor_1655_nl;
  assign mux_828_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1209_nl : mux_827_cse;
  assign mux_826_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_825_nl : or_1196_cse;
  assign mux_825_nl = and_2191_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1198_cse : mux_823_nl;
  assign mux_823_nl = cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1201_nl : nand_4_nl;
  assign mux_822_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_229_nl : and_230_nl;
  assign mux_821_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_3_nl;
  assign mux_819_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1658_nl;
  assign mux_815_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_227_nl : and_228_nl;
  assign mux_814_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : nand_2_nl;
  assign mux_812_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1664_cse : nor_1665_nl;
  assign mux_811_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_807_nl : nor_1671_nl;
  assign mux_810_nl = or_1157_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_808_nl : mux_809_nl;
  assign mux_809_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1672_cse : or_4532_nl;
  assign mux_808_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nand_208_nl;
  assign mux_807_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_806_nl : mux_805_nl;
  assign mux_806_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1669_cse : nor_1670_nl;
  assign mux_805_nl = cvt_unequal_tmp_20 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1666_cse : nor_1667_nl;
  assign mux_794_nl = or_400_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_793_nl : mux_792_nl;
  assign mux_793_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_8 : and_136_nl;
  assign mux_792_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_8 : _00060_;
  assign mux_2223_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2222_nl : or_tmp_3849;
  assign mux_2222_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2219_nl : or_tmp_3849;
  assign mux_2219_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3849 : nor_2287_nl;
  assign mux_746_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_737_nl : mux_745_nl;
  assign mux_745_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_744_nl : main_stage_v_2;
  assign mux_744_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_743 : nor_1698_nl;
  assign mux_737_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_736_nl : main_stage_v_1;
  assign mux_736_nl = cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_720 : nor_1697_nl;
  assign mux_730_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_722_nl : mux_729_nl;
  assign mux_729_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_728_nl : main_stage_v_2;
  assign mux_728_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_727 : nor_1709_nl;
  assign mux_722_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_721_nl : main_stage_v_1;
  assign mux_721_nl = cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_720 : nor_1708_nl;
  assign mux_715_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_219_nl : and_221_nl;
  assign mux_714_nl = IsNaN_5U_10U_nor_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_417_cse : and_2196_nl;
  assign mux_2218_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2217_nl : or_tmp_3840;
  assign mux_2217_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2215_nl : or_tmp_3840;
  assign mux_2215_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3840 : nor_2290_nl;
  assign mux_698_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_690_nl : mux_697_nl;
  assign mux_697_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_696_nl : main_stage_v_2;
  assign mux_696_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_695 : nor_1737_nl;
  assign mux_690_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_689_nl : main_stage_v_1;
  assign mux_689_nl = cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_634 : nor_1772_cse;
  assign mux_684_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_677_nl : mux_683_nl;
  assign mux_683_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_682_nl : main_stage_v_2;
  assign mux_682_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_681 : nor_1746_nl;
  assign mux_677_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_676_nl : main_stage_v_1;
  assign mux_676_nl = cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_634 : nor_1745_nl;
  assign mux_671_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_216_nl : and_218_nl;
  assign mux_670_nl = IsNaN_5U_10U_nor_14_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_417_cse : and_2201_nl;
  assign mux_2214_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00046_ : mux_2213_nl;
  assign mux_2213_nl = and_2487_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2212_nl : _00046_;
  assign mux_2212_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2211_nl : _00046_;
  assign mux_2211_nl = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2208_nl : mux_2210_nl;
  assign mux_2210_nl = cfg_proc_precision_1_sva_st_64[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00046_ : mux_2208_nl;
  assign mux_644_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_636_nl : mux_643_nl;
  assign mux_643_nl = or_425_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_642_nl : main_stage_v_2;
  assign mux_642_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_641 : nor_1773_nl;
  assign mux_636_nl = or_961_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_635_nl : main_stage_v_1;
  assign mux_635_nl = cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_634 : nor_1772_cse;
  assign mux_630_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_213_nl : and_215_nl;
  assign mux_629_nl = IsNaN_5U_10U_nor_1_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_417_cse : and_2203_nl;
  assign mux_617_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_610_nl : mux_616_nl;
  assign mux_616_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_615_nl : main_stage_v_2;
  assign mux_615_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_614 : nor_1794_nl;
  assign mux_610_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_609_nl : main_stage_v_1;
  assign mux_609_nl = cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_597 : nor_1793_nl;
  assign mux_605_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_599_nl : mux_604_nl;
  assign mux_604_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_603_nl : main_stage_v_2;
  assign mux_603_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_602 : nor_1801_nl;
  assign mux_599_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_598_nl : main_stage_v_1;
  assign mux_598_nl = cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_597 : nor_1800_nl;
  assign mux_594_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_210_nl : and_212_nl;
  assign mux_593_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_592 : nor_1809_nl;
  assign mux_583_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_575_nl : mux_582_nl;
  assign mux_582_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_581_nl : main_stage_v_2;
  assign mux_581_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_580 : nor_1814_nl;
  assign mux_575_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_574_nl : main_stage_v_1;
  assign mux_574_nl = cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_435 : nor_1898_cse;
  assign mux_569_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_562_nl : mux_568_nl;
  assign mux_568_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_567_nl : main_stage_v_2;
  assign mux_567_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_566 : nor_1823_nl;
  assign mux_562_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_561_nl : main_stage_v_1;
  assign mux_561_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_560 : nor_1822_nl;
  assign mux_556_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_203_nl : and_205_nl;
  assign mux_555_nl = IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_417_cse : and_2213_nl;
  assign mux_544_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_533_nl : mux_543_nl;
  assign mux_543_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_541 : mux_542_nl;
  assign mux_542_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00037_ : mux_tmp_541;
  assign mux_533_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_532_nl : main_stage_v_1;
  assign mux_532_nl = cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_305 : nor_1980_cse;
  assign mux_528_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_521_nl : mux_527_nl;
  assign mux_527_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_526_nl : main_stage_v_2;
  assign mux_526_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_525 : nor_1848_nl;
  assign mux_521_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_520_nl : main_stage_v_1;
  assign mux_520_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_519 : nor_1847_nl;
  assign mux_516_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_199_nl : mux_515_nl;
  assign mux_515_nl = IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_174_cse : and_2217_nl;
  assign mux_505_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_495_nl : mux_504_nl;
  assign mux_504_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_502 : mux_503_nl;
  assign mux_503_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00037_ : mux_tmp_502;
  assign mux_495_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_494_nl : main_stage_v_1;
  assign mux_494_nl = cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_305 : nor_1980_cse;
  assign mux_490_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_483_nl : mux_489_nl;
  assign mux_489_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_488_nl : main_stage_v_2;
  assign mux_488_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_487 : nor_1869_nl;
  assign mux_483_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_482_nl : main_stage_v_1;
  assign mux_482_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_481 : nor_1868_nl;
  assign mux_478_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_195_nl : mux_477_nl;
  assign mux_477_nl = IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_174_cse : and_2221_nl;
  assign mux_472_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2005_cse : mux_471_nl;
  assign mux_471_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2004_cse : and_tmp_94;
  assign mux_467_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_462_nl : mux_466_nl;
  assign mux_466_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_465_nl : main_stage_v_2;
  assign mux_465_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_194_nl : mux_tmp_263;
  assign mux_462_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_461_nl : main_stage_v_1;
  assign mux_461_nl = cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_2011_cse;
  assign mux_458_nl = cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_456_nl : and_2856_nl;
  assign mux_456_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_93 : and_tmp_94;
  assign mux_453_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_18 : and_2230_cse;
  assign mux_450_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_129 : and_178_itm;
  assign mux_2186_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2185_nl : or_tmp_3763;
  assign mux_2185_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2183_nl : or_tmp_3763;
  assign mux_2183_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3763 : nor_2326_cse;
  assign mux_444_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_437_nl : mux_443_nl;
  assign mux_443_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_442_nl : main_stage_v_2;
  assign mux_442_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_185_nl : mux_tmp_441;
  assign mux_437_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_436_nl : main_stage_v_1;
  assign mux_436_nl = cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_435 : nor_1898_cse;
  assign mux_431_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_424_nl : mux_430_nl;
  assign mux_430_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_429_nl : main_stage_v_2;
  assign mux_429_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_428 : nor_1908_nl;
  assign mux_424_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_423_nl : main_stage_v_1;
  assign mux_423_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_422 : nor_1907_nl;
  assign mux_418_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_182_nl : and_183_nl;
  assign mux_408_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_399_nl : mux_407_nl;
  assign mux_407_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_405 : mux_406_nl;
  assign mux_406_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00037_ : mux_tmp_405;
  assign mux_399_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_398_nl : main_stage_v_1;
  assign mux_398_nl = cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_305 : nor_1980_cse;
  assign mux_394_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_388_nl : mux_393_nl;
  assign mux_393_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_392_nl : main_stage_v_2;
  assign mux_392_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_391 : nor_1932_nl;
  assign mux_388_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_387_nl : main_stage_v_1;
  assign mux_387_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_386 : nor_1931_nl;
  assign mux_383_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_179_nl : and_180_nl;
  assign mux_373_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_364_nl : mux_372_nl;
  assign mux_372_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_370 : mux_371_nl;
  assign mux_371_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00037_ : mux_tmp_370;
  assign mux_364_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_363_nl : main_stage_v_1;
  assign mux_363_nl = cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_305 : nor_1980_cse;
  assign mux_359_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_353_nl : mux_358_nl;
  assign mux_358_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_357_nl : main_stage_v_2;
  assign mux_357_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_356 : nor_1952_nl;
  assign mux_353_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_352_nl : main_stage_v_1;
  assign mux_352_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_351 : nor_1951_nl;
  assign mux_348_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_173_nl : mux_347_nl;
  assign mux_347_nl = cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_174_cse : and_2229_nl;
  assign mux_342_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1962_nl : mux_341_nl;
  assign mux_341_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00059_ : and_2230_cse;
  assign mux_2176_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2175_nl : or_4569_nl;
  assign mux_2175_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2265_nl : or_tmp_3768;
  assign mux_338_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_333_nl : mux_337_nl;
  assign mux_337_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_336_nl : main_stage_v_2;
  assign mux_336_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_172_nl : mux_tmp_263;
  assign mux_333_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_332_nl : main_stage_v_1;
  assign mux_332_nl = cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_2011_cse;
  assign mux_329_nl = IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_327_nl : mux_328_nl;
  assign mux_328_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_71 : and_171_nl;
  assign mux_327_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_71 : and_2230_cse;
  assign mux_322_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_16 : and_168_nl;
  assign mux_316_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_307_nl : mux_315_nl;
  assign mux_315_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_313 : mux_314_nl;
  assign mux_314_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00037_ : mux_tmp_313;
  assign mux_307_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_306_nl : main_stage_v_1;
  assign mux_306_nl = cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_305 : nor_1980_cse;
  assign mux_302_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_296_nl : mux_301_nl;
  assign mux_301_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_300_nl : main_stage_v_2;
  assign mux_300_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_299 : nor_1985_nl;
  assign mux_296_nl = or_513_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_295_nl : main_stage_v_1;
  assign mux_295_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_294 : nor_1984_nl;
  assign mux_291_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_164_nl : and_166_nl;
  assign mux_290_nl = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_67 : nor_1991_nl;
  assign mux_289_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1993_nl : mux_288_nl;
  assign mux_288_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1992_nl : and_1078_cse;
  assign mux_285_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_280_nl : mux_284_nl;
  assign mux_284_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_283_nl : main_stage_v_2;
  assign mux_283_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_161_nl : mux_tmp_263;
  assign mux_280_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_279_nl : main_stage_v_1;
  assign mux_279_nl = cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_2011_cse;
  assign mux_275_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_156_nl : and_160_nl;
  assign mux_271_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2005_cse : mux_270_nl;
  assign mux_270_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2004_cse : and_1078_cse;
  assign mux_267_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_261_nl : mux_266_nl;
  assign mux_266_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_265_nl : main_stage_v_2;
  assign mux_265_nl = cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_263 : mux_264_nl;
  assign mux_264_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2233_nl : mux_tmp_263;
  assign mux_261_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_260_nl : main_stage_v_1;
  assign mux_260_nl = cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_2011_cse;
  assign mux_257_nl = cfg_out_precision_1_sva_st_149[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_253 : mux_256_nl;
  assign mux_256_nl = and_2234_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_253 : mux_255_nl;
  assign mux_255_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_251 : mux_254_nl;
  assign mux_254_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_1078_cse : main_stage_v_2;
  assign mux_248_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_147_nl : and_tmp_52;
  assign mux_247_nl = or_1198_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2017_nl : mux_246_nl;
  assign mux_246_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2016_nl : and_2237_cse;
  assign mux_243_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_238_nl : mux_242_nl;
  assign mux_242_nl = or_423_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_241_nl : main_stage_v_2;
  assign mux_241_nl = cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_239 : and_2857_nl;
  assign mux_238_nl = or_419_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_237_nl : main_stage_v_1;
  assign mux_237_nl = cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_236 : nor_2020_nl;
  assign mux_235_nl = cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_232_nl : and_145_nl;
  assign mux_232_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_143_nl : and_2237_cse;
  assign mux_192_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_306_cse : or_tmp_378;
  assign mux_191_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_189 : mux_190_nl;
  assign mux_190_nl = cfg_mode_eql_1_sva_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_378 : _00058_;
  assign mux_167_nl = or_300_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_303_cse : mux_166_cse;
  assign mux_162_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2047_cse : nor_2048_nl;
  assign mux_159_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_in_rsci_bawt : and_132_nl;
  assign mux_155_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_110_cse : mux_154_nl;
  assign mux_154_nl = reg_cfg_proc_precision_1_sva_st_40_cse[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_8_cse : mux_110_cse;
  assign FpMantRNE_24U_11U_else_mux_1_nl = or_dcpl_350 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_1_FpMantRNE_24U_11U_else_and_svs : cvt_1_FpMantRNE_24U_11U_else_and_tmp;
  assign FpMantRNE_24U_11U_else_mux_3_nl = or_dcpl_348 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_2_FpMantRNE_24U_11U_else_and_1_svs : cvt_2_FpMantRNE_24U_11U_else_and_1_tmp;
  assign FpMantRNE_24U_11U_else_mux_5_nl = or_dcpl_346 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_3_FpMantRNE_24U_11U_else_and_1_svs : cvt_3_FpMantRNE_24U_11U_else_and_1_tmp;
  assign FpMantRNE_24U_11U_else_mux_7_nl = or_dcpl_344 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpMantRNE_24U_11U_else_and_2_svs : cvt_4_FpMantRNE_24U_11U_else_and_2_tmp;
  assign FpMantRNE_24U_11U_else_mux_9_nl = or_dcpl_342 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_FpMantRNE_24U_11U_else_and_1_svs : cvt_5_FpMantRNE_24U_11U_else_and_1_tmp;
  assign FpMantRNE_24U_11U_else_mux_11_nl = or_dcpl_340 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpMantRNE_24U_11U_else_and_2_svs : cvt_6_FpMantRNE_24U_11U_else_and_2_tmp;
  assign FpMantRNE_24U_11U_else_mux_13_nl = or_dcpl_338 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpMantRNE_24U_11U_else_and_2_svs : cvt_7_FpMantRNE_24U_11U_else_and_2_tmp;
  assign FpMantRNE_24U_11U_else_mux_15_nl = or_dcpl_336 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpMantRNE_24U_11U_else_and_3_svs : cvt_8_FpMantRNE_24U_11U_else_and_3_tmp;
  assign FpMantRNE_24U_11U_else_mux_17_nl = or_dcpl_334 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_9_FpMantRNE_24U_11U_else_and_1_svs : cvt_9_FpMantRNE_24U_11U_else_and_1_tmp;
  assign FpMantRNE_24U_11U_else_mux_19_nl = or_dcpl_332 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpMantRNE_24U_11U_else_and_2_svs : cvt_10_FpMantRNE_24U_11U_else_and_2_tmp;
  assign FpMantRNE_24U_11U_else_mux_21_nl = or_dcpl_330 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpMantRNE_24U_11U_else_and_2_svs : cvt_11_FpMantRNE_24U_11U_else_and_2_tmp;
  assign FpMantRNE_24U_11U_else_mux_23_nl = or_dcpl_328 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpMantRNE_24U_11U_else_and_3_svs : cvt_12_FpMantRNE_24U_11U_else_and_3_tmp;
  assign FpMantRNE_24U_11U_else_mux_25_nl = or_dcpl_326 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpMantRNE_24U_11U_else_and_2_svs : cvt_13_FpMantRNE_24U_11U_else_and_2_tmp;
  assign FpMantRNE_24U_11U_else_mux_27_nl = or_dcpl_324 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpMantRNE_24U_11U_else_and_3_svs : cvt_14_FpMantRNE_24U_11U_else_and_3_tmp;
  assign FpMantRNE_24U_11U_else_mux_29_nl = or_dcpl_322 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpMantRNE_24U_11U_else_and_3_svs : cvt_15_FpMantRNE_24U_11U_else_and_3_tmp;
  assign FpMantRNE_24U_11U_else_mux_31_nl = or_dcpl_320 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpMantRNE_24U_11U_else_and_4_svs : cvt_16_FpMantRNE_24U_11U_else_and_4_tmp;
  assign mux_91_nl = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_90_nl : or_181_nl;
  assign mux_90_nl = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_89_nl = _07623_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_179_nl : mux_88_nl;
  assign mux_88_nl = _08290_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_87_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2057_nl : nor_2058_nl;
  assign mux_86_nl = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_85_nl : or_173_nl;
  assign mux_85_nl = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_84_nl = _07624_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_171_nl : mux_83_nl;
  assign mux_83_nl = _08276_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_82_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2059_nl : nor_2060_nl;
  assign mux_81_nl = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_80_nl : or_165_nl;
  assign mux_80_nl = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_79_nl = _07625_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_163_nl : mux_78_nl;
  assign mux_78_nl = _08262_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_77_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2061_nl : nor_2062_nl;
  assign mux_76_nl = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_75_nl : or_157_nl;
  assign mux_75_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : nand_231_nl;
  assign mux_74_nl = _07626_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_152_nl : mux_73_nl;
  assign mux_73_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_150_nl;
  assign mux_72_nl = _08247_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_147_nl : mux_71_nl;
  assign mux_71_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_145_nl;
  assign mux_70_nl = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_69_nl : or_142_nl;
  assign mux_69_nl = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_68_nl = _07627_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_140_nl : mux_67_nl;
  assign mux_67_nl = _08232_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_66_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2063_nl : nor_2064_nl;
  assign mux_65_nl = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_64_nl : or_134_nl;
  assign mux_64_nl = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_63_nl = _07628_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_132_nl : mux_62_nl;
  assign mux_62_nl = _08218_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_61_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2065_nl : nor_2066_nl;
  assign mux_60_nl = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_59_nl : or_126_nl;
  assign mux_59_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : nand_232_nl;
  assign mux_58_nl = _07629_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_121_nl : mux_57_nl;
  assign mux_57_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_119_nl;
  assign mux_56_nl = _08203_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_116_nl : mux_55_nl;
  assign mux_55_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_114_nl;
  assign mux_54_nl = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_53_nl : or_111_nl;
  assign mux_53_nl = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_52_nl = _07630_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_109_nl : mux_51_nl;
  assign mux_51_nl = _08188_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_50_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2067_nl : nor_2068_nl;
  assign mux_49_nl = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_48_nl : or_103_nl;
  assign mux_48_nl = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_47_nl = _07631_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_101_nl : mux_46_nl;
  assign mux_46_nl = _08174_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_45_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2069_nl : nor_2070_nl;
  assign mux_44_nl = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_43_nl : or_95_nl;
  assign mux_43_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : nand_233_nl;
  assign mux_42_nl = _07632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_90_nl : mux_tmp_39;
  assign mux_41_nl = _08162_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_88_nl : mux_40_nl;
  assign mux_40_nl = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_39;
  assign mux_38_nl = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_37_nl : or_83_nl;
  assign mux_37_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : nand_234_nl;
  assign mux_36_nl = _07633_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_78_nl : mux_35_nl;
  assign mux_35_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_76_nl;
  assign mux_34_nl = _08148_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_73_nl : mux_33_nl;
  assign mux_33_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_71_nl;
  assign mux_32_nl = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_31_nl : or_68_nl;
  assign mux_31_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : nand_235_nl;
  assign mux_30_nl = _07634_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_63_nl : mux_29_nl;
  assign mux_29_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_61_nl;
  assign mux_28_nl = _08132_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_58_nl : mux_27_nl;
  assign mux_27_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_56_nl;
  assign mux_26_nl = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_25_nl : or_53_nl;
  assign mux_25_nl = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_24_nl = _07635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_51_nl : mux_23_nl;
  assign mux_23_nl = _08117_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_22_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2071_nl : nor_2072_nl;
  assign mux_21_nl = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_20_nl : or_45_nl;
  assign mux_20_nl = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_19_nl = _07636_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_43_nl : mux_18_nl;
  assign mux_18_nl = _08103_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_17_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2073_nl : nor_2074_nl;
  assign mux_16_nl = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_15_nl : or_37_nl;
  assign mux_15_nl = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_14_nl = _07637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_35_nl : mux_13_nl;
  assign mux_13_nl = _08089_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_11_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2075_nl : nor_2076_nl;
  assign mux_10_nl = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_9_nl : or_28_nl;
  assign mux_9_nl = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_8_nl = or_17_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_19_nl : mux_7_nl;
  assign mux_7_nl = or_14_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_24 : mux_tmp_6;
  assign mux_5_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_98_nl : mux_4_nl;
  assign mux_4_nl = _08075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2242_nl : mux_3_nl;
  assign mux_3_nl = or_14_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2239_cse : and_2240_nl;
  assign mux_2_nl = _05732_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1_nl : or_9_nl;
  assign mux_1_nl = or_17_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_13_nl : or_11_nl;
  assign mux_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2081_nl : nor_2082_nl;
  assign cvt_mux_2341_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_292_nl : cvt_if_mux_232_nl;
  assign cvt_if_mux_232_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[4] : IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3;
  assign cvt_mux_2340_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_295_nl : cvt_if_mux_235_nl;
  assign cvt_if_mux_235_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_15_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_109_nl = cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_47_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_47_nl = IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_sva_3;
  assign cvt_mux_2356_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_274_nl : cvt_if_mux_218_nl;
  assign cvt_if_mux_218_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_495_479_1[0];
  assign cvt_mux_2336_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_463_447_1[1] : cvt_else_mux1h_276_nl;
  assign cvt_mux_2337_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_463_447_1[1] : cvt_if_mux_220_nl;
  assign cvt_if_mux_220_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_14_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_102_nl = cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 : FpFloatToInt_16U_5U_10U_else_mux_44_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_44_nl = chn_idata_data_sva_3_495_479_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 : FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  assign cvt_mux_2368_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_255_nl : cvt_if_mux_203_nl;
  assign cvt_if_mux_203_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_463_447_1[0];
  assign cvt_mux_2332_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_431_415_1[1] : chn_odata_data_mux_1_nl;
  assign chn_odata_data_mux_1_nl = or_dcpl_195 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_odata_data_13_0_lpi_1_dfm_1 : chn_odata_data_13_0_lpi_1_dfm_1_mx0w0;
  assign cvt_mux_2333_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_431_415_1[1] : cvt_if_mux_205_nl;
  assign cvt_if_mux_205_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_13_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_95_nl = cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_41_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_41_nl = chn_idata_data_sva_3_463_447_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  assign cvt_mux_2372_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_236_nl : cvt_if_mux_188_nl;
  assign cvt_if_mux_188_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_431_415_1[0];
  assign cvt_mux_2328_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_399_383_1[1] : cvt_else_mux1h_238_nl;
  assign cvt_mux_2329_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_399_383_1[1] : cvt_if_mux_190_nl;
  assign cvt_if_mux_190_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_12_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_88_nl = cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_38_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_38_nl = chn_idata_data_sva_3_431_415_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  assign cvt_mux_2370_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_217_nl : cvt_if_mux_173_nl;
  assign cvt_if_mux_173_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_399_383_1[0];
  assign cvt_mux_2324_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_367_351_1[1] : cvt_else_mux1h_219_nl;
  assign cvt_mux_2325_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_367_351_1[1] : cvt_if_mux_175_nl;
  assign cvt_if_mux_175_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_11_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_81_nl = cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_35_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_35_nl = chn_idata_data_sva_3_399_383_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  assign cvt_mux_2366_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_198_nl : cvt_if_mux_158_nl;
  assign cvt_if_mux_158_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_367_351_1[0];
  assign cvt_mux_2320_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_335_319_1[1] : cvt_else_mux1h_200_nl;
  assign cvt_mux_2321_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_335_319_1[1] : cvt_if_mux_160_nl;
  assign cvt_if_mux_160_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_10_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_74_nl = cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_32_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_32_nl = chn_idata_data_sva_3_367_351_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  assign cvt_mux_2364_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_179_nl : cvt_if_mux_143_nl;
  assign cvt_if_mux_143_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_335_319_1[0];
  assign cvt_mux_2316_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_303_287_1[1] : cvt_else_mux1h_181_nl;
  assign cvt_mux_2317_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_303_287_1[1] : cvt_if_mux_145_nl;
  assign cvt_if_mux_145_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_9_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_67_nl = cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_29_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_29_nl = chn_idata_data_sva_3_335_319_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  assign cvt_mux_2362_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_160_nl : cvt_if_mux_128_nl;
  assign cvt_if_mux_128_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_303_287_1[0];
  assign cvt_mux_2312_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_271_255_1[1] : cvt_else_mux1h_162_nl;
  assign cvt_mux_2313_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_271_255_1[1] : cvt_if_mux_130_nl;
  assign cvt_if_mux_130_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_8_nl : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1[0];
  assign FpFloatToInt_16U_5U_10U_mux_60_nl = cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_26_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_26_nl = chn_idata_data_sva_3_303_287_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  assign cvt_mux_2360_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_141_nl : cvt_if_mux_113_nl;
  assign cvt_if_mux_113_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_271_255_1[0];
  assign cvt_mux_2308_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_239_223_1[1] : cvt_else_mux1h_143_nl;
  assign cvt_mux_2309_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_239_223_1[1] : cvt_if_mux_115_nl;
  assign cvt_if_mux_115_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_7_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_53_nl = cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 : FpFloatToInt_16U_5U_10U_else_mux_23_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_23_nl = chn_idata_data_sva_3_271_255_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2 : FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  assign cvt_mux_2358_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_122_nl : cvt_if_mux_98_nl;
  assign cvt_if_mux_98_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_239_223_1[0];
  assign cvt_mux_2304_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_207_191_1[1] : cvt_else_mux1h_124_nl;
  assign cvt_mux_2305_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_207_191_1[1] : cvt_if_mux_100_nl;
  assign cvt_if_mux_100_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_6_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_46_nl = cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2 : FpFloatToInt_16U_5U_10U_else_mux_20_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_20_nl = chn_idata_data_sva_3_239_223_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2 : FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  assign cvt_mux_2354_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_103_nl : cvt_if_mux_83_nl;
  assign cvt_if_mux_83_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_207_191_1[0];
  assign cvt_mux_2300_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_175_159_1[1] : cvt_else_mux1h_105_nl;
  assign cvt_mux_2301_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_175_159_1[1] : cvt_if_mux_85_nl;
  assign cvt_if_mux_85_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_5_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_39_nl = cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_17_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_17_nl = chn_idata_data_sva_3_207_191_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  assign cvt_mux_2352_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_84_nl : cvt_if_mux_68_nl;
  assign cvt_if_mux_68_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_175_159_1[0];
  assign cvt_mux_2296_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_143_127_1[1] : cvt_else_mux1h_86_nl;
  assign cvt_mux_2297_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_143_127_1[1] : cvt_if_mux_70_nl;
  assign cvt_if_mux_70_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_4_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_32_nl = cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2 : FpFloatToInt_16U_5U_10U_else_mux_14_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_14_nl = chn_idata_data_sva_3_175_159_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2 : FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  assign cvt_mux_2350_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_65_nl : cvt_if_mux_53_nl;
  assign cvt_if_mux_53_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[14] : chn_idata_data_sva_3_143_127_1[0];
  assign cvt_mux_2292_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_111_95_1[1] : cvt_else_mux1h_67_nl;
  assign cvt_mux_2293_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_111_95_1[1] : cvt_if_mux_55_nl;
  assign cvt_if_mux_55_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_3_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_25_nl = cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_11_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_11_nl = chn_idata_data_sva_3_143_127_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  assign cvt_mux_2348_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_46_nl : cvt_if_mux_38_nl;
  assign cvt_if_mux_38_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_111_95_1[0];
  assign cvt_mux_2288_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_79_63_1[1] : cvt_else_mux1h_48_nl;
  assign cvt_mux_2289_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_79_63_1[1] : cvt_if_mux_40_nl;
  assign cvt_if_mux_40_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_2_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_18_nl = cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_8_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_8_nl = chn_idata_data_sva_3_111_95_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  assign cvt_mux_2346_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_27_nl : cvt_if_mux_23_nl;
  assign cvt_if_mux_23_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[4] : chn_idata_data_sva_3_79_63_1[0];
  assign cvt_mux_2284_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_47_31_1[1] : cvt_else_mux1h_29_nl;
  assign cvt_mux_2285_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_47_31_1[1] : cvt_if_mux_25_nl;
  assign cvt_if_mux_25_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_1_nl : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_11_nl = cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 : FpFloatToInt_16U_5U_10U_else_mux_5_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_5_nl = chn_idata_data_sva_3_79_63_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1 : FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  assign cvt_mux_2373_nl = cvt_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_mux1h_8_nl : cvt_if_mux_8_nl;
  assign cvt_if_mux_8_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_chn_idata_data_sva_3_15_0_1_reg[4] : chn_idata_data_sva_3_47_31_1[0];
  assign cvt_mux_2280_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_chn_idata_data_sva_3_15_0_2_reg[0] : cvt_else_mux1h_10_nl;
  assign cvt_mux_2281_nl = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_chn_idata_data_sva_3_15_0_2_reg[0] : cvt_if_mux_10_nl;
  assign cvt_if_mux_10_nl = cvt_else_equal_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_nl : reg_chn_idata_data_sva_3_15_0_2_reg[0];
  assign FpFloatToInt_16U_5U_10U_mux_4_nl = cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2 : FpFloatToInt_16U_5U_10U_else_mux_2_nl;
  assign FpFloatToInt_16U_5U_10U_else_mux_2_nl = chn_idata_data_sva_3_47_31_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2 : FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  assign mux_2362_nl = or_5254_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00057_ : or_tmp_4097;
  assign mux_2361_nl = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2353 : mux_2360_nl;
  assign mux_2360_nl = cfg_proc_precision_1_sva_st_102[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00056_ : mux_tmp_2353;
  assign mux_2349_nl = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2341 : mux_2348_nl;
  assign mux_2348_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00054_ : mux_tmp_2341;
  assign mux_2344_nl = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2336 : mux_2343_nl;
  assign mux_2343_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00051_ : mux_tmp_2336;
  assign mux_2338_nl = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2330 : mux_2337_nl;
  assign mux_2337_nl = cfg_proc_precision_1_sva_st_102[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00053_ : mux_tmp_2330;
  assign mux_2332_nl = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2324 : mux_2331_nl;
  assign mux_2331_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00052_ : mux_tmp_2324;
  assign mux_2327_nl = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2319 : mux_2326_nl;
  assign mux_2326_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00051_ : mux_tmp_2319;
  assign mux_2320_nl = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2312 : mux_2319_nl;
  assign mux_2319_nl = cfg_proc_precision_1_sva_st_102[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00050_ : mux_tmp_2312;
  assign mux_2314_nl = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2306 : mux_2313_nl;
  assign mux_2313_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00049_ : mux_tmp_2306;
  assign mux_2308_nl = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2300 : mux_2307_nl;
  assign mux_2307_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00048_ : mux_tmp_2300;
  assign mux_2302_nl = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2294 : mux_2301_nl;
  assign mux_2301_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00047_ : mux_tmp_2294;
  assign mux_tmp_2353 = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2351 : mux_2358_nl;
  assign mux_2358_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00056_ : mux_tmp_2351;
  assign mux_tmp_2351 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : mux_2356_nl;
  assign mux_2356_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00056_ : and_2136_cse;
  assign mux_tmp_2347 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2345 : mux_2352_nl;
  assign mux_2352_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00055_ : mux_tmp_2345;
  assign mux_tmp_2345 = or_3542_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2350_nl : _00055_;
  assign mux_2350_nl = or_5254_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : _00055_;
  assign mux_tmp_2341 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2339 : mux_2346_nl;
  assign mux_2346_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00054_ : mux_tmp_2339;
  assign mux_tmp_2339 = or_3542_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : _00054_;
  assign mux_tmp_2336 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2334 : mux_2341_nl;
  assign mux_2341_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00051_ : mux_tmp_2334;
  assign mux_tmp_2334 = or_3542_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2315 : _00051_;
  assign mux_tmp_2330 = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2328 : mux_2335_nl;
  assign mux_2335_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00053_ : mux_tmp_2328;
  assign mux_tmp_2328 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : mux_2333_nl;
  assign mux_2333_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00053_ : and_2136_cse;
  assign mux_tmp_2324 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2322 : mux_2329_nl;
  assign mux_2329_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00052_ : mux_tmp_2322;
  assign mux_tmp_2322 = or_3542_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : _00052_;
  assign mux_tmp_2319 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2317 : mux_2324_nl;
  assign mux_2324_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00051_ : mux_tmp_2317;
  assign mux_tmp_2317 = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2315 : mux_2322_nl;
  assign mux_2322_nl = cfg_proc_precision_1_sva_st_102[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00051_ : mux_tmp_2315;
  assign mux_tmp_2315 = or_5254_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : _00051_;
  assign mux_tmp_2312 = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2310 : mux_2317_nl;
  assign mux_2317_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00050_ : mux_tmp_2310;
  assign mux_tmp_2310 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : mux_2315_nl;
  assign mux_2315_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00050_ : and_2136_cse;
  assign mux_tmp_2306 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2304 : mux_2311_nl;
  assign mux_2311_nl = cfg_proc_precision_1_sva_st_66[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00049_ : mux_tmp_2304;
  assign mux_tmp_2304 = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : mux_2309_nl;
  assign mux_2309_nl = cfg_proc_precision_1_sva_st_102[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00049_ : and_2136_cse;
  assign mux_tmp_2300 = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2298 : mux_2305_nl;
  assign mux_2305_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00048_ : mux_tmp_2298;
  assign mux_tmp_2298 = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : mux_2303_nl;
  assign mux_2303_nl = cfg_proc_precision_1_sva_st_102[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00048_ : and_2136_cse;
  assign mux_tmp_2294 = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2136_cse : mux_2299_nl;
  assign mux_2299_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00047_ : and_2136_cse;
  assign mux_2208_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2207_nl : or_tmp_3832;
  assign mux_2207_nl = or_4714_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4675_nl : or_tmp_3832;
  assign mux_tmp_2203 = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2205_nl : or_tmp_3826;
  assign mux_2205_nl = or_4714_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2204_nl : or_tmp_3826;
  assign mux_2204_nl = or_4667_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3826 : mux_2203_nl;
  assign mux_2203_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2201_nl : mux_2202_nl;
  assign mux_2202_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2040_cse : or_tmp_3826;
  assign mux_2201_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2200_nl : or_tmp_3826;
  assign mux_2200_nl = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2040_cse : fsm_output[1];
  assign mux_1964_nl = and_2145_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1953_nl = and_2146_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1943_nl = and_2147_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1940_nl = and_2148_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1927_nl = and_2150_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1903_nl = and_2152_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1876_nl = and_2155_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1846_nl = and_2157_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1836_nl = and_2158_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1966_itm = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_unequal_tmp_20 : cvt_unequal_tmp_21;
  assign mux_tmp_1899 = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_165 : nor_1025_nl;
  assign not_tmp_2422 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1839_nl : mux_1841_nl;
  assign mux_1841_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1053_nl : or_1157_cse;
  assign mux_1839_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_57_cse : nor_2099_cse;
  assign mux_tmp_1813 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_225 : nor_1063_nl;
  assign mux_tmp_1622 = cvt_1_FpMantRNE_24U_11U_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1618 = cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1614 = cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1610 = cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1606 = cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1600 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : nand_230_nl;
  assign mux_tmp_1596 = cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1592 = cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1586 = cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1582 = cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1578 = cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1574 = cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1570 = cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1566 = cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_6 : or_tmp_24;
  assign mux_tmp_1469 = or_2306_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : and_306_nl;
  assign mux_tmp_1435 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : mux_1434_nl;
  assign mux_1434_nl = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1433_nl : nor_1320_cse;
  assign mux_1433_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1432_nl : or_tmp_2136;
  assign mux_1432_nl = or_4714_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1431_nl : or_tmp_2136;
  assign mux_1431_nl = or_400_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1430_nl : or_tmp_2136;
  assign mux_1430_nl = cfg_out_precision_1_sva_st_149[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : and_2246_cse;
  assign mux_tmp_1419 = or_1198_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1418_nl : or_2246_nl;
  assign mux_1418_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1417_nl : or_5189_cse;
  assign mux_1417_nl = or_4714_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1416_nl : or_5189_cse;
  assign mux_1416_nl = or_400_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_2245_nl : or_5189_cse;
  assign mux_tmp_1409 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : mux_1408_nl;
  assign mux_1408_nl = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1407_nl : nor_1320_cse;
  assign mux_1407_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1406_nl : or_tmp_2136;
  assign mux_1406_nl = or_4714_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1405_nl : or_tmp_2136;
  assign mux_1405_nl = or_2232_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : and_2246_cse;
  assign mux_tmp_1337 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_1 : mux_1494_cse;
  assign mux_tmp_1332 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : mux_1331_nl;
  assign mux_1331_nl = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1330_nl : nor_1320_cse;
  assign mux_1330_nl = or_2140_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : mux_1329_nl;
  assign mux_1329_nl = cfg_out_precision_1_sva_st_149[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00044_ : or_tmp_2136;
  assign mux_1328_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1326 : mux_1327_nl;
  assign mux_1327_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00042_ : mux_tmp_1326;
  assign mux_tmp_1326 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1270 : mux_1325_nl;
  assign mux_1325_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00042_ : mux_tmp_1270;
  assign mux_tmp_1280 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_1 : mux_1464_cse;
  assign mux_tmp_1276 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : mux_1275_nl;
  assign mux_1275_nl = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1274_nl : nor_1320_cse;
  assign mux_1274_nl = or_2140_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2136 : mux_1273_nl;
  assign mux_1273_nl = cfg_out_precision_1_sva_st_149[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00043_ : or_tmp_2136;
  assign mux_1272_nl = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1270 : mux_1271_nl;
  assign mux_1271_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00042_ : mux_tmp_1270;
  assign mux_tmp_1270 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2139 : mux_1269_nl;
  assign mux_1269_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00042_ : or_tmp_2139;
  assign mux_tmp_1264 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_94 : and_283_cse;
  assign mux_tmp_1227 = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1226 : nor_1373_nl;
  assign mux_tmp_1226 = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1225 : nor_1372_nl;
  assign mux_tmp_1225 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_3 : nor_1371_nl;
  assign mux_tmp_1197 = cfg_proc_precision_1_sva_st_66[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1196 : nor_1388_nl;
  assign mux_tmp_1196 = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3538_cse : nor_1387_nl;
  assign mux_tmp_1152 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1041 : mux_1151_nl;
  assign mux_1151_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00040_ : mux_tmp_1041;
  assign mux_tmp_1111 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1109 : mux_1110_nl;
  assign mux_1110_nl = reg_cfg_proc_precision_1_sva_st_40_cse[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00041_ : mux_tmp_1109;
  assign mux_tmp_1105 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1103 : mux_1104_nl;
  assign mux_1104_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00041_ : mux_tmp_1103;
  assign mux_tmp_1103 = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1101 : mux_1102_nl;
  assign mux_1102_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00041_ : mux_tmp_1101;
  assign mux_tmp_1101 = or_1773_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1109 : nor_1446_nl;
  assign mux_tmp_1100 = or_1774_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_987 : nor_1486_cse;
  assign mux_tmp_1088 = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1087_nl : mux_976_nl;
  assign mux_976_nl = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_169 : mux_tmp_962;
  assign mux_1087_nl = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1086_nl : mux_tmp_962;
  assign mux_1086_nl = or_1745_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_169 : nor_1455_nl;
  assign mux_tmp_1074 = or_1918_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_963 : mux_1073_nl;
  assign mux_1073_nl = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1072_nl : mux_tmp_962;
  assign mux_1072_nl = or_1919_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_168 : nor_1464_nl;
  assign mux_tmp_1049 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1047 : mux_1048_nl;
  assign mux_1048_nl = reg_cfg_proc_precision_1_sva_st_40_cse[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00040_ : mux_tmp_1047;
  assign mux_tmp_1043 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1041 : mux_1042_nl;
  assign mux_1042_nl = cfg_proc_precision_1_sva_st_89[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00040_ : mux_tmp_1041;
  assign mux_tmp_1041 = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1039 : mux_1040_nl;
  assign mux_1040_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00040_ : mux_tmp_1039;
  assign mux_tmp_1039 = or_1643_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1047 : nor_1487_nl;
  assign mux_tmp_1038 = or_1644_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_987 : nor_1486_cse;
  assign mux_tmp_1015 = _07544_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_947 : mux_1014_nl;
  assign mux_1014_nl = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1013_nl : mux_tmp_946;
  assign mux_1013_nl = or_1919_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_165 : and_2247_nl;
  assign mux_tmp_994 = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_987 : mux_989_cse;
  assign mux_tmp_992 = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1142_cse : mux_tmp_944;
  assign mux_tmp_987 = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_986 : nor_1535_nl;
  assign mux_tmp_986 = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nor_1534_nl;
  assign mux_969_nl = cfg_proc_precision_1_sva_st_102[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1159_cse : nor_1545_nl;
  assign mux_tmp_963 = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_168 : mux_tmp_962;
  assign mux_tmp_962 = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_79 : and_tmp_19;
  assign mux_tmp_961 = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_79 : mux_tmp_960;
  assign mux_tmp_960 = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_123 : and_2186_cse;
  assign mux_tmp_947 = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_165 : mux_tmp_946;
  assign mux_tmp_946 = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_50 : and_1386_cse;
  assign mux_tmp_945 = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_50 : mux_tmp_944;
  assign mux_tmp_944 = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_12 : and_2186_cse;
  assign mux_tmp_766 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_765 : nor_1686_nl;
  assign mux_tmp_765 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_658 : nor_1685_nl;
  assign not_tmp_989 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1687_nl : nor_1689_nl;
  assign mux_tmp_743 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_742 : nor_1702_nl;
  assign mux_tmp_742 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_741 : nor_1701_nl;
  assign mux_tmp_741 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_740 : nor_1700_nl;
  assign mux_tmp_740 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_739 : nor_1699_nl;
  assign mux_tmp_739 = IsNaN_5U_10U_nor_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : mux_738_nl;
  assign mux_738_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2194_cse : main_stage_v_2;
  assign mux_tmp_727 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_726 : nor_1714_nl;
  assign mux_tmp_726 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_725 : nor_1713_nl;
  assign mux_tmp_725 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_724 : nor_1712_nl;
  assign mux_tmp_724 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_723 : nor_1711_nl;
  assign mux_tmp_723 = or_1072_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : and_2194_cse;
  assign mux_tmp_720 = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_719 : nor_1719_nl;
  assign mux_tmp_719 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1489_cse : nor_1718_nl;
  assign not_tmp_899 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1728_nl : nor_1730_nl;
  assign mux_tmp_695 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_694 : nor_1740_nl;
  assign mux_tmp_694 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_693 : nor_1739_nl;
  assign mux_tmp_693 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_692 : nor_1738_nl;
  assign mux_tmp_692 = IsNaN_5U_10U_nor_14_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : mux_691_nl;
  assign mux_691_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2199_cse : main_stage_v_2;
  assign mux_tmp_681 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_680 : nor_1750_nl;
  assign mux_tmp_680 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_679 : nor_1749_nl;
  assign mux_tmp_679 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_678 : nor_1748_nl;
  assign mux_tmp_678 = or_1015_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : and_2199_cse;
  assign mux_tmp_658 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : nor_1762_nl;
  assign not_tmp_811 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1764_nl : nor_1766_nl;
  assign mux_tmp_641 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_640 : nor_1776_nl;
  assign mux_tmp_640 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_639 : nor_1775_nl;
  assign mux_tmp_639 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_638 : nor_1774_nl;
  assign mux_tmp_638 = IsNaN_5U_10U_nor_1_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : mux_637_nl;
  assign mux_637_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2202_nl : main_stage_v_2;
  assign mux_tmp_634 = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1489_cse : nor_1780_nl;
  assign not_tmp_757 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1787_nl : nor_1789_nl;
  assign mux_tmp_614 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_613 : nor_1796_nl;
  assign mux_tmp_613 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_612 : nor_1795_nl;
  assign mux_tmp_612 = IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : mux_611_nl;
  assign mux_611_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2206_cse : main_stage_v_2;
  assign mux_tmp_602 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_601 : nor_1804_nl;
  assign mux_tmp_601 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_600 : nor_1803_nl;
  assign mux_tmp_600 = or_921_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : and_2206_cse;
  assign mux_tmp_597 = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1460_cse : nor_1807_nl;
  assign mux_tmp_592 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_591 : nor_1810_nl;
  assign mux_tmp_591 = IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_400_cse_1 : and_2208_nl;
  assign mux_tmp_585 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_894_nl : or_898_nl;
  assign mux_tmp_580 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_579 : nor_1817_nl;
  assign mux_tmp_579 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_578 : nor_1816_nl;
  assign mux_tmp_578 = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_577 : nor_1815_nl;
  assign mux_tmp_577 = IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : mux_576_nl;
  assign mux_576_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2209_nl : main_stage_v_2;
  assign mux_tmp_566 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_565 : nor_1827_nl;
  assign mux_tmp_565 = or_871_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_298 : and_2210_nl;
  assign mux_tmp_560 = cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_305 : nor_1828_nl;
  assign not_tmp_638 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1838_nl : nor_1840_nl;
  assign mux_tmp_541 = IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_311 : mux_540_nl;
  assign mux_540_nl = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_538_nl : mux_tmp_311;
  assign mux_538_nl = IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_311 : _00037_;
  assign mux_tmp_525 = IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_298 : mux_524_nl;
  assign mux_524_nl = or_828_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2214_nl : mux_tmp_298;
  assign mux_tmp_519 = cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_1851_nl;
  assign not_tmp_580 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1858_nl : nor_1860_nl;
  assign mux_tmp_502 = or_795_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_311 : mux_500_nl;
  assign mux_500_nl = IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_311 : _00037_;
  assign mux_tmp_487 = IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_298 : mux_486_nl;
  assign mux_486_nl = or_784_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2218_nl : mux_tmp_298;
  assign mux_tmp_481 = cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_1872_nl;
  assign not_tmp_520 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1882_nl : nor_1884_nl;
  assign mux_tmp_455 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_1891_nl;
  assign not_tmp_497 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1892_nl : nor_1894_nl;
  assign mux_tmp_441 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_440 : nor_1902_nl;
  assign mux_tmp_440 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_298 : nor_1901_nl;
  assign mux_tmp_435 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_305 : nor_1906_nl;
  assign mux_tmp_428 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_427 : nor_1911_nl;
  assign mux_tmp_427 = or_690_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_184_nl : mux_tmp_298;
  assign mux_tmp_422 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_421 : nor_1915_nl;
  assign mux_tmp_421 = cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_1912_nl;
  assign mux_tmp_416 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_415 : nor_1919_nl;
  assign mux_tmp_415 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_400_cse_1 : _00039_;
  assign not_tmp_436 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1922_nl : nor_1924_nl;
  assign mux_tmp_405 = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_404_nl : mux_tmp_311;
  assign mux_404_nl = or_4536_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_311 : _00037_;
  assign mux_tmp_391 = or_645_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_181_nl : mux_tmp_298;
  assign mux_tmp_386 = cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_1935_nl;
  assign not_tmp_388 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1942_nl : nor_1944_nl;
  assign mux_tmp_370 = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_369_nl : mux_tmp_311;
  assign mux_369_nl = or_600_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_311 : _00037_;
  assign mux_tmp_356 = or_599_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_176_nl : mux_tmp_298;
  assign mux_tmp_351 = cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_1955_nl;
  assign mux_tmp_345 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_400_cse_1 : nor_1959_nl;
  assign not_tmp_336 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1964_nl : nor_1966_nl;
  assign mux_tmp_321 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_50 : nor_1974_nl;
  assign not_tmp_312 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1975_nl : nor_1977_nl;
  assign mux_tmp_317 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_183_cse_1 : _00038_;
  assign mux_tmp_313 = or_461_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_312_nl : mux_tmp_311;
  assign mux_312_nl = or_510_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_311 : _00037_;
  assign mux_tmp_311 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_309 : mux_310_nl;
  assign mux_310_nl = cfg_proc_precision_1_sva_st_101[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00037_ : mux_tmp_309;
  assign mux_tmp_309 = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : mux_308_nl;
  assign mux_308_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00037_ : main_stage_v_2;
  assign mux_tmp_305 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_1983_nl;
  assign mux_tmp_299 = or_520_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_167_nl : mux_tmp_298;
  assign mux_tmp_298 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_239 : nor_1987_nl;
  assign mux_tmp_294 = cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_259 : nor_1988_nl;
  assign not_tmp_269 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1995_nl : nor_1997_nl;
  assign not_tmp_249 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2007_nl : nor_2009_nl;
  assign mux_tmp_263 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_239 : nor_2013_nl;
  assign mux_tmp_259 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_236 : nor_2015_nl;
  assign mux_tmp_253 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_251 : mux_252_nl;
  assign mux_252_nl = or_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_52 : main_stage_v_2;
  assign mux_tmp_251 = or_445_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_152_nl : and_153_nl;
  assign mux_250_nl = cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_249 : _00036_;
  assign mux_tmp_249 = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_448_nl : _00036_;
  assign mux_tmp_245 = or_1198_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_434_nl : mux_244_nl;
  assign mux_244_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_429_nl : or_431_nl;
  assign mux_tmp_239 = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : nor_2021_nl;
  assign mux_tmp_236 = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_1 : nor_2022_nl;
  assign mux_tmp_200 = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_199 : nor_2028_nl;
  assign mux_tmp_199 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : nor_2027_nl;
  assign mux_tmp_189 = _04006_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_378_nl : nand_nl;
  assign mux_188_nl = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_4 : nor_2029_nl;
  assign mux_tmp_161 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_1 : main_stage_v_2;
  assign mux_tmp_151 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_33 : nor_2049_nl;
  assign mux_148_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_117 : nor_2050_nl;
  assign mux_tmp_129 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_19 : nor_2052_nl;
  assign mux_tmp_123 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_120 : nor_2054_nl;
  assign mux_tmp_122 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_tmp_18;
  assign mux_tmp_120 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4550_cse : nor_2055_nl;
  assign mux_tmp_117 = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_12 : nor_2056_nl;
  assign mux_tmp_114 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_tmp_11;
  assign mux_110_cse = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_186_cse : mux_109_nl;
  assign mux_109_nl = reg_cfg_proc_precision_1_sva_st_40_cse[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_8_cse : or_186_cse;
  assign mux_tmp_39 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_86_nl;
  assign mux_tmp_6 = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_19 : or_23_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_1_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_27_0_1[9:0] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_2_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_59_31_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_3_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_91_63_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_4_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_123_95_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_5_mx0 = or_tmp_2469 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1 : chn_idata_data_sva_1_155_127_1[10:1];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_6_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_187_159_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_7_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_219_191_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_8_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_251_223_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_9_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_283_255_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_10_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_315_287_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_11_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_347_319_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_12_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_379_351_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_13_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_411_383_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_14_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_443_415_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_15_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_475_447_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_5_mx0 = IsNaN_8U_23U_land_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) chn_idata_data_sva_1_507_479_1[10:1] : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1;
  assign FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0 = chn_idata_data_sva_2_511_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0 = chn_idata_data_sva_2_495_479_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0 = chn_idata_data_sva_2_463_447_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0 = chn_idata_data_sva_2_431_415_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0 = chn_idata_data_sva_2_399_383_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0 = chn_idata_data_sva_2_367_351_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0 = chn_idata_data_sva_2_335_319_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0 = chn_idata_data_sva_2_303_287_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0 = chn_idata_data_sva_2_271_255_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0 = chn_idata_data_sva_2_239_223_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0 = chn_idata_data_sva_2_207_191_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0 = chn_idata_data_sva_2_175_159_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0 = chn_idata_data_sva_2_143_127_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0 = chn_idata_data_sva_2_111_95_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0 = chn_idata_data_sva_2_79_63_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0 = chn_idata_data_sva_2_47_31_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24490|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24489" *) 16'b1000000000000000 : 16'b0111111111111111;
  assign FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1;
  assign FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg;
  assign FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1 = FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : reg_chn_idata_data_sva_3_15_0_2_reg;
  assign _00170_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_22_nl;
  assign _00169_ = _07252_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[24:1] : 24'b111111111111111111111111;
  assign _00168_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  assign _00167_ = _07221_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[24:1] : 24'b111111111111111111111111;
  assign _00166_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  assign _00165_ = _07190_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[24:1] : 24'b111111111111111111111111;
  assign _00164_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  assign _00163_ = _07159_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[24:1] : 24'b111111111111111111111111;
  assign _00162_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  assign _00161_ = _07128_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[24:1] : 24'b111111111111111111111111;
  assign _00160_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  assign _00159_ = _07097_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[24:1] : 24'b111111111111111111111111;
  assign _00158_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  assign _00157_ = _07066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[24:1] : 24'b111111111111111111111111;
  assign _00156_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  assign _00155_ = _07035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[24:1] : 24'b111111111111111111111111;
  assign _00154_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  assign _00153_ = _07004_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[24:1] : 24'b111111111111111111111111;
  assign _00152_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  assign _00151_ = _06973_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[24:1] : 24'b111111111111111111111111;
  assign _00150_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  assign _00149_ = _06942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[24:1] : 24'b111111111111111111111111;
  assign _00148_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  assign _00147_ = _06911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[24:1] : 24'b111111111111111111111111;
  assign _00146_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  assign _00145_ = _06880_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[24:1] : 24'b111111111111111111111111;
  assign _00144_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  assign _00143_ = _06849_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[24:1] : 24'b111111111111111111111111;
  assign _00142_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  assign _00141_ = _06818_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[24:1] : 24'b111111111111111111111111;
  assign _00140_ = IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) 24'b111111111111111111111111 : cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_2_nl;
  assign _00139_ = _06787_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24507|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24506" *) IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[24:1] : 24'b111111111111111111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_47_nl = cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9[4] : _00035_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_46_nl = cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9[4] : _00034_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_45_nl = cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9[4] : _00033_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_44_nl = cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9[4] : _00032_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_43_nl = cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9[4] : _00031_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_42_nl = cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9[4] : _00030_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_41_nl = cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9[4] : _00029_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_40_nl = cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9[4] : _00028_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_39_nl = cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9[4] : _00027_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_38_nl = cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9[4] : _00026_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_37_nl = cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9[4] : _00025_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_36_nl = cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9[4] : _00024_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_35_nl = cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9[4] : _00023_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_34_nl = cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9[4] : _00022_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_33_nl = cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9[4] : _00021_;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_32_nl = cvt_1_FpMantRNE_24U_11U_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9[4] : _00020_;
  assign FpIntToFloat_17U_5U_10U_else_mux_46_nl = FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_15 : or_5086_cse;
  assign FpMantRNE_17U_11U_else_mux_31_nl = or_3999_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpMantRNE_17U_11U_else_and_4_svs : cvt_16_FpMantRNE_17U_11U_else_and_4_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0 = cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_16_FpMantRNE_17U_11U_else_acc_4_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_43_nl = FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_14 : or_5069_cse;
  assign FpMantRNE_17U_11U_else_mux_29_nl = or_3989_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpMantRNE_17U_11U_else_and_3_svs : cvt_15_FpMantRNE_17U_11U_else_and_3_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0 = cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_15_FpMantRNE_17U_11U_else_acc_3_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_40_nl = FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_13 : or_5053_cse;
  assign FpMantRNE_17U_11U_else_mux_27_nl = or_3977_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpMantRNE_17U_11U_else_and_3_svs : cvt_14_FpMantRNE_17U_11U_else_and_3_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0 = cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_14_FpMantRNE_17U_11U_else_acc_3_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_37_nl = FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_12 : or_5038_cse;
  assign FpMantRNE_17U_11U_else_mux_25_nl = or_3965_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpMantRNE_17U_11U_else_and_2_svs : cvt_13_FpMantRNE_17U_11U_else_and_2_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0 = cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_13_FpMantRNE_17U_11U_else_acc_2_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_34_nl = FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_11 : or_1925_cse_1;
  assign FpMantRNE_17U_11U_else_mux_23_nl = or_3953_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpMantRNE_17U_11U_else_and_3_svs : cvt_12_FpMantRNE_17U_11U_else_and_3_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0 = cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_12_FpMantRNE_17U_11U_else_acc_3_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_31_nl = FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_10 : or_1892_cse_1;
  assign FpMantRNE_17U_11U_else_mux_21_nl = or_3942_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpMantRNE_17U_11U_else_and_2_svs : cvt_11_FpMantRNE_17U_11U_else_and_2_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0 = cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_11_FpMantRNE_17U_11U_else_acc_2_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_28_nl = FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_9 : or_1851_cse_1;
  assign FpMantRNE_17U_11U_else_mux_19_nl = or_3932_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpMantRNE_17U_11U_else_and_2_svs : cvt_10_FpMantRNE_17U_11U_else_and_2_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0 = cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_10_FpMantRNE_17U_11U_else_acc_2_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_22_nl = FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_7 : or_1789_cse_1;
  assign FpMantRNE_17U_11U_else_mux_15_nl = or_3911_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpMantRNE_17U_11U_else_and_3_svs : cvt_8_FpMantRNE_17U_11U_else_and_3_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0 = cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_8_FpMantRNE_17U_11U_else_acc_3_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_19_nl = FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_6 : or_1752_cse_1;
  assign FpMantRNE_17U_11U_else_mux_13_nl = or_3900_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpMantRNE_17U_11U_else_and_2_svs : cvt_7_FpMantRNE_17U_11U_else_and_2_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0 = cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_7_FpMantRNE_17U_11U_else_acc_2_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_16_nl = FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_5 : or_1720_cse_1;
  assign FpMantRNE_17U_11U_else_mux_11_nl = or_3891_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpMantRNE_17U_11U_else_and_2_svs : cvt_6_FpMantRNE_17U_11U_else_and_2_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0 = cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_6_FpMantRNE_17U_11U_else_acc_2_nl;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0 = cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_5_FpMantRNE_17U_11U_else_acc_1_nl;
  assign FpIntToFloat_17U_5U_10U_else_mux_10_nl = FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_else_unequal_tmp_3 : or_1659_cse_1;
  assign FpMantRNE_17U_11U_else_mux_7_nl = or_3872_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpMantRNE_17U_11U_else_and_2_svs : cvt_4_FpMantRNE_17U_11U_else_and_2_tmp;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0 = cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_4_FpMantRNE_17U_11U_else_acc_2_nl;
  assign cvt_else_equal_tmp_36_mx0 = or_dcpl_195 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 : cvt_else_equal_tmp;
  assign cvt_else_equal_tmp_37_mx0 = or_dcpl_195 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 : cvt_else_equal_tmp_1;
  assign cvt_else_mux_59_nl = and_1059_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_46 : cvt_else_equal_tmp_1;
  assign cvt_else_mux_62_nl = and_1059_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_45 : cvt_else_equal_tmp;
  assign cvt_else_mux_56_nl = and_1059_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs_15 : cvt_else_nor_dfs;
  assign cvt_else_equal_tmp_42_mx0 = and_tmp_248 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  assign cvt_else_equal_tmp_43_mx0 = and_tmp_248 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  assign cvt_else_nor_dfs_14_mx1 = and_tmp_248 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs : cvt_else_nor_dfs_15;
  assign cvt_else_equal_tmp_39_mx1 = or_dcpl_197 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_45 : cvt_else_equal_tmp;
  assign cvt_else_equal_tmp_40_mx1 = or_dcpl_197 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_46 : cvt_else_equal_tmp_1;
  assign cvt_else_nor_dfs_13_mx1 = or_dcpl_197 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs_15 : cvt_else_nor_dfs;
  assign cvt_else_equal_tmp_30_mx0 = mux_tmp_987 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  assign cvt_else_equal_tmp_31_mx0 = mux_tmp_987 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  assign cvt_else_nor_dfs_10_mx1 = mux_tmp_987 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs : cvt_else_nor_dfs_10;
  assign cvt_else_equal_tmp_33_mx1 = or_dcpl_197 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_33 : cvt_else_equal_tmp;
  assign cvt_else_equal_tmp_34_mx1 = or_dcpl_197 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_34 : cvt_else_equal_tmp_1;
  assign cvt_else_nor_dfs_11_mx1 = or_dcpl_197 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs_11 : cvt_else_nor_dfs;
  assign cvt_else_equal_tmp_27_mx0 = or_dcpl_195 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 : cvt_else_equal_tmp;
  assign cvt_else_equal_tmp_28_mx1 = or_dcpl_195 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_28 : cvt_else_equal_tmp_1;
  assign cvt_else_nor_dfs_9_mx1 = or_dcpl_195 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_cvt_else_nor_dfs_9_cse : cvt_else_nor_dfs;
  assign cvt_else_equal_tmp_18_mx0 = mux_tmp_1899 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  assign cvt_else_equal_tmp_19_mx0 = mux_tmp_1899 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  assign cvt_else_nor_dfs_6_mx1 = mux_tmp_1899 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs : cvt_else_nor_dfs_10;
  assign cvt_else_equal_tmp_21_mx1 = or_dcpl_188 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_33 : cvt_else_equal_tmp;
  assign cvt_else_equal_tmp_22_mx1 = or_dcpl_188 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_34 : cvt_else_equal_tmp_1;
  assign cvt_else_nor_dfs_7_mx1 = or_dcpl_188 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs_11 : cvt_else_nor_dfs;
  assign cvt_else_equal_tmp_15_mx0 = or_dcpl_184 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 : cvt_else_equal_tmp;
  assign cvt_else_equal_tmp_16_mx1 = or_dcpl_184 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_16 : cvt_else_equal_tmp_1;
  assign cvt_else_nor_dfs_5_mx1 = or_dcpl_184 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs_10 : cvt_else_nor_dfs;
  assign cvt_else_equal_tmp_9_mx1 = or_dcpl_181 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_9 : cvt_else_equal_tmp;
  assign cvt_else_equal_tmp_10_mx0 = or_dcpl_181 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 : cvt_else_equal_tmp_1;
  assign cvt_else_nor_dfs_3_mx1 = or_dcpl_181 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs_10 : cvt_else_nor_dfs;
  assign cvt_else_equal_tmp_3_mx0 = _01591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  assign cvt_else_equal_tmp_4_mx1 = _01591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : cvt_else_equal_tmp_5;
  assign cvt_else_nor_dfs_1_mx1 = _01591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_nor_dfs : cvt_else_nor_dfs_2;
  assign _00138_ = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_22_nl;
  assign _00137_ = _04873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[15:1] : 15'b111111111111111;
  assign _00136_ = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  assign _00135_ = _04871_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1] : 15'b111111111111111;
  assign _00134_ = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  assign _00133_ = _04869_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1] : 15'b111111111111111;
  assign _00132_ = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  assign _00131_ = _04868_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1] : 15'b111111111111111;
  assign _00130_ = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  assign _00129_ = _04866_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1] : 15'b111111111111111;
  assign _00128_ = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  assign _00127_ = _04865_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1] : 15'b111111111111111;
  assign _00126_ = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  assign _00125_ = _04864_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1] : 15'b111111111111111;
  assign _00124_ = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  assign _00123_ = _05324_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1] : 15'b111111111111111;
  assign _00122_ = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  assign _00121_ = _04863_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1] : 15'b111111111111111;
  assign _00120_ = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  assign _00119_ = _04861_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1] : 15'b111111111111111;
  assign _00118_ = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  assign _00117_ = _04860_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1] : 15'b111111111111111;
  assign _00116_ = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  assign _00115_ = _04859_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1] : 15'b111111111111111;
  assign _00114_ = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  assign _00113_ = _04857_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1] : 15'b111111111111111;
  assign _00112_ = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  assign _00111_ = _05320_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1] : 15'b111111111111111;
  assign _00110_ = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  assign _00109_ = _05319_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1] : 15'b111111111111111;
  assign _00108_ = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) 15'b111111111111111 : cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_2_nl;
  assign _00107_ = _05318_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[15:1] : 15'b111111111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_30_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_30_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_15_nl;
  assign _00106_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_nl;
  assign _00105_ = _03839_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_181_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_181_nl = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_16_FpMantRNE_24U_11U_else_acc_4_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_15_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_28_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_28_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_14_nl;
  assign _00104_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_nl;
  assign _00103_ = _03838_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_169_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_169_nl = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_15_FpMantRNE_24U_11U_else_acc_3_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_14_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_26_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_26_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_13_nl;
  assign _00102_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_nl;
  assign _00101_ = _03837_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_157_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_157_nl = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_14_FpMantRNE_24U_11U_else_acc_3_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_13_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_24_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_24_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_12_nl;
  assign _00100_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_nl;
  assign _00099_ = _03836_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_145_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_145_nl = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_13_FpMantRNE_24U_11U_else_acc_2_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_12_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_22_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_22_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_11_nl;
  assign _00098_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_nl;
  assign _00097_ = _03835_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_133_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_133_nl = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_12_FpMantRNE_24U_11U_else_acc_3_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_11_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_20_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_20_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_10_nl;
  assign _00096_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_nl;
  assign _00095_ = _03834_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_121_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_121_nl = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_11_FpMantRNE_24U_11U_else_acc_2_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_10_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_18_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_18_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_9_nl;
  assign _00094_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_nl;
  assign _00093_ = _03833_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_109_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_109_nl = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_10_FpMantRNE_24U_11U_else_acc_2_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_9_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_16_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_16_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_8_nl;
  assign _00092_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_nl;
  assign _00091_ = _03832_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_97_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_97_nl = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_9_FpMantRNE_24U_11U_else_acc_1_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_8_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_14_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_14_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_7_nl;
  assign _00090_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_nl;
  assign _00089_ = _03831_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_85_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_85_nl = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_8_FpMantRNE_24U_11U_else_acc_3_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_7_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_12_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_12_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_6_nl;
  assign _00088_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_nl;
  assign _00087_ = _03830_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_73_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_73_nl = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_7_FpMantRNE_24U_11U_else_acc_2_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_6_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_10_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_10_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_5_nl;
  assign _00086_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_nl;
  assign _00085_ = _03829_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_61_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_61_nl = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_6_FpMantRNE_24U_11U_else_acc_2_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0 = or_tmp_2469 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_8_nl : 4'b1111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_8_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_4_nl;
  assign _00084_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_nl;
  assign _00083_ = _03828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_49_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_49_nl = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_5_FpMantRNE_24U_11U_else_acc_1_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_4_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_6_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_6_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_3_nl;
  assign _00082_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_nl;
  assign _00081_ = _03827_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_37_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_37_nl = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_4_FpMantRNE_24U_11U_else_acc_2_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_3_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_4_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_4_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_2_nl;
  assign _00080_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl;
  assign _00079_ = _03826_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_25_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_25_nl = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_3_FpMantRNE_24U_11U_else_acc_1_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_2_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_2_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_2_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_1_nl;
  assign _00078_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_nl;
  assign _00077_ = _03825_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_13_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_13_nl = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_2_FpMantRNE_24U_11U_else_acc_1_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0 = IsNaN_8U_23U_land_1_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b1111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24541|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24540" *) 4'b0000 : FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl;
  assign _00076_ = FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b1111111111 : FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl;
  assign _00075_ = _03824_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl : 10'b1111111111;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) cvt_1_FpMantRNE_24U_11U_else_acc_nl : FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[9:0];
  assign mux_134_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_243_nl;
  assign mux_125_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_226_nl;
  assign mux_119_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_213 : or_217_nl;
  assign mux_1286_nl = or_3623_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1276 : mux_1285_nl;
  assign mux_1285_nl = cfg_out_precision_1_sva_st_154[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00019_ : mux_tmp_1276;
  assign mux_1284_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1280 : mux_1283_nl;
  assign mux_1283_nl = reg_cfg_proc_precision_1_sva_st_40_cse[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00018_ : mux_tmp_1280;
  assign mux_377_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : or_626_nl;
  assign mux_320_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : or_547_nl;
  assign mux_272_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_5379_cse : or_479_nl;
  assign mux_1654_cse = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1489_cse : mux_1653_nl;
  assign mux_1653_nl = cfg_proc_precision_1_sva_st_64[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1185_cse : mux_1489_cse;
  assign mux_1626_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1195_nl : nor_1556_cse;
  assign mux_152_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : mux_tmp_151;
  assign mux_149_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_tmp_33;
  assign mux_118_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_tmp_16;
  assign mux_133_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_1386_cse;
  assign mux_130_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : mux_tmp_129;
  assign mux_124_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_tmp_19;
  assign mux_1521_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1519_nl : mux_1436_cse;
  assign mux_1519_nl = or_2289_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1271_nl : main_stage_v_1;
  assign mux_1495_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1490_nl : mux_1494_cse;
  assign mux_1490_nl = or_2289_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2110_nl : main_stage_v_1;
  assign mux_1489_cse = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1460_cse : nor_1287_nl;
  assign mux_1494_cse = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2127_nl : main_stage_v_2;
  assign mux_1466_cse = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_1 : nor_1301_nl;
  assign mux_1465_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1461_nl : mux_1464_cse;
  assign mux_1461_nl = or_2289_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2114_nl : main_stage_v_1;
  assign mux_1460_cse = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1466_cse : nor_1305_nl;
  assign mux_1464_cse = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2130_nl : main_stage_v_2;
  assign mux_1463_cse = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_658 : nor_1306_nl;
  assign mux_1458_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1309_cse : nor_1310_cse;
  assign mux_1442_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1441_nl : mux_tmp_1435;
  assign mux_1441_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1439_nl : mux_tmp_1435;
  assign mux_1439_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1435 : mux_1438_nl;
  assign mux_1438_nl = cfg_out_precision_1_sva_st_154[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00067_ : mux_tmp_1435;
  assign mux_1437_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_1 : mux_1436_cse;
  assign mux_1436_cse = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1314_nl : main_stage_v_2;
  assign mux_1345_nl = or_3623_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1332 : mux_1344_nl;
  assign mux_1344_nl = cfg_out_precision_1_sva_st_154[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00074_ : mux_tmp_1332;
  assign mux_1343_nl = reg_cfg_proc_precision_1_sva_st_40_cse[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1337 : mux_1342_nl;
  assign mux_1342_nl = reg_cfg_proc_precision_1_sva_st_40_cse[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00045_ : mux_tmp_1337;
  assign mux_2020_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3606_nl : mux_2019_nl;
  assign mux_2019_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3607_nl : mux_2018_nl;
  assign mux_2018_nl = or_1159_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : or_3609_nl;
  assign mux_2017_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_1198_cse : or_4709_cse;
  assign mux_2015_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3597_nl : mux_2014_nl;
  assign mux_2014_nl = or_1159_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2013_nl : mux_2012_nl;
  assign mux_2013_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3600_nl : cfg_mode_eql_1_sva_6;
  assign mux_2012_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : or_1176_cse;
  assign mux_2011_nl = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_out_precision_1_sva_st_113[1] : mux_2010_nl;
  assign mux_2010_nl = cfg_proc_precision_1_sva_st_65[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_300_cse : cfg_out_precision_1_sva_st_113[1];
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_14_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_1_nl;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_1_nl = IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_1_FpMantRNE_17U_11U_else_acc_nl;
  assign mux_1268_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2237_cse : and_295_nl;
  assign mux_1267_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_94 : and_271_nl;
  assign IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt = mux_2000_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) { 5'b00000, FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0 } : IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2;
  assign mux_2000_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_out_precision_1_sva_st_149[1] : cfg_out_precision_1_sva_6[1];
  assign mux_1142_cse = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_455 : nor_1415_nl;
  assign mux_1126_cse = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4714_cse : nor_1434_nl;
  assign mux_1071_cse = or_1587_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_961 : nor_1463_nl;
  assign mux_1053_cse = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1051_nl : mux_1052_nl;
  assign mux_1052_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2186_cse : and_tmp_171;
  assign mux_1051_nl = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_1049 : mux_1050_nl;
  assign mux_1050_nl = cfg_proc_precision_1_sva_st_64[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00040_ : mux_tmp_1049;
  assign mux_1027_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1498_nl : nor_1500_cse;
  assign mux_1003_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1001_nl : mux_1002_nl;
  assign mux_1002_nl = or_1159_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1525_nl : nor_1524_nl;
  assign mux_1001_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1523_nl : nor_1556_cse;
  assign mux_991_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_985_nl : mux_990_nl;
  assign mux_990_nl = main_stage_v_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_988_nl : mux_989_cse;
  assign mux_988_nl = cfg_proc_precision_1_sva_st_108[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_987 : nor_1536_nl;
  assign mux_985_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1142_cse : mux_984_nl;
  assign mux_984_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_944 : _00073_;
  assign mux_989_cse = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1142_cse : and_1386_cse;
  assign mux_948_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_945 : mux_tmp_947;
  assign mux_938_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) main_stage_v_2 : main_stage_v_3;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_13_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_12_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_11_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_25_nl;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_25_nl = cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_9_FpMantRNE_17U_11U_else_acc_1_nl;
  assign mux_1933_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1930_nl : mux_1851_cse;
  assign mux_1930_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2149_nl : nor_2099_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_10_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_9_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0;
  assign mux_1916_nl = and_2151_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_2236_nl = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4714_cse : nor_2269_nl;
  assign mux_1909_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1864_cse : mux_1881_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_8_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_7_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0;
  assign mux_1892_nl = and_2153_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1889_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2142_nl : nor_2143_nl;
  assign mux_1888_nl = or_300_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_1886_nl = and_2154_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_2233_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2395_nl : or_4709_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_6_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0;
  assign mux_1882_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1849_cse : mux_1881_cse;
  assign mux_1881_cse = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1033_nl : mux_827_cse;
  assign mux_2232_nl = cfg_out_precision_1_sva_st_113[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4755_nl : and_2388_cse;
  assign mux_2231_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2388_cse : mux_2230_cse;
  assign mux_2230_cse = cfg_out_precision_1_sva_st_113[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_unequal_tmp_20 : or_4745_nl;
  assign mux_1867_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1864_cse : mux_1851_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_5_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0;
  assign mux_1864_cse = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1040_nl : nor_2099_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_4_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0;
  assign mux_1859_nl = and_2156_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_4862_cse : nor_50_cse;
  assign mux_2227_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_2371_nl : or_4709_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_3_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0;
  assign mux_1852_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1849_cse : mux_1851_cse;
  assign mux_1849_cse = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1048_cse : nor_2099_cse;
  assign mux_1851_cse = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1049_nl : mux_827_cse;
  assign mux_2226_nl = cfg_out_precision_1_sva_st_113[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2225_nl : or_4718_nl;
  assign mux_2225_nl = cfg_out_precision_1_sva_st_113[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_unequal_tmp_20 : nor_2284_nl;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_2_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0;
  assign mux_1831_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1828_nl : mux_1830_nl;
  assign mux_1830_nl = cvt_unequal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2101_nl : mux_827_cse;
  assign mux_1828_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2100_nl : nor_2099_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_1_nl = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_4_nl;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_4_nl = cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : cvt_2_FpMantRNE_17U_11U_else_acc_1_nl;
  assign mux_827_cse = or_1157_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1672_cse : or_1159_cse;
  assign mux_818_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_816_nl : mux_817_nl;
  assign mux_817_nl = or_1159_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1630_cse : nor_1661_nl;
  assign mux_816_nl = or_4862_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_1626_cse : nor_1659_nl;
  assign mux_813_cse = or_1159_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cfg_mode_eql_1_sva_6 : or_1176_cse;
  assign mux_800_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_11 : and_2237_cse;
  assign mux_796_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_1386_cse : and_tmp_94;
  assign mux_786_cse_1 = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_765 : nor_1674_nl;
  assign mux_767_cse = cfg_proc_precision_1_sva_st_89[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_766 : nor_1683_nl;
  assign mux_1817_nl = or_400_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1816_nl : or_3063_cse;
  assign mux_1816_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3696_cse : mux_1815_nl;
  assign mux_1815_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3220_nl : mux_1814_nl;
  assign mux_1814_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00072_ : or_3696_cse;
  assign mux_1808_nl = or_400_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1807_nl : or_3063_cse;
  assign mux_1807_nl = _07612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3696_cse : or_3196_nl;
  assign mux_660_cse = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1463_cse : nor_1761_nl;
  assign mux_1799_nl = or_400_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1798_nl : mux_1794_nl;
  assign mux_1798_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3032 : mux_1797_nl;
  assign mux_1797_nl = cfg_out_precision_1_sva_st_154[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nand_225_nl : mux_1796_nl;
  assign mux_1796_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3151_cse : not_tmp_270;
  assign mux_1794_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3032 : or_3170_nl;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_63_nl = fsm_output[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) 10'b0000000000 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0;
  assign mux_1791_nl = or_400_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_1790_nl : or_3063_cse;
  assign mux_1790_nl = _07612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3696_cse : nand_51_nl;
  assign mux_2196_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2195_nl : or_tmp_3379;
  assign mux_2195_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2193_nl : or_tmp_3379;
  assign mux_2193_nl = or_4559_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3379 : nor_2300_nl;
  assign mux_1788_nl = _07612_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3696_cse : or_3151_cse;
  assign mux_1780_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3063_cse : mux_1779_cse;
  assign mux_1779_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3696_cse : mux_2171_nl;
  assign mux_2171_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00071_ : or_3696_cse;
  assign mux_474_cse = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_317 : nor_1875_nl;
  assign mux_1762_cse = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3063_cse : mux_1761_cse;
  assign mux_417_cse = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_416 : nor_1917_nl;
  assign mux_382_cse = cfg_proc_precision_1_sva_st_65[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_345 : nor_1939_nl;
  assign mux_378_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_tmp_19 : and_178_itm;
  assign mux_2179_nl = or_4550_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2178_nl : or_tmp_3763;
  assign mux_2178_nl = or_183_cse_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_2177_nl : or_tmp_3763;
  assign mux_2177_nl = cfg_out_precision_1_sva_st_154[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_3763 : nor_2326_cse;
  assign mux_1761_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3696_cse : mux_1760_nl;
  assign mux_1760_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00070_ : or_3696_cse;
  assign mux_344_cse = cfg_proc_precision_1_sva_st_64[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_183_cse_1 : nor_1958_nl;
  assign mux_1758_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3070_nl : mux_1757_nl;
  assign mux_1757_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_tmp_2960 : mux_2170_nl;
  assign mux_2170_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00069_ : or_tmp_2960;
  assign mux_1752_nl = or_578_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3063_cse : mux_1751_nl;
  assign mux_1751_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_3696_cse : mux_1750_nl;
  assign mux_1750_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00068_ : or_3696_cse;
  assign mux_273_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) and_1386_cse : and_1078_cse;
  assign mux_201_cse = cfg_proc_precision_1_sva_st_101[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_200 : nor_2026_nl;
  assign mux_169_nl = or_309_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_303_cse : mux_166_cse;
  assign mux_166_cse = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) or_306_cse : or_tmp_306;
  assign mux_163_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) nor_2047_cse : nor_2046_nl;
  assign mux_12_nl = or_5189_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_in_rsci_bawt : main_stage_v_1;
  assign mux_2355_nl = cfg_proc_precision_1_sva_st_90[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) mux_tmp_2347 : mux_2354_nl;
  assign mux_2354_nl = cfg_proc_precision_1_sva_st_90[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) _00055_ : mux_tmp_2347;
  assign _00987_ = _02624_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21412" *) cvt_16_FpMantRNE_24U_11U_else_and_4_tmp : cvt_16_FpMantRNE_24U_11U_else_and_4_svs;
  assign _00974_ = _02623_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21402" *) cvt_15_FpMantRNE_24U_11U_else_and_3_tmp : cvt_15_FpMantRNE_24U_11U_else_and_3_svs;
  assign _00960_ = _02622_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21392" *) cvt_14_FpMantRNE_24U_11U_else_and_3_tmp : cvt_14_FpMantRNE_24U_11U_else_and_3_svs;
  assign _00947_ = _02621_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21382" *) cvt_13_FpMantRNE_24U_11U_else_and_2_tmp : cvt_13_FpMantRNE_24U_11U_else_and_2_svs;
  assign _00934_ = _02620_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21372" *) cvt_12_FpMantRNE_24U_11U_else_and_3_tmp : cvt_12_FpMantRNE_24U_11U_else_and_3_svs;
  assign _00921_ = _02619_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21362" *) cvt_11_FpMantRNE_24U_11U_else_and_2_tmp : cvt_11_FpMantRNE_24U_11U_else_and_2_svs;
  assign _00908_ = _02618_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21352" *) cvt_10_FpMantRNE_24U_11U_else_and_2_tmp : cvt_10_FpMantRNE_24U_11U_else_and_2_svs;
  assign _01115_ = _02617_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21342" *) cvt_9_FpMantRNE_24U_11U_else_and_1_tmp : cvt_9_FpMantRNE_24U_11U_else_and_1_svs;
  assign _01101_ = _02616_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21332" *) cvt_8_FpMantRNE_24U_11U_else_and_3_tmp : cvt_8_FpMantRNE_24U_11U_else_and_3_svs;
  assign _01087_ = _02615_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21322" *) cvt_7_FpMantRNE_24U_11U_else_and_2_tmp : cvt_7_FpMantRNE_24U_11U_else_and_2_svs;
  assign _01073_ = _02614_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21312" *) cvt_6_FpMantRNE_24U_11U_else_and_2_tmp : cvt_6_FpMantRNE_24U_11U_else_and_2_svs;
  assign _01058_ = _02613_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21302" *) cvt_5_FpMantRNE_24U_11U_else_and_1_tmp : cvt_5_FpMantRNE_24U_11U_else_and_1_svs;
  assign _01043_ = _02612_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21292" *) cvt_4_FpMantRNE_24U_11U_else_and_2_tmp : cvt_4_FpMantRNE_24U_11U_else_and_2_svs;
  assign _01028_ = _02611_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21282" *) cvt_3_FpMantRNE_24U_11U_else_and_1_tmp : cvt_3_FpMantRNE_24U_11U_else_and_1_svs;
  assign _01014_ = _02610_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21272" *) cvt_2_FpMantRNE_24U_11U_else_and_1_tmp : cvt_2_FpMantRNE_24U_11U_else_and_1_svs;
  assign _00999_ = _02609_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21262" *) cvt_1_FpMantRNE_24U_11U_else_and_tmp : cvt_1_FpMantRNE_24U_11U_else_and_svs;
  assign _00983_ = _02608_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21252" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp : cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs;
  assign _00970_ = _02607_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21243" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  assign _00956_ = _02606_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21234" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  assign _00930_ = _02604_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21226" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  assign _00917_ = FpIntToFloat_17U_5U_10U_if_and_36_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21216" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  assign _00904_ = FpIntToFloat_17U_5U_10U_if_and_36_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21216" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  assign _01097_ = _02603_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21207" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  assign _01083_ = FpIntToFloat_17U_5U_10U_if_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21197" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  assign _01069_ = FpIntToFloat_17U_5U_10U_if_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21197" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  assign _00625_ = _02601_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21188" *) IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_5_sva;
  assign _01053_ = _02599_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21180" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs;
  assign _00943_ = FpIntToFloat_17U_5U_10U_if_and_31_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21170" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  assign _01039_ = FpIntToFloat_17U_5U_10U_if_and_31_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21170" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  assign _00617_ = _02597_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21161" *) IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_1_sva;
  assign _01384_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0;
  assign _00311_ = _02595_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21152" *) _01384_ : FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign _01383_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0;
  assign _01382_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0;
  assign _01381_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0;
  assign _01380_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0;
  assign _01379_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp : FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0;
  assign _00307_ = FpIntToFloat_17U_5U_10U_is_inf_and_28_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21134" *) _01383_ : FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign _00305_ = FpIntToFloat_17U_5U_10U_is_inf_and_28_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21134" *) _01382_ : FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign _00325_ = FpIntToFloat_17U_5U_10U_is_inf_and_28_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21134" *) _01381_ : FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign _00323_ = FpIntToFloat_17U_5U_10U_is_inf_and_28_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21134" *) _01380_ : FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign _00320_ = FpIntToFloat_17U_5U_10U_is_inf_and_28_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21134" *) _01379_ : FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign _00295_ = _02594_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21122" *) or_5086_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_15;
  assign _00986_ = _02592_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21112" *) cvt_16_FpMantRNE_17U_11U_else_and_4_tmp : cvt_16_FpMantRNE_17U_11U_else_and_4_svs;
  assign _00294_ = _02591_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21103" *) or_5069_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_14;
  assign _00973_ = _02589_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21094" *) cvt_15_FpMantRNE_17U_11U_else_and_3_tmp : cvt_15_FpMantRNE_17U_11U_else_and_3_svs;
  assign _00293_ = _02588_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21084" *) or_5053_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_13;
  assign _00959_ = _02586_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21075" *) cvt_14_FpMantRNE_17U_11U_else_and_3_tmp : cvt_14_FpMantRNE_17U_11U_else_and_3_svs;
  assign _00292_ = _02585_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21065" *) or_5038_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_12;
  assign _00946_ = _02583_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21055" *) cvt_13_FpMantRNE_17U_11U_else_and_2_tmp : cvt_13_FpMantRNE_17U_11U_else_and_2_svs;
  assign _00291_ = _02582_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21045" *) or_1925_cse_1 : FpIntToFloat_17U_5U_10U_else_unequal_tmp_11;
  assign _00933_ = _02580_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21035" *) cvt_12_FpMantRNE_17U_11U_else_and_3_tmp : cvt_12_FpMantRNE_17U_11U_else_and_3_svs;
  assign _00290_ = _02579_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21024" *) or_1892_cse_1 : FpIntToFloat_17U_5U_10U_else_unequal_tmp_10;
  assign _00920_ = _02577_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21016" *) cvt_11_FpMantRNE_17U_11U_else_and_2_tmp : cvt_11_FpMantRNE_17U_11U_else_and_2_svs;
  assign _00304_ = _02576_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:21007" *) or_1851_cse_1 : FpIntToFloat_17U_5U_10U_else_unequal_tmp_9;
  assign _00907_ = _02574_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20998" *) cvt_10_FpMantRNE_17U_11U_else_and_2_tmp : cvt_10_FpMantRNE_17U_11U_else_and_2_svs;
  assign _00303_ = _02573_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20989" *) or_1829_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_8;
  assign _01114_ = _02571_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20979" *) cvt_9_FpMantRNE_17U_11U_else_and_1_tmp : cvt_9_FpMantRNE_17U_11U_else_and_1_svs;
  assign _00302_ = _02570_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20969" *) or_1789_cse_1 : FpIntToFloat_17U_5U_10U_else_unequal_tmp_7;
  assign _01100_ = _02568_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20960" *) cvt_8_FpMantRNE_17U_11U_else_and_3_tmp : cvt_8_FpMantRNE_17U_11U_else_and_3_svs;
  assign _00301_ = _02567_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20949" *) or_1752_cse_1 : FpIntToFloat_17U_5U_10U_else_unequal_tmp_6;
  assign _01086_ = _02565_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20941" *) cvt_7_FpMantRNE_17U_11U_else_and_2_tmp : cvt_7_FpMantRNE_17U_11U_else_and_2_svs;
  assign _00300_ = _02564_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20931" *) or_1720_cse_1 : FpIntToFloat_17U_5U_10U_else_unequal_tmp_5;
  assign _01072_ = _02562_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20923" *) cvt_6_FpMantRNE_17U_11U_else_and_2_tmp : cvt_6_FpMantRNE_17U_11U_else_and_2_svs;
  assign _00299_ = _02561_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20914" *) or_1693_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_4;
  assign _01057_ = _02559_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20904" *) cvt_5_FpMantRNE_17U_11U_else_and_1_tmp : cvt_5_FpMantRNE_17U_11U_else_and_1_svs;
  assign _00298_ = _02558_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20893" *) or_1659_cse_1 : FpIntToFloat_17U_5U_10U_else_unequal_tmp_3;
  assign _01042_ = _02556_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20885" *) cvt_4_FpMantRNE_17U_11U_else_and_2_tmp : cvt_4_FpMantRNE_17U_11U_else_and_2_svs;
  assign _00297_ = _02555_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20876" *) or_1625_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_2;
  assign _01027_ = _02553_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20867" *) cvt_3_FpMantRNE_17U_11U_else_and_1_tmp : cvt_3_FpMantRNE_17U_11U_else_and_1_svs;
  assign _00296_ = _02552_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20858" *) or_1596_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp_1;
  assign _01013_ = _02550_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20849" *) cvt_2_FpMantRNE_17U_11U_else_and_1_tmp : cvt_2_FpMantRNE_17U_11U_else_and_1_svs;
  assign _00289_ = _02549_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20840" *) or_1202_cse : FpIntToFloat_17U_5U_10U_else_unequal_tmp;
  assign _00998_ = _02547_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20831" *) cvt_1_FpMantRNE_17U_11U_else_and_tmp : cvt_1_FpMantRNE_17U_11U_else_and_svs;
  assign _01378_ = and_1467_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0;
  assign _00566_ = _02546_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20820" *) _01378_ : IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm;
  assign _01377_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0;
  assign _00559_ = _02542_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20809" *) _01377_ : IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm;
  assign _01376_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0;
  assign _00565_ = _02541_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20798" *) _01376_ : IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm;
  assign _01375_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp : IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0;
  assign _00574_ = _02540_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20787" *) _01375_ : IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm;
  assign _01374_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0;
  assign _01373_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0;
  assign _00564_ = IntShiftRightSat_49U_6U_17U_oelse_and_25_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20773" *) _01373_ : IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm;
  assign _00563_ = IntShiftRightSat_49U_6U_17U_oelse_and_25_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20773" *) _01374_ : IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm;
  assign _01372_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0;
  assign _00562_ = _02538_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20762" *) _01372_ : IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm;
  assign _01371_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0;
  assign _01370_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0;
  assign _00561_ = IntShiftRightSat_49U_6U_17U_oelse_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20748" *) _01371_ : IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm;
  assign _00560_ = IntShiftRightSat_49U_6U_17U_oelse_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20748" *) _01370_ : IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm;
  assign _01369_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp : IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0;
  assign _00570_ = _02537_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20737" *) _01369_ : IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm;
  assign _01368_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0;
  assign _00573_ = _02536_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20726" *) _01368_ : IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm;
  assign _01367_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0;
  assign _01366_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0;
  assign _00572_ = IntShiftRightSat_49U_6U_17U_oelse_and_18_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20712" *) _01367_ : IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm;
  assign _00571_ = IntShiftRightSat_49U_6U_17U_oelse_and_18_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20712" *) _01366_ : IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm;
  assign _01365_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0;
  assign _00569_ = _02534_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20701" *) _01365_ : IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm;
  assign _01364_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp : IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0;
  assign _01363_ = and_1385_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp : IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0;
  assign _00568_ = IntShiftRightSat_49U_6U_17U_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20687" *) _01364_ : IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm;
  assign _00567_ = IntShiftRightSat_49U_6U_17U_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20687" *) _01363_ : IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm;
  assign _01362_ = and_dcpl_204 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : IsNaN_5U_10U_IsNaN_5U_10U_nand_14_nl;
  assign _00681_ = _02533_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20676" *) _01362_ : IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2;
  assign _01361_ = and_dcpl_204 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : IsNaN_5U_10U_nor_14_nl;
  assign _00713_ = _02532_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20666" *) _01361_ : IsNaN_5U_10U_nor_14_itm_2;
  assign _01360_ = and_dcpl_204 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp : IsNaN_5U_10U_IsNaN_5U_10U_nand_1_nl;
  assign _00682_ = _02531_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20656" *) _01360_ : IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  assign _01359_ = and_dcpl_204 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : IsNaN_5U_10U_nor_1_nl;
  assign _00714_ = _02530_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20646" *) _01359_ : IsNaN_5U_10U_nor_1_itm_2;
  assign _01358_ = and_dcpl_204 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : IsNaN_5U_10U_IsNaN_5U_10U_nand_nl;
  assign _00683_ = _02529_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20635" *) _01358_ : IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2;
  assign _01357_ = and_dcpl_204 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp : IsNaN_5U_10U_nor_nl;
  assign _00715_ = _02528_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20625" *) _01357_ : IsNaN_5U_10U_nor_itm_2;
  assign _00771_ = _02527_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20616" *) chn_idata_data_sva_1_27_0_1[15:0] : chn_idata_data_sva_2_15_0_1;
  assign _00526_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07866_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2;
  assign _00516_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07877_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2;
  assign _00518_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07865_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2;
  assign _00519_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07876_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2;
  assign _00520_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07864_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2;
  assign _00521_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07875_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2;
  assign _00522_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07874_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2;
  assign _00523_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07873_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2;
  assign _00524_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07863_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2;
  assign _00525_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07872_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2;
  assign _00508_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07871_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2;
  assign _00509_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07870_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2;
  assign _00510_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07869_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2;
  assign _00514_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07868_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2;
  assign _00515_ = IntSaturation_17U_16U_and_33_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20579" *) _07867_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2;
  assign _00533_ = _02511_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20555" *) _09166_ : IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5;
  assign _00534_ = _02509_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20543" *) _09165_ : IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6;
  assign _00535_ = _02507_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20531" *) _09164_ : IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6;
  assign _00536_ = _02505_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20519" *) _09163_ : IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7;
  assign _00537_ = _02503_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20507" *) _09162_ : IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6;
  assign _00538_ = _02501_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20495" *) _09161_ : IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7;
  assign _00539_ = _02499_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20483" *) _09160_ : IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7;
  assign _00540_ = _02497_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20471" *) _09159_ : IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8;
  assign _00541_ = _02495_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20459" *) _09158_ : IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6;
  assign _00527_ = _02493_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20447" *) _09157_ : IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7;
  assign _00528_ = _02491_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20435" *) _09156_ : IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7;
  assign _00529_ = _02489_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20423" *) _09155_ : IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8;
  assign _00530_ = _02487_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20411" *) _09154_ : IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7;
  assign _00531_ = _02485_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20399" *) _09153_ : IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8;
  assign _00532_ = _02483_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20387" *) _09152_ : IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8;
  assign _00542_ = _02481_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20375" *) _09151_ : IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9;
  assign _01356_ = and_1381_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_1_FpMantRNE_24U_11U_else_and_svs : cvt_1_FpMantRNE_24U_11U_else_and_tmp;
  assign _01000_ = _02479_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20364" *) _01356_ : cvt_1_FpMantRNE_24U_11U_else_and_svs_2;
  assign _00448_ = _02474_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20354" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9;
  assign _01355_ = and_1377_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_2_FpMantRNE_24U_11U_else_and_1_svs : cvt_2_FpMantRNE_24U_11U_else_and_1_tmp;
  assign _01015_ = _02473_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20345" *) _01355_ : cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign _00451_ = _02468_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20335" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9;
  assign _01354_ = and_1373_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_3_FpMantRNE_24U_11U_else_and_1_svs : cvt_3_FpMantRNE_24U_11U_else_and_1_tmp;
  assign _01029_ = _02467_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20326" *) _01354_ : cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign _00454_ = _02462_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20316" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9;
  assign _01353_ = and_1369_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpMantRNE_24U_11U_else_and_2_svs : cvt_4_FpMantRNE_24U_11U_else_and_2_tmp;
  assign _01044_ = _02461_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20307" *) _01353_ : cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign _00457_ = _02456_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20297" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9;
  assign _01352_ = and_1365_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_FpMantRNE_24U_11U_else_and_1_svs : cvt_5_FpMantRNE_24U_11U_else_and_1_tmp;
  assign _01059_ = _02455_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20288" *) _01352_ : cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign _00460_ = _02450_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20278" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9;
  assign _01351_ = and_1361_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpMantRNE_24U_11U_else_and_2_svs : cvt_6_FpMantRNE_24U_11U_else_and_2_tmp;
  assign _01074_ = _02449_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20269" *) _01351_ : cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign _00463_ = _02444_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20259" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9;
  assign _01350_ = and_1357_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpMantRNE_24U_11U_else_and_2_svs : cvt_7_FpMantRNE_24U_11U_else_and_2_tmp;
  assign _01088_ = _02443_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20250" *) _01350_ : cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign _00466_ = _02438_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20240" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9;
  assign _01349_ = and_1353_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpMantRNE_24U_11U_else_and_3_svs : cvt_8_FpMantRNE_24U_11U_else_and_3_tmp;
  assign _01102_ = _02437_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20231" *) _01349_ : cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign _00469_ = _02432_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20221" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9;
  assign _01348_ = and_1349_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_9_FpMantRNE_24U_11U_else_and_1_svs : cvt_9_FpMantRNE_24U_11U_else_and_1_tmp;
  assign _01116_ = _02431_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20212" *) _01348_ : cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2;
  assign _00472_ = _02426_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20202" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9;
  assign _01347_ = and_1345_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpMantRNE_24U_11U_else_and_2_svs : cvt_10_FpMantRNE_24U_11U_else_and_2_tmp;
  assign _00909_ = _02425_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20193" *) _01347_ : cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign _00430_ = _02420_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20183" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9;
  assign _01346_ = and_1341_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpMantRNE_24U_11U_else_and_2_svs : cvt_11_FpMantRNE_24U_11U_else_and_2_tmp;
  assign _00922_ = _02419_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20174" *) _01346_ : cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign _00433_ = _02414_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20164" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9;
  assign _01345_ = and_1337_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpMantRNE_24U_11U_else_and_3_svs : cvt_12_FpMantRNE_24U_11U_else_and_3_tmp;
  assign _00935_ = _02413_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20155" *) _01345_ : cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign _00436_ = _02408_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20145" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9;
  assign _01344_ = and_1333_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpMantRNE_24U_11U_else_and_2_svs : cvt_13_FpMantRNE_24U_11U_else_and_2_tmp;
  assign _00948_ = _02407_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20136" *) _01344_ : cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2;
  assign _00439_ = _02402_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20126" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9;
  assign _01343_ = and_1329_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpMantRNE_24U_11U_else_and_3_svs : cvt_14_FpMantRNE_24U_11U_else_and_3_tmp;
  assign _00961_ = _02401_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20117" *) _01343_ : cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign _00442_ = _02396_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20107" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9;
  assign _01342_ = and_1325_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpMantRNE_24U_11U_else_and_3_svs : cvt_15_FpMantRNE_24U_11U_else_and_3_tmp;
  assign _00975_ = _02395_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20098" *) _01342_ : cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2;
  assign _00445_ = _02390_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20088" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9;
  assign _01341_ = and_1321_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpMantRNE_24U_11U_else_and_4_svs : cvt_16_FpMantRNE_24U_11U_else_and_4_tmp;
  assign _00988_ = _02389_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20079" *) _01341_ : cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2;
  assign _00475_ = _02384_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20069" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9;
  assign _00363_ = _02383_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20061" *) FpMantRNE_24U_11U_else_carry_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_sva_2;
  assign _00347_ = _02382_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20053" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2;
  assign _00353_ = _02381_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20045" *) FpMantRNE_24U_11U_else_carry_15_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_15_sva_2;
  assign _00337_ = _02380_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20037" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2;
  assign _00352_ = _02379_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20029" *) FpMantRNE_24U_11U_else_carry_14_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_14_sva_2;
  assign _00336_ = _02378_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20021" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2;
  assign _00351_ = _02377_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20013" *) FpMantRNE_24U_11U_else_carry_13_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_13_sva_2;
  assign _00335_ = _02376_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:20005" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2;
  assign _00350_ = _02375_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19997" *) FpMantRNE_24U_11U_else_carry_12_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_12_sva_2;
  assign _00334_ = _02374_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19989" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2;
  assign _00349_ = _02373_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19981" *) FpMantRNE_24U_11U_else_carry_11_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_11_sva_2;
  assign _00333_ = _02372_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19973" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2;
  assign _00348_ = _02371_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19965" *) FpMantRNE_24U_11U_else_carry_10_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_10_sva_2;
  assign _00332_ = _02370_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19957" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2;
  assign _00362_ = _02369_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19949" *) FpMantRNE_24U_11U_else_carry_9_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_9_sva_2;
  assign _00346_ = _02368_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19941" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2[4:0] : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2;
  assign _00361_ = _02367_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19933" *) FpMantRNE_24U_11U_else_carry_8_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_8_sva_2;
  assign _00345_ = _02366_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19925" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2[4:0] : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2;
  assign _00360_ = _02365_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19917" *) FpMantRNE_24U_11U_else_carry_7_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_7_sva_2;
  assign _00344_ = _02364_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19909" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2;
  assign _00359_ = _02363_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19901" *) FpMantRNE_24U_11U_else_carry_6_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_6_sva_2;
  assign _00343_ = _02362_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19893" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2;
  assign _00358_ = _02361_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19885" *) FpMantRNE_24U_11U_else_carry_5_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_5_sva_2;
  assign _00342_ = _02360_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19877" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2;
  assign _00357_ = _02359_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19869" *) FpMantRNE_24U_11U_else_carry_4_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_4_sva_2;
  assign _00341_ = _02358_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19861" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2;
  assign _00356_ = _02357_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19853" *) FpMantRNE_24U_11U_else_carry_3_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_3_sva_2;
  assign _00340_ = _02356_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19845" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2;
  assign _00355_ = _02355_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19837" *) FpMantRNE_24U_11U_else_carry_2_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_2_sva_2;
  assign _00339_ = _02354_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19829" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2;
  assign _00354_ = _02353_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19821" *) FpMantRNE_24U_11U_else_carry_1_sva_mx0w0 : FpMantRNE_24U_11U_else_carry_1_sva_2;
  assign _00338_ = _02352_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19813" *) nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 : FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2;
  assign _00766_ = _02351_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19805" *) chn_in_rsci_d_mxwt[511] : chn_idata_data_sva_1_511_1;
  assign _00678_ = IntShiftRightSat_49U_6U_17U_o_and_115_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19796" *) IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_sva;
  assign _00635_ = IntShiftRightSat_49U_6U_17U_o_and_115_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19796" *) IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_sva;
  assign _00652_ = IntShiftRightSat_49U_6U_17U_o_and_114_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19786" *) IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_15_sva;
  assign _00615_ = IntShiftRightSat_49U_6U_17U_o_and_114_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19786" *) IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_15_sva;
  assign _00511_ = IntShiftRightSat_49U_6U_17U_o_and_112_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19771" *) IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0 : IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm;
  assign _00649_ = IntShiftRightSat_49U_6U_17U_o_and_112_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19771" *) IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_14_sva;
  assign _00613_ = IntShiftRightSat_49U_6U_17U_o_and_112_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19771" *) IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_14_sva;
  assign _00646_ = IntShiftRightSat_49U_6U_17U_o_and_112_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19771" *) IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_13_sva;
  assign _00611_ = IntShiftRightSat_49U_6U_17U_o_and_112_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19771" *) IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_13_sva;
  assign _00662_ = IntShiftRightSat_49U_6U_17U_o_and_112_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19771" *) IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_4_sva;
  assign _00623_ = IntShiftRightSat_49U_6U_17U_o_and_112_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19771" *) IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_4_sva;
  assign _00643_ = IntShiftRightSat_49U_6U_17U_o_and_111_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19756" *) IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_12_sva;
  assign _00609_ = IntShiftRightSat_49U_6U_17U_o_and_111_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19756" *) IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_12_sva;
  assign _00640_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_11_sva;
  assign _00607_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_11_sva;
  assign _00637_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_10_sva;
  assign _00605_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_10_sva;
  assign _00633_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_9_sva;
  assign _00621_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_3_sva;
  assign _00657_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_2_sva;
  assign _00619_ = IntShiftRightSat_49U_6U_17U_o_and_109_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19740" *) IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_2_sva;
  assign _00673_ = IntShiftRightSat_49U_6U_17U_o_and_108_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19724" *) IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_8_sva;
  assign _00631_ = IntShiftRightSat_49U_6U_17U_o_and_108_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19724" *) IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_8_sva;
  assign _00670_ = IntShiftRightSat_49U_6U_17U_o_and_107_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19712" *) IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_7_sva;
  assign _00629_ = IntShiftRightSat_49U_6U_17U_o_and_107_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19712" *) IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_7_sva;
  assign _00667_ = IntShiftRightSat_49U_6U_17U_o_and_107_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19712" *) IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_6_sva;
  assign _00627_ = IntShiftRightSat_49U_6U_17U_o_and_107_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19712" *) IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_15_1_6_sva;
  assign _01340_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs : cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign _00957_ = FpIntToFloat_17U_5U_10U_if_and_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19700" *) _01340_ : cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _01339_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs : cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp;
  assign _01338_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs : cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign _01337_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs : cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign _00984_ = FpIntToFloat_17U_5U_10U_if_and_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19686" *) _01339_ : cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2;
  assign _00971_ = FpIntToFloat_17U_5U_10U_if_and_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19686" *) _01338_ : cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _00944_ = FpIntToFloat_17U_5U_10U_if_and_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19686" *) _01337_ : cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _01336_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs : cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign _01335_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs : cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  assign _00931_ = FpIntToFloat_17U_5U_10U_if_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19673" *) _01336_ : cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _01098_ = FpIntToFloat_17U_5U_10U_if_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19673" *) _01335_ : cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign _01334_ = and_1250_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs : cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  assign _01054_ = _02348_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19663" *) _01334_ : cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _01333_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs : cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign _01332_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs : cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign _01331_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs : cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign _01330_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs : cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign _01329_ = and_1247_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs : cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  assign _00918_ = FpIntToFloat_17U_5U_10U_if_and_18_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19646" *) _01333_ : cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _00905_ = FpIntToFloat_17U_5U_10U_if_and_18_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19646" *) _01332_ : cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _01084_ = FpIntToFloat_17U_5U_10U_if_and_18_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19646" *) _01331_ : cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _01070_ = FpIntToFloat_17U_5U_10U_if_and_18_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19646" *) _01330_ : cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _01040_ = FpIntToFloat_17U_5U_10U_if_and_18_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19646" *) _01329_ : cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign _01111_ = FpIntToFloat_17U_5U_10U_if_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19632" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _01024_ = FpIntToFloat_17U_5U_10U_if_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19632" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _01010_ = FpIntToFloat_17U_5U_10U_if_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19632" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign _01328_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp : FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0;
  assign _01327_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0;
  assign _00330_ = FpIntToFloat_17U_5U_10U_is_inf_and_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19619" *) _01328_ : FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign _00315_ = FpIntToFloat_17U_5U_10U_is_inf_and_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19619" *) _01327_ : FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign _01326_ = and_1213_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0;
  assign _00313_ = _02346_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19609" *) _01326_ : FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign _01325_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0;
  assign _01324_ = and_1249_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp : FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0;
  assign _00309_ = FpIntToFloat_17U_5U_10U_is_inf_and_23_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19596" *) _01325_ : FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign _00327_ = FpIntToFloat_17U_5U_10U_is_inf_and_23_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19596" *) _01324_ : FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign _01229_ = _02338_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19587" *) chn_idata_data_mux1h_65_rgt[9:0] : reg_chn_idata_data_sva_3_15_0_2_reg;
  assign _01228_ = _02336_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19578" *) chn_idata_data_mux1h_65_rgt[14:10] : reg_chn_idata_data_sva_3_15_0_1_reg;
  assign _01230_ = _02334_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19568" *) chn_idata_data_mux1h_65_rgt[15] : reg_chn_idata_data_sva_3_15_0_reg;
  assign _00750_ = cfg_proc_precision_and_43_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19559" *) cfg_proc_precision_1_sva_st_89 : cfg_proc_precision_1_sva_st_90;
  assign _00738_ = cfg_proc_precision_and_43_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19559" *) cfg_out_precision_1_sva_st_113 : cfg_out_precision_1_sva_st_136;
  assign _00744_ = cfg_proc_precision_and_40_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19549" *) cfg_proc_precision_1_sva_st_101 : cfg_proc_precision_1_sva_st_102;
  assign _00739_ = cfg_proc_precision_and_40_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19549" *) cfg_out_precision_1_sva_st_149 : cfg_out_precision_1_sva_st_144;
  assign _00745_ = _02333_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19540" *) cfg_proc_precision_1_sva_st_101 : cfg_proc_precision_1_sva_st_108;
  assign _00742_ = _02332_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19532" *) cfg_out_precision_1_sva_st_149 : cfg_out_precision_1_sva_st_156;
  assign _01223_ = _02331_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19524" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm;
  assign _01224_ = _02327_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19515" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm;
  assign _01203_ = _02315_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19503" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm;
  assign _01204_ = _02312_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19494" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm;
  assign _01323_ = and_dcpl_648 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0;
  assign _01322_ = and_dcpl_648 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0;
  assign _00331_ = FpIntToFloat_17U_5U_10U_is_inf_and_10_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19479" *) _01323_ : FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  assign _00316_ = FpIntToFloat_17U_5U_10U_is_inf_and_10_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19479" *) _01322_ : FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  assign _01226_ = _02299_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19470" *) IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt[9:0] : reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg;
  assign _01225_ = _02300_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19461" *) IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt[14:10] : reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg;
  assign _01201_ = _02298_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19453" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm;
  assign _01202_ = _02295_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19444" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm;
  assign _00513_ = _02283_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19432" *) IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3 : IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4;
  assign _00583_ = _02282_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19424" *) IntShiftRightSat_49U_6U_17U_o_0_14_sva_3 : IntShiftRightSat_49U_6U_17U_o_0_14_sva_4;
  assign _01199_ = _02281_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19416" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm;
  assign _01200_ = _02277_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19407" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm;
  assign _01321_ = and_dcpl_631 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0;
  assign _01320_ = and_dcpl_631 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0;
  assign _00314_ = FpIntToFloat_17U_5U_10U_is_inf_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19392" *) _01321_ : FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  assign _00312_ = FpIntToFloat_17U_5U_10U_is_inf_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19392" *) _01320_ : FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7;
  assign _01197_ = _02265_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19383" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm;
  assign _01198_ = _02261_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19374" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm;
  assign _01319_ = and_dcpl_617 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0;
  assign _00310_ = _02249_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19361" *) _01319_ : FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  assign _01195_ = _02248_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19352" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm;
  assign _01196_ = _02244_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19343" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm;
  assign _01318_ = and_dcpl_617 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0;
  assign _00308_ = _02232_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19330" *) _01318_ : FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  assign _01193_ = _02230_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19321" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm;
  assign _01194_ = _02226_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19312" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm;
  assign _01317_ = and_dcpl_617 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0;
  assign _00306_ = _02214_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19299" *) _01317_ : FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7;
  assign _01120_ = _02213_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19290" *) cvt_9_IntSaturation_17U_8U_if_acc_1_nl[10] : cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  assign _01221_ = _02212_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19281" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm;
  assign _01222_ = _02208_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19272" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm;
  assign _00329_ = _02195_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19258" *) _04930_ : FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7;
  assign _01219_ = _02194_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19250" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm;
  assign _01220_ = _02190_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19241" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm;
  assign _01316_ = and_1104_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0;
  assign _00328_ = _02178_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19228" *) _01316_ : FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  assign _01217_ = _02177_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19219" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm;
  assign _01218_ = _02173_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19210" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm;
  assign _01315_ = and_1104_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0;
  assign _00326_ = _02161_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19197" *) _01315_ : FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  assign _01215_ = _02160_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19188" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm;
  assign _01216_ = _02156_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19179" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm;
  assign _01314_ = and_1104_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0;
  assign _00324_ = _02144_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19166" *) _01314_ : FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  assign _01063_ = _02142_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19156" *) cvt_5_IntSaturation_17U_8U_if_acc_1_nl[10] : cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  assign _01213_ = _02141_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19147" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm;
  assign _01214_ = _02137_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19138" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm;
  assign _01211_ = _02126_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19126" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm;
  assign _01212_ = _02123_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19117" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm;
  assign _01313_ = and_1091_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp_1 : FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0;
  assign _00321_ = _02111_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19104" *) _01313_ : FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7;
  assign _01033_ = _02108_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19094" *) cvt_3_IntSaturation_17U_8U_if_acc_1_nl[10] : cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  assign _01209_ = _02107_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19085" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm;
  assign _01210_ = _02103_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19076" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm;
  assign _00322_ = FpIntToFloat_17U_5U_10U_is_inf_and_14_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19059" *) _04912_ : FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7;
  assign _00319_ = FpIntToFloat_17U_5U_10U_is_inf_and_14_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19059" *) _04909_ : FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7;
  assign _01207_ = _02088_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19050" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm;
  assign _01208_ = _02084_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19041" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm;
  assign _01312_ = and_1077_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_else_equal_tmp : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_nor_1_nl;
  assign _00318_ = _02073_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19028" *) _01312_ : FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  assign _01004_ = _02070_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19018" *) cvt_1_IntSaturation_17U_8U_if_acc_nl[10] : cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2;
  assign _01205_ = _02069_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19009" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm[3:0] : reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm;
  assign _01206_ = _02065_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:19000" *) FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm[4] : reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm;
  assign _00317_ = _02054_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18987" *) _04900_ : FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6;
  assign _00590_ = IntShiftRightSat_49U_6U_17U_o_and_103_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18977" *) IntShiftRightSat_49U_6U_17U_o_0_3_sva_3 : IntShiftRightSat_49U_6U_17U_o_0_3_sva_4;
  assign _00594_ = IntShiftRightSat_49U_6U_17U_o_and_103_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18977" *) IntShiftRightSat_49U_6U_17U_o_0_5_sva_3 : IntShiftRightSat_49U_6U_17U_o_0_5_sva_4;
  assign _00602_ = IntShiftRightSat_49U_6U_17U_o_and_103_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18977" *) IntShiftRightSat_49U_6U_17U_o_0_9_sva_3 : IntShiftRightSat_49U_6U_17U_o_0_9_sva_4;
  assign _00677_ = _02053_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18967" *) IntShiftRightSat_49U_6U_17U_o_16_9_sva_3 : IntShiftRightSat_49U_6U_17U_o_16_9_sva_4;
  assign _00803_ = _02052_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18959" *) chn_odata_data_13_0_lpi_1_dfm_1_mx0w0 : chn_odata_data_13_0_lpi_1_dfm_1;
  assign _01133_ = cvt_else_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18949" *) cvt_else_nor_dfs : cvt_else_nor_dfs_15;
  assign _01128_ = cvt_else_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18949" *) cvt_else_equal_tmp_1 : cvt_else_equal_tmp_46;
  assign _01127_ = cvt_else_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18949" *) cvt_else_equal_tmp : cvt_else_equal_tmp_45;
  assign _01131_ = _02051_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18939" *) cvt_else_nor_dfs : cvt_else_nor_dfs_10;
  assign _01132_ = cvt_else_and_34_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18928" *) cvt_else_nor_dfs : cvt_else_nor_dfs_11;
  assign _01126_ = cvt_else_and_34_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18928" *) cvt_else_equal_tmp_1 : cvt_else_equal_tmp_34;
  assign _01125_ = cvt_else_and_34_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18928" *) cvt_else_equal_tmp : cvt_else_equal_tmp_33;
  assign _01232_ = cvt_else_and_10_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18917" *) cvt_else_nor_dfs : reg_cvt_else_nor_dfs_9_cse;
  assign _01124_ = cvt_else_and_10_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18917" *) cvt_else_equal_tmp_1 : cvt_else_equal_tmp_28;
  assign _00666_ = _02049_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18908" *) IntShiftRightSat_49U_6U_17U_o_16_5_sva_3 : IntShiftRightSat_49U_6U_17U_o_16_5_sva_4;
  assign _01123_ = _02048_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18900" *) cvt_else_equal_tmp_1 : cvt_else_equal_tmp_16;
  assign _00661_ = _02046_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18891" *) IntShiftRightSat_49U_6U_17U_o_16_3_sva_3 : IntShiftRightSat_49U_6U_17U_o_16_3_sva_4;
  assign _01130_ = _02045_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18883" *) cvt_else_equal_tmp : cvt_else_equal_tmp_9;
  assign _01134_ = cvt_else_and_24_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18873" *) cvt_else_nor_dfs : cvt_else_nor_dfs_2;
  assign _01129_ = cvt_else_and_24_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18873" *) cvt_else_equal_tmp_1 : cvt_else_equal_tmp_5;
  assign _00680_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_sva_3;
  assign _00654_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_15_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_15_sva_3;
  assign _00651_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_14_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_14_sva_3;
  assign _00648_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_13_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_13_sva_3;
  assign _00645_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_12_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_12_sva_3;
  assign _00642_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_11_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_11_sva_3;
  assign _00639_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_10_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_10_sva_3;
  assign _00675_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_8_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_8_sva_3;
  assign _00672_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_7_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_7_sva_3;
  assign _00669_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_6_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_6_sva_3;
  assign _00664_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_4_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_4_sva_3;
  assign _00659_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_16_2_sva_2 : IntShiftRightSat_49U_6U_17U_o_16_2_sva_3;
  assign _00588_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_2_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_2_sva_3;
  assign _00592_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_4_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_4_sva_3;
  assign _00596_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_6_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_6_sva_3;
  assign _00600_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_8_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_8_sva_3;
  assign _00579_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_12_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_12_sva_3;
  assign _00965_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) cvt_14_IntSaturation_17U_8U_if_acc_3_nl[10] : cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1;
  assign _00604_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_sva_3;
  assign _00585_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_15_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_15_sva_3;
  assign _00581_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_13_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_13_sva_3;
  assign _00577_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_11_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_11_sva_3;
  assign _00598_ = IntShiftRightSat_49U_6U_17U_o_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18841" *) IntShiftRightSat_49U_6U_17U_o_0_7_sva_2 : IntShiftRightSat_49U_6U_17U_o_0_7_sva_3;
  assign _00656_ = _02043_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18810" *) IntShiftRightSat_49U_6U_17U_o_16_1_sva_3 : IntShiftRightSat_49U_6U_17U_o_16_1_sva_4;
  assign _00748_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) cfg_proc_precision_1_sva_st_65 : cfg_proc_precision_1_sva_st_66;
  assign _01005_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04891_ : cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01019_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04890_ : cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01034_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04889_ : cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01048_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04888_ : cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01064_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04887_ : cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01078_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04886_ : cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01092_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04885_ : cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01106_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04884_ : cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01121_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04883_ : cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _00913_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04882_ : cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _00926_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04881_ : cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _00939_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04880_ : cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _00952_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04879_ : cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _00966_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04878_ : cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _00979_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04877_ : cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _00992_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) _04876_ : cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  assign _01137_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) cvt_unequal_tmp_20 : cvt_unequal_tmp_21;
  assign _00735_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) cfg_mode_eql_1_sva_5 : cfg_mode_eql_1_sva_6;
  assign _00736_ = cfg_out_precision_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18751" *) cfg_out_precision_1_sva_st_113 : cfg_out_precision_1_sva_6;
  assign _00914_ = _02042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18703" *) _09058_ : cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  assign _00901_ = _02041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18687" *) _09057_ : cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  assign _00793_ = _02040_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18676" *) chn_idata_data_sva_2_335_319_1 : chn_idata_data_sva_3_335_319_1;
  assign _00927_ = _02039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18663" *) _09056_ : cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1;
  assign _00792_ = _02038_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18652" *) chn_idata_data_sva_2_303_287_1 : chn_idata_data_sva_3_303_287_1;
  assign _01108_ = _02037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18639" *) _09055_ : cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  assign _00794_ = _02036_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18628" *) chn_idata_data_sva_2_367_351_1 : chn_idata_data_sva_3_367_351_1;
  assign _00940_ = _02035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18615" *) _09054_ : cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  assign _00791_ = _02034_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18604" *) chn_idata_data_sva_2_271_255_1 : chn_idata_data_sva_3_271_255_1;
  assign _01094_ = _02033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18593" *) _09053_ : cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2;
  assign _00795_ = _02031_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18583" *) chn_idata_data_sva_2_399_383_1 : chn_idata_data_sva_3_399_383_1;
  assign _01147_ = _02030_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18575" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg;
  assign _01148_ = _02028_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18567" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg;
  assign _01311_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 : IsNaN_5U_10U_land_14_lpi_1_dfm_5;
  assign _00693_ = _02026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18557" *) _01311_ : IsNaN_5U_10U_land_14_lpi_1_dfm_6;
  assign _00953_ = _02025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18544" *) _09052_ : cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1;
  assign _01310_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 : IsNaN_5U_10U_land_7_lpi_1_dfm_5;
  assign _00706_ = _02024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18532" *) _01310_ : IsNaN_5U_10U_land_7_lpi_1_dfm_6;
  assign _00790_ = _02023_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18524" *) chn_idata_data_sva_2_239_223_1 : chn_idata_data_sva_3_239_223_1;
  assign _01080_ = _02022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18513" *) _09051_ : cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2;
  assign _00796_ = _02020_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18503" *) chn_idata_data_sva_2_431_415_1 : chn_idata_data_sva_3_431_415_1;
  assign _01149_ = _02019_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18495" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg;
  assign _01150_ = _02017_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18486" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg;
  assign _00967_ = _02014_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18474" *) _09050_ : cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2;
  assign _01141_ = and_2402_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18461" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg;
  assign _01143_ = and_2402_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18461" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg;
  assign _01161_ = and_2402_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18461" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg;
  assign _01159_ = and_2402_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18461" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg;
  assign _01164_ = and_2396_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18448" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg;
  assign _01162_ = and_2396_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18448" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg;
  assign _01160_ = and_2396_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18448" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg;
  assign _00789_ = _02012_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18438" *) chn_idata_data_sva_2_207_191_1 : chn_idata_data_sva_3_207_191_1;
  assign _01066_ = _02011_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18425" *) _09049_ : cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  assign _00797_ = _02010_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18414" *) chn_idata_data_sva_2_463_447_1 : chn_idata_data_sva_3_463_447_1;
  assign _01145_ = and_2393_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18405" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg;
  assign _01151_ = and_2393_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18405" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg;
  assign _01146_ = and_2389_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18395" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg;
  assign _01152_ = and_2389_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18395" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg;
  assign _00980_ = _02009_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18381" *) _09048_ : cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1;
  assign _01309_ = and_957_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1 : FpFloatToInt_16U_5U_10U_internal_int_0_sva_mx0w0;
  assign _00266_ = _02008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18369" *) _01309_ : FpFloatToInt_16U_5U_10U_internal_int_0_sva_3;
  assign _00788_ = _02006_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18361" *) chn_idata_data_sva_2_175_159_1 : chn_idata_data_sva_3_175_159_1;
  assign _01050_ = _02005_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18350" *) _09047_ : cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2;
  assign _00799_ = _02003_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18340" *) chn_idata_data_sva_2_495_479_1 : chn_idata_data_sva_3_495_479_1;
  assign _01163_ = and_2380_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18331" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg;
  assign _01167_ = and_2380_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18331" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg;
  assign _01142_ = and_2372_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18320" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg;
  assign _01144_ = and_2372_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18320" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg;
  assign _01168_ = and_2372_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18320" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg;
  assign _00267_ = _02002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18305" *) _09179_ : FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5;
  assign _00787_ = _02001_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18296" *) chn_idata_data_sva_2_143_127_1 : chn_idata_data_sva_3_143_127_1;
  assign _01036_ = _02000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18283" *) _09046_ : cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  assign _01165_ = and_2369_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18270" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg;
  assign _01157_ = and_2369_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18270" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg;
  assign _01155_ = and_2369_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18270" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg;
  assign _01166_ = and_2365_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18258" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg;
  assign _01158_ = and_2365_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18258" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg;
  assign _01156_ = and_2365_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18258" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg;
  assign _01401_ = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8 : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_nl;
  assign _01308_ = and_dcpl_408 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_2_511_1 : IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2;
  assign _01307_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 : IsNaN_5U_10U_land_11_lpi_1_dfm_4;
  assign _01306_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 : IsNaN_5U_10U_land_10_lpi_1_dfm_4;
  assign _01305_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 : IsNaN_5U_10U_land_12_lpi_1_dfm_4;
  assign _01304_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 : IsNaN_5U_10U_land_9_lpi_1_dfm_4;
  assign _01303_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 : IsNaN_5U_10U_land_13_lpi_1_dfm_4;
  assign _01302_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 : IsNaN_5U_10U_land_8_lpi_1_dfm_4;
  assign _01301_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 : IsNaN_5U_10U_land_6_lpi_1_dfm_4;
  assign _01300_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 : IsNaN_5U_10U_land_lpi_1_dfm_4;
  assign _01299_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 : IsNaN_5U_10U_land_5_lpi_1_dfm_4;
  assign _01298_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 : IsNaN_5U_10U_land_4_lpi_1_dfm_4;
  assign _01297_ = and_dcpl_420 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 : IsNaN_5U_10U_land_3_lpi_1_dfm_4;
  assign _00517_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01308_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3;
  assign _00268_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01401_ : FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1;
  assign _00698_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01297_ : IsNaN_5U_10U_land_3_lpi_1_dfm_5;
  assign _00702_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01299_ : IsNaN_5U_10U_land_5_lpi_1_dfm_5;
  assign _00704_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01301_ : IsNaN_5U_10U_land_6_lpi_1_dfm_5;
  assign _00710_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01304_ : IsNaN_5U_10U_land_9_lpi_1_dfm_5;
  assign _00685_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01306_ : IsNaN_5U_10U_land_10_lpi_1_dfm_5;
  assign _00689_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01305_ : IsNaN_5U_10U_land_12_lpi_1_dfm_5;
  assign _00712_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01300_ : IsNaN_5U_10U_land_lpi_1_dfm_5;
  assign _00691_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01303_ : IsNaN_5U_10U_land_13_lpi_1_dfm_5;
  assign _00687_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01307_ : IsNaN_5U_10U_land_11_lpi_1_dfm_5;
  assign _00708_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01302_ : IsNaN_5U_10U_land_8_lpi_1_dfm_5;
  assign _00700_ = IsNaN_5U_10U_aelse_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18219" *) _01298_ : IsNaN_5U_10U_land_4_lpi_1_dfm_5;
  assign _00786_ = _01999_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18199" *) chn_idata_data_sva_2_111_95_1 : chn_idata_data_sva_3_111_95_1;
  assign _01021_ = _01998_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18186" *) _09045_ : cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  assign _01153_ = _01997_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18175" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt[9:0] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg;
  assign _01154_ = _01994_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18166" *) FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt[14:10] : reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg;
  assign _01296_ = and_dcpl_424 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 : IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0;
  assign _00696_ = _01992_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18157" *) _01296_ : IsNaN_5U_10U_land_2_lpi_1_dfm_4;
  assign _00800_ = _01991_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18149" *) chn_idata_data_sva_2_79_63_1 : chn_idata_data_sva_3_79_63_1;
  assign _01007_ = _01990_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18136" *) _09044_ : cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  assign _01295_ = and_dcpl_424 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2 : IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0;
  assign _01294_ = and_dcpl_424 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 : IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0;
  assign _00694_ = IsNaN_5U_10U_aelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18120" *) _01295_ : IsNaN_5U_10U_land_15_lpi_1_dfm_3;
  assign _00695_ = IsNaN_5U_10U_aelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18120" *) _01294_ : IsNaN_5U_10U_land_1_lpi_1_dfm_3;
  assign _01022_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] : cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  assign _01051_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] : cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  assign _01067_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] : cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  assign _01109_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] : cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  assign _00902_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] : cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  assign _00928_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] : cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  assign _00968_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] : cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  assign _00981_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11] : cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2;
  assign _00954_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] : cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  assign _00941_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] : cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  assign _00915_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] : cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  assign _01095_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11] : cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  assign _01081_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] : cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  assign _01037_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11] : cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  assign _01008_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11] : cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  assign _00994_ = FpFloatToInt_16U_5U_10U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18080" *) cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl[11] : cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2;
  assign _00798_ = _01989_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18041" *) chn_idata_data_sva_2_47_31_1 : chn_idata_data_sva_3_47_31_1;
  assign _00993_ = _01988_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:18030" *) _09043_ : cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2;
  assign _00257_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09028_ : FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  assign _00258_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09029_ : FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  assign _00259_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09030_ : FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  assign _00260_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09031_ : FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  assign _00261_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09032_ : FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  assign _00262_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09033_ : FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  assign _00263_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09035_ : FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  assign _00264_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09037_ : FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  assign _00265_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09039_ : FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  assign _00251_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09041_ : FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  assign _00252_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09042_ : FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  assign _00253_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09040_ : FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  assign _00254_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09038_ : FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  assign _00255_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09036_ : FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  assign _00256_ = FpFloatToInt_16U_5U_10U_internal_int_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17976" *) _09034_ : FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  assign _01140_ = _01986_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17954" *) _04874_ : main_stage_v_3;
  assign _00749_ = cfg_proc_precision_and_27_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17944" *) reg_cfg_proc_precision_1_sva_st_40_cse : cfg_proc_precision_1_sva_st_89;
  assign _01006_ = cfg_proc_precision_and_27_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17944" *) cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp : cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2;
  assign _00743_ = cfg_proc_precision_and_24_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17932" *) reg_cfg_proc_precision_1_sva_st_40_cse : cfg_proc_precision_1_sva_st_101;
  assign _01122_ = cfg_proc_precision_and_24_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17932" *) cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp : cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2;
  assign _00740_ = _01985_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17922" *) cfg_out_precision_1_sva_st_154 : cfg_out_precision_1_sva_st_149;
  assign _00985_ = _01984_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17913" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[16] : cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2;
  assign _01293_ = and_881_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[0];
  assign _00284_ = _01983_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17903" *) _01293_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9;
  assign _01191_ = _01979_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17894" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg;
  assign _01421_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_sva : IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0;
  assign _00636_ = _01978_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17885" *) _01421_ : IntShiftRightSat_49U_6U_17U_o_15_1_sva_2;
  assign _01292_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_sva : IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0;
  assign _00679_ = _01977_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17875" *) _01292_ : IntShiftRightSat_49U_6U_17U_o_16_sva_2;
  assign _00558_ = _01976_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17866" *) IntShiftRightSat_49U_6U_17U_i_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_sva_2;
  assign _00972_ = _01975_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17857" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[16] : cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  assign _01291_ = and_866_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[0];
  assign _00274_ = _01974_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17847" *) _01291_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8;
  assign _01179_ = _01970_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17838" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg;
  assign _01420_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_15_sva : IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0;
  assign _00616_ = _01969_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17829" *) _01420_ : IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2;
  assign _01290_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_15_sva : IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0;
  assign _00653_ = _01968_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17819" *) _01290_ : IntShiftRightSat_49U_6U_17U_o_16_15_sva_2;
  assign _00548_ = _01967_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17810" *) IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_15_sva_2;
  assign _00958_ = _01966_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17801" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[16] : cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  assign _01289_ = and_849_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[0];
  assign _00273_ = _01965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17791" *) _01289_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8;
  assign _01177_ = _01961_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17782" *) FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg;
  assign _01178_ = _01960_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17774" *) FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg;
  assign _01419_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_14_sva : IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0;
  assign _00614_ = _01957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17764" *) _01419_ : IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2;
  assign _01288_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm : IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0;
  assign _01287_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_14_sva : IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0;
  assign _00512_ = IntShiftRightSat_49U_6U_17U_o_and_90_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17752" *) _01288_ : IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3;
  assign _00650_ = IntShiftRightSat_49U_6U_17U_o_and_90_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17752" *) _01287_ : IntShiftRightSat_49U_6U_17U_o_16_14_sva_2;
  assign _00547_ = _01956_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17743" *) IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_14_sva_2;
  assign _00945_ = _01955_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17734" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[16] : cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  assign _01286_ = and_830_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[0];
  assign _00272_ = _01954_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17724" *) _01286_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7;
  assign _01418_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_13_sva : IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0;
  assign _00612_ = _01950_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17714" *) _01418_ : IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2;
  assign _01285_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_13_sva : IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0;
  assign _00647_ = _01949_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17704" *) _01285_ : IntShiftRightSat_49U_6U_17U_o_16_13_sva_2;
  assign _00546_ = _01948_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17695" *) IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_13_sva_2;
  assign _00932_ = _01947_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17686" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[16] : cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  assign _01284_ = and_816_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[0];
  assign _00271_ = _01946_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17676" *) _01284_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8;
  assign _01175_ = and_2317_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17666" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg;
  assign _01173_ = and_2317_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17666" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg;
  assign _01417_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_12_sva : IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0;
  assign _00610_ = _01942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17656" *) _01417_ : IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2;
  assign _01283_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_12_sva : IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0;
  assign _00644_ = _01941_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17646" *) _01283_ : IntShiftRightSat_49U_6U_17U_o_16_12_sva_2;
  assign _00545_ = _01940_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17637" *) IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_12_sva_2;
  assign _00919_ = _01939_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17628" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[16] : cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  assign _01282_ = and_801_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[0];
  assign _00270_ = _01938_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17618" *) _01282_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7;
  assign _01416_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_11_sva : IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0;
  assign _00608_ = _01934_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17608" *) _01416_ : IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2;
  assign _01281_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_11_sva : IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0;
  assign _00641_ = _01933_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17598" *) _01281_ : IntShiftRightSat_49U_6U_17U_o_16_11_sva_2;
  assign _00544_ = _01932_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17589" *) IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_11_sva_2;
  assign _00906_ = _01931_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17580" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[16] : cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  assign _01280_ = and_787_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[0];
  assign _00269_ = _01930_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17570" *) _01280_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7;
  assign _01415_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_10_sva : IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0;
  assign _00606_ = _01926_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17560" *) _01415_ : IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2;
  assign _01279_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_10_sva : IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0;
  assign _00638_ = _01925_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17550" *) _01279_ : IntShiftRightSat_49U_6U_17U_o_16_10_sva_2;
  assign _00543_ = _01924_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17541" *) IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_10_sva_2;
  assign _01112_ = _01923_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17532" *) cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _01113_ = _01922_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17522" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[16] : cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  assign _01278_ = and_dcpl_301 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[0];
  assign _01414_ = and_dcpl_301 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[15:1];
  assign _00283_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17510" *) _01278_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6;
  assign _00288_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17510" *) _01414_ : FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6;
  assign _01413_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_9_sva : IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0;
  assign _00634_ = _01921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17500" *) _01413_ : IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2;
  assign _00557_ = _01920_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17491" *) IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_i_9_sva_2;
  assign _01065_ = _01919_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17482" *) cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp : cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  assign _01107_ = _01918_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17472" *) cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp : cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2;
  assign _01099_ = _01917_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17462" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[16] : cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  assign _01277_ = and_766_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[0];
  assign _00282_ = _01916_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17452" *) _01277_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8;
  assign _01189_ = and_2259_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17443" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg;
  assign _01412_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_8_sva : IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0;
  assign _00632_ = _01912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17434" *) _01412_ : IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2;
  assign _01276_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_8_sva : IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0;
  assign _00674_ = _01911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17424" *) _01276_ : IntShiftRightSat_49U_6U_17U_o_16_8_sva_2;
  assign _00556_ = _01910_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17415" *) IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_8_sva_2;
  assign _01085_ = _01909_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17406" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[16] : cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  assign _01275_ = and_749_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[0];
  assign _00281_ = _01908_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17396" *) _01275_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7;
  assign _01411_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_7_sva : IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0;
  assign _00630_ = _01904_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17386" *) _01411_ : IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2;
  assign _01274_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_7_sva : IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0;
  assign _00671_ = _01903_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17376" *) _01274_ : IntShiftRightSat_49U_6U_17U_o_16_7_sva_2;
  assign _00555_ = _01902_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17367" *) IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_7_sva_2;
  assign _01093_ = IntShiftRightSat_49U_6U_17U_if_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17356" *) cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign _01079_ = IntShiftRightSat_49U_6U_17U_if_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17356" *) cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign _01071_ = _01901_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17344" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[16] : cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  assign _01273_ = and_734_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[0];
  assign _00280_ = _01900_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17334" *) _01273_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7;
  assign _01187_ = and_2275_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17324" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg;
  assign _01185_ = and_2275_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17324" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg;
  assign _01410_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_6_sva : IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0;
  assign _00628_ = _01896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17314" *) _01410_ : IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2;
  assign _01272_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_6_sva : IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0;
  assign _00668_ = _01895_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17304" *) _01272_ : IntShiftRightSat_49U_6U_17U_o_16_6_sva_2;
  assign _00554_ = _01894_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17295" *) IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_6_sva_2;
  assign _01055_ = _01893_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17286" *) cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _01056_ = _01892_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17276" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[16] : cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  assign _01271_ = and_719_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[0];
  assign _00279_ = _01891_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17266" *) _01271_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6;
  assign _01183_ = _01887_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17257" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg;
  assign _01409_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_5_sva : IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0;
  assign _00626_ = _01886_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17248" *) _01409_ : IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2;
  assign _00553_ = _01885_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17239" *) IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_i_5_sva_2;
  assign _01049_ = _01884_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17230" *) cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp : cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign _01041_ = _01883_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17220" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[16] : cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  assign _01270_ = and_704_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[0];
  assign _00278_ = _01882_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17210" *) _01270_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7;
  assign _01171_ = and_2259_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17199" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg;
  assign _01169_ = and_2259_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17199" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg;
  assign _01181_ = and_2259_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17199" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt[9:0] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg;
  assign _01192_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg;
  assign _01180_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg;
  assign _01176_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg;
  assign _01174_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg;
  assign _01172_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg;
  assign _01170_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg;
  assign _01190_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg;
  assign _01188_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg;
  assign _01186_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg;
  assign _01184_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg;
  assign _01182_ = and_2257_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17179" *) FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt[14:10] : reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg;
  assign _01408_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_4_sva : IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0;
  assign _00624_ = _01878_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17160" *) _01408_ : IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2;
  assign _01269_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_4_sva : IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0;
  assign _00663_ = _01877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17150" *) _01269_ : IntShiftRightSat_49U_6U_17U_o_16_4_sva_2;
  assign _00552_ = _01876_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17141" *) IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1 : IntShiftRightSat_49U_6U_17U_i_4_sva_2;
  assign _01025_ = _01875_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17132" *) cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _01026_ = _01874_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17122" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[16] : cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  assign _01268_ = and_dcpl_224 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[0];
  assign _01407_ = and_dcpl_224 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[15:1];
  assign _00277_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17110" *) _01268_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6;
  assign _00287_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17110" *) _01407_ : FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6;
  assign _01406_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_3_sva : IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0;
  assign _00622_ = _01873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17100" *) _01406_ : IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2;
  assign _00551_ = _01872_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17091" *) IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_i_3_sva_2;
  assign _01035_ = IntShiftRightSat_49U_6U_17U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17080" *) cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp : cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  assign _01020_ = IntShiftRightSat_49U_6U_17U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17080" *) cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp : cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  assign _01011_ = _01871_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17068" *) cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp : cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign _01012_ = _01870_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17058" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[16] : cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  assign _01267_ = and_dcpl_217 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[0];
  assign _01405_ = and_dcpl_217 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[15:1];
  assign _00276_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17046" *) _01267_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6;
  assign _00286_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17046" *) _01405_ : FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6;
  assign _01404_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_2_sva : IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0;
  assign _00620_ = _01869_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17036" *) _01404_ : IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2;
  assign _01266_ = and_685_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_16_2_sva : IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0;
  assign _00658_ = _01868_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17026" *) _01266_ : IntShiftRightSat_49U_6U_17U_o_16_2_sva_2;
  assign _00550_ = _01866_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17017" *) IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_i_2_sva_2;
  assign _00996_ = _01865_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17009" *) cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp : cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign _00997_ = _01864_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:17000" *) FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[16] : cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2;
  assign _01265_ = and_dcpl_209 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[0];
  assign _01403_ = and_dcpl_209 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0 : FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[15:1];
  assign _00275_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16988" *) _01265_ : FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5;
  assign _00285_ = FpIntToFloat_17U_5U_10U_else_i_abs_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16988" *) _01403_ : FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5;
  assign _01402_ = and_dcpl_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24473|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24472" *) IntShiftRightSat_49U_6U_17U_o_15_1_1_sva : IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0;
  assign _00618_ = _01863_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16978" *) _01402_ : IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2;
  assign _00549_ = _01861_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16969" *) IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_i_1_sva_2;
  assign _00982_ = _01860_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16961" *) nl_cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2 : cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2;
  assign _01400_ = and_668_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1 : chn_idata_data_sva_1_507_479_1[10:1];
  assign _00491_ = _01859_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16951" *) _01400_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9;
  assign _00784_ = _01856_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16942" *) chn_idata_data_sva_1_511_1 : chn_idata_data_sva_2_511_1;
  assign _01399_ = and_666_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1 : chn_idata_data_sva_1_475_447_1[10:1];
  assign _00481_ = _01855_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16932" *) _01399_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8;
  assign _01398_ = and_664_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1 : chn_idata_data_sva_1_443_415_1[10:1];
  assign _00480_ = _01852_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16921" *) _01398_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8;
  assign _01397_ = and_662_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1 : chn_idata_data_sva_1_411_383_1[10:1];
  assign _00479_ = _01849_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16910" *) _01397_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8;
  assign _01396_ = and_660_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1 : chn_idata_data_sva_1_379_351_1[10:1];
  assign _00478_ = _01846_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16899" *) _01396_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8;
  assign _01395_ = and_658_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1 : chn_idata_data_sva_1_347_319_1[10:1];
  assign _00477_ = _01843_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16888" *) _01395_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8;
  assign _01394_ = and_656_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1 : chn_idata_data_sva_1_315_287_1[10:1];
  assign _00476_ = _01840_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16877" *) _01394_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8;
  assign _00955_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16866" *) nl_cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 : cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign _00929_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16866" *) nl_cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 : cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign _01110_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16866" *) nl_cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0] : cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign _01393_ = and_654_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1 : chn_idata_data_sva_1_283_255_1[10:1];
  assign _00490_ = _01837_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16854" *) _01393_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8;
  assign _01392_ = and_652_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1 : chn_idata_data_sva_1_251_223_1[10:1];
  assign _00489_ = _01834_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16843" *) _01392_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8;
  assign _01391_ = and_650_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1 : chn_idata_data_sva_1_219_191_1[10:1];
  assign _00488_ = _01831_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16832" *) _01391_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8;
  assign _00969_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16817" *) nl_cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 : cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign _00942_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16817" *) nl_cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 : cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign _00916_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16817" *) nl_cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 : cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign _00903_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16817" *) nl_cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 : cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign _01096_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16817" *) nl_cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2[4:0] : cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign _01082_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16817" *) nl_cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0] : cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign _01068_ = FpFloatToInt_16U_5U_10U_shift_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16817" *) nl_cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0] : cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign _01390_ = and_648_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1 : chn_idata_data_sva_1_187_159_1[10:1];
  assign _00487_ = _01828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16801" *) _01390_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8;
  assign _01052_ = _01825_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16792" *) nl_cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0] : cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign _01389_ = and_646_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1 : chn_idata_data_sva_1_155_127_1[10:1];
  assign _00486_ = _01824_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16782" *) _01389_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8;
  assign _01388_ = and_643_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1 : chn_idata_data_sva_1_123_95_1[10:1];
  assign _00485_ = _01821_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16771" *) _01388_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8;
  assign _01387_ = and_641_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1 : chn_idata_data_sva_1_91_63_1[10:1];
  assign _00484_ = _01818_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16760" *) _01387_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8;
  assign _01038_ = FpFloatToInt_16U_5U_10U_shift_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16749" *) nl_cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 : cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign _01023_ = FpFloatToInt_16U_5U_10U_shift_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16749" *) nl_cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 : cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign _01009_ = FpFloatToInt_16U_5U_10U_shift_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16749" *) nl_cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 : cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign _01386_ = and_639_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1 : chn_idata_data_sva_1_59_31_1[10:1];
  assign _00483_ = _01815_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16737" *) _01386_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8;
  assign _00995_ = _01812_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16728" *) nl_cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2 : cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2;
  assign _01385_ = and_637_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24456|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24455" *) FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1 : chn_idata_data_sva_1_27_0_1[9:0];
  assign _00482_ = _01811_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16718" *) _01385_ : FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8;
  assign _00782_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_59_31_1[16:0] : chn_idata_data_sva_2_47_31_1;
  assign _00785_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_91_63_1[16:0] : chn_idata_data_sva_2_79_63_1;
  assign _00769_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_123_95_1[16:0] : chn_idata_data_sva_2_111_95_1;
  assign _00770_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_155_127_1[16:0] : chn_idata_data_sva_2_143_127_1;
  assign _00772_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_187_159_1[16:0] : chn_idata_data_sva_2_175_159_1;
  assign _00773_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_219_191_1[16:0] : chn_idata_data_sva_2_207_191_1;
  assign _00774_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_251_223_1[16:0] : chn_idata_data_sva_2_239_223_1;
  assign _00775_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_283_255_1[16:0] : chn_idata_data_sva_2_271_255_1;
  assign _00776_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_315_287_1[16:0] : chn_idata_data_sva_2_303_287_1;
  assign _00777_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_347_319_1[16:0] : chn_idata_data_sva_2_335_319_1;
  assign _00778_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_379_351_1[16:0] : chn_idata_data_sva_2_367_351_1;
  assign _00779_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_411_383_1[16:0] : chn_idata_data_sva_2_399_383_1;
  assign _00780_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_443_415_1[16:0] : chn_idata_data_sva_2_431_415_1;
  assign _00781_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_475_447_1[16:0] : chn_idata_data_sva_2_463_447_1;
  assign _00783_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) chn_idata_data_sva_1_507_479_1[16:0] : chn_idata_data_sva_2_495_479_1;
  assign _00473_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1;
  assign _00474_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1;
  assign _00443_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1;
  assign _00444_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1;
  assign _00440_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1;
  assign _00441_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1;
  assign _00437_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1;
  assign _00438_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1;
  assign _00434_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1;
  assign _00435_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1;
  assign _00431_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1;
  assign _00432_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1;
  assign _00428_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1;
  assign _00429_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1;
  assign _00470_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1;
  assign _00471_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1;
  assign _00467_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1;
  assign _00468_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1;
  assign _00464_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1;
  assign _00465_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1;
  assign _00461_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1;
  assign _00462_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1;
  assign _00458_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1;
  assign _00459_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1;
  assign _00455_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1;
  assign _00456_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1;
  assign _00452_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1;
  assign _00453_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1;
  assign _00449_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1;
  assign _00450_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1;
  assign _00446_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1;
  assign _00447_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1;
  assign _00737_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) cfg_out_precision_1_sva_st_154 : cfg_out_precision_1_sva_st_113;
  assign _00747_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) cfg_proc_precision_1_sva_st_64 : cfg_proc_precision_1_sva_st_65;
  assign _01136_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) cvt_unequal_tmp_19 : cvt_unequal_tmp_20;
  assign _00734_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) cfg_mode_eql_1_sva_4 : cfg_mode_eql_1_sva_5;
  assign _00587_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_2_sva_2;
  assign _00591_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_4_sva_2;
  assign _00595_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_6_sva_2;
  assign _00599_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_8_sva_2;
  assign _00575_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_10_sva_2;
  assign _00578_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_12_sva_2;
  assign _00582_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_14_sva_3;
  assign _00603_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_sva_2;
  assign _00660_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_3_sva_3;
  assign _00665_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_5_sva_3;
  assign _00676_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_9_sva_3;
  assign _00655_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_16_1_sva_3;
  assign _00589_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_3_sva_3;
  assign _00697_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04816_ : IsNaN_5U_10U_land_3_lpi_1_dfm_4;
  assign _00593_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_5_sva_3;
  assign _00701_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04822_ : IsNaN_5U_10U_land_5_lpi_1_dfm_4;
  assign _00703_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04825_ : IsNaN_5U_10U_land_6_lpi_1_dfm_4;
  assign _00601_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_9_sva_3;
  assign _00709_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04834_ : IsNaN_5U_10U_land_9_lpi_1_dfm_4;
  assign _00684_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04837_ : IsNaN_5U_10U_land_10_lpi_1_dfm_4;
  assign _00688_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04843_ : IsNaN_5U_10U_land_12_lpi_1_dfm_4;
  assign _00584_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_15_sva_2;
  assign _00711_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04852_ : IsNaN_5U_10U_land_lpi_1_dfm_4;
  assign _00692_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04849_ : IsNaN_5U_10U_land_14_lpi_1_dfm_5;
  assign _00580_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_13_sva_2;
  assign _00690_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04846_ : IsNaN_5U_10U_land_13_lpi_1_dfm_4;
  assign _00576_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_11_sva_2;
  assign _00686_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04840_ : IsNaN_5U_10U_land_11_lpi_1_dfm_4;
  assign _00707_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04831_ : IsNaN_5U_10U_land_8_lpi_1_dfm_4;
  assign _00597_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_7_sva_2;
  assign _00705_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04828_ : IsNaN_5U_10U_land_7_lpi_1_dfm_5;
  assign _00699_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) _04819_ : IsNaN_5U_10U_land_4_lpi_1_dfm_4;
  assign _00586_ = chn_idata_data_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16613" *) IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0 : IntShiftRightSat_49U_6U_17U_o_0_1_sva_2;
  assign _01139_ = _01795_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16522" *) _04813_ : main_stage_v_2;
  assign _01227_ = cfg_proc_precision_and_11_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16512" *) cfg_proc_precision_rsci_d : reg_cfg_proc_precision_1_sva_st_40_cse;
  assign _00498_ = cfg_proc_precision_and_11_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16512" *) _04005_ : IntMulExt_33U_16U_49U_return_1_sva_2;
  assign _00741_ = _01794_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16503" *) cfg_out_precision_rsci_d : cfg_out_precision_1_sva_st_154;
  assign _00502_ = _01793_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16494" *) _04004_ : IntMulExt_33U_16U_49U_return_5_sva_2;
  assign _01432_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1 : cvt_13_IntMulExt_33U_16U_49U_o_mul_2_nl;
  assign _01431_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1 : cvt_15_IntMulExt_33U_16U_49U_o_mul_3_nl;
  assign _01430_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_sva_mx0w1 : cvt_16_IntMulExt_33U_16U_49U_o_mul_4_nl;
  assign _01429_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1 : cvt_14_IntMulExt_33U_16U_49U_o_mul_3_nl;
  assign _01428_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1 : cvt_11_IntMulExt_33U_16U_49U_o_mul_2_nl;
  assign _01427_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1 : cvt_12_IntMulExt_33U_16U_49U_o_mul_3_nl;
  assign _01426_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1 : cvt_10_IntMulExt_33U_16U_49U_o_mul_2_nl;
  assign _01425_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1 : cvt_7_IntMulExt_33U_16U_49U_o_mul_2_nl;
  assign _01424_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1 : cvt_8_IntMulExt_33U_16U_49U_o_mul_3_nl;
  assign _01423_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1 : cvt_6_IntMulExt_33U_16U_49U_o_mul_2_nl;
  assign _00507_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01430_ : IntMulExt_33U_16U_49U_return_sva_1;
  assign _00497_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01431_ : IntMulExt_33U_16U_49U_return_15_sva_1;
  assign _00496_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01429_ : IntMulExt_33U_16U_49U_return_14_sva_1;
  assign _00495_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01432_ : IntMulExt_33U_16U_49U_return_13_sva_1;
  assign _00494_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01427_ : IntMulExt_33U_16U_49U_return_12_sva_1;
  assign _00493_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01428_ : IntMulExt_33U_16U_49U_return_11_sva_1;
  assign _00492_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01426_ : IntMulExt_33U_16U_49U_return_10_sva_1;
  assign _00505_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01424_ : IntMulExt_33U_16U_49U_return_8_sva_1;
  assign _00504_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01425_ : IntMulExt_33U_16U_49U_return_7_sva_1;
  assign _00503_ = IntMulExt_33U_16U_49U_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16467" *) _01423_ : IntMulExt_33U_16U_49U_return_6_sva_1;
  assign _01422_ = IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24524|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24523" *) IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1 : cvt_4_IntMulExt_33U_16U_49U_o_mul_2_nl;
  assign _00501_ = _01792_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16449" *) _01422_ : IntMulExt_33U_16U_49U_return_4_sva_1;
  assign _00506_ = IntMulExt_33U_16U_49U_and_11_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16435" *) _04003_ : IntMulExt_33U_16U_49U_return_9_sva_2;
  assign _00500_ = IntMulExt_33U_16U_49U_and_11_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16435" *) _04002_ : IntMulExt_33U_16U_49U_return_3_sva_2;
  assign _00499_ = IntMulExt_33U_16U_49U_and_11_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16435" *) _04001_ : IntMulExt_33U_16U_49U_return_2_sva_2;
  assign _00991_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl[8] : cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2;
  assign _00978_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] : cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign _00964_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] : cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign _00951_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] : cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign _00938_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] : cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign _00925_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] : cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign _00912_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] : cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign _01119_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] : cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign _01105_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8] : cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign _01091_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] : cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign _01077_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] : cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign _01062_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] : cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign _01047_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8] : cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign _01032_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] : cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign _01018_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8] : cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign _01003_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8] : cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2;
  assign _00417_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04782_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2;
  assign _00416_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04784_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2;
  assign _00415_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04786_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2;
  assign _00414_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04788_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2;
  assign _00413_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04790_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2;
  assign _00412_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04792_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2;
  assign _00426_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04794_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2;
  assign _00425_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04796_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2;
  assign _00424_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04798_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2;
  assign _00423_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04800_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2;
  assign _00422_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04802_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2;
  assign _00716_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp : IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2;
  assign _00732_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_nor_4_tmp : IsNaN_8U_23U_nor_4_itm_2;
  assign _00421_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04804_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2;
  assign _00420_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04806_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2;
  assign _00419_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04808_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2;
  assign _00418_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04810_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2;
  assign _00427_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) _04812_ : FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2;
  assign _00731_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp : IsNaN_8U_23U_land_lpi_1_dfm_3;
  assign _00722_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp : IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  assign _00721_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp : IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  assign _00720_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp : IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  assign _00719_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp : IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  assign _00718_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp : IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  assign _00717_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp : IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  assign _00730_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp : IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  assign _00729_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp : IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  assign _00728_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp : IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  assign _00727_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp : IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  assign _00726_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp : IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  assign _00725_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp : IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  assign _00724_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp : IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  assign _00723_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp : IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  assign _00392_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2;
  assign _01001_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8] : cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2;
  assign _00394_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2;
  assign _01016_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _00396_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2;
  assign _01030_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _00398_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2;
  assign _01045_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _00400_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2;
  assign _01060_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _00402_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2;
  assign _01075_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _00404_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2;
  assign _01089_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _00406_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2;
  assign _01103_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _00408_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2;
  assign _01117_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  assign _00380_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2;
  assign _00910_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _00382_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2;
  assign _00923_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _00384_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2;
  assign _00936_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _00386_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2;
  assign _00949_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  assign _00388_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2;
  assign _00962_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _00390_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2;
  assign _00976_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  assign _00410_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2;
  assign _00989_ = FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16265" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8] : cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2;
  assign _00411_ = _01742_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16128" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2;
  assign _00990_ = _01741_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16118" *) cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8] : cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2;
  assign _00371_ = _01740_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16109" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2;
  assign _00391_ = _01739_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16100" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2;
  assign _00977_ = _01738_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16090" *) cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _00370_ = _01737_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16081" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2;
  assign _00389_ = _01736_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16072" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2;
  assign _00963_ = _01735_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16062" *) cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _00369_ = _01734_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16053" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2;
  assign _00387_ = _01733_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16044" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2;
  assign _00950_ = _01732_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16034" *) cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _00368_ = _01731_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16025" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2;
  assign _00385_ = _01730_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16016" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2;
  assign _00937_ = _01729_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:16006" *) cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _00367_ = _01728_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15997" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2;
  assign _00383_ = _01727_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15988" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2;
  assign _00924_ = _01726_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15978" *) cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _00366_ = _01725_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15969" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2;
  assign _00381_ = _01724_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15960" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2;
  assign _00911_ = _01723_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15950" *) cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _00365_ = _01722_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15941" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2;
  assign _00409_ = _01721_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15932" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2;
  assign _01118_ = _01720_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15922" *) cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _00364_ = _01719_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15913" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2;
  assign _00407_ = _01718_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15904" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2;
  assign _01104_ = _01717_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15894" *) cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8] : cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  assign _00379_ = _01716_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15885" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2;
  assign _00405_ = _01715_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15876" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2;
  assign _01090_ = _01714_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15866" *) cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _00378_ = _01713_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15857" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2;
  assign _00403_ = _01712_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15848" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2;
  assign _01076_ = _01711_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15838" *) cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _00377_ = _01710_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15829" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2;
  assign _00401_ = _01709_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15820" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2;
  assign _01061_ = _01708_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15810" *) cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _00376_ = _01707_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15801" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2;
  assign _00399_ = _01706_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15792" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2;
  assign _01046_ = _01705_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15782" *) cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8] : cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  assign _00375_ = _01704_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15773" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2;
  assign _00397_ = _01703_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15764" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2;
  assign _01031_ = _01702_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15754" *) cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _00374_ = _01701_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15745" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2;
  assign _00395_ = _01700_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15736" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2;
  assign _01017_ = _01699_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15726" *) cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8] : cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  assign _00767_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[59:31] : chn_idata_data_sva_1_59_31_1;
  assign _00768_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[91:63] : chn_idata_data_sva_1_91_63_1;
  assign _00752_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[123:95] : chn_idata_data_sva_1_123_95_1;
  assign _00753_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[155:127] : chn_idata_data_sva_1_155_127_1;
  assign _00754_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[187:159] : chn_idata_data_sva_1_187_159_1;
  assign _00755_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[219:191] : chn_idata_data_sva_1_219_191_1;
  assign _00756_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[251:223] : chn_idata_data_sva_1_251_223_1;
  assign _00758_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[283:255] : chn_idata_data_sva_1_283_255_1;
  assign _00759_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[315:287] : chn_idata_data_sva_1_315_287_1;
  assign _00760_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[347:319] : chn_idata_data_sva_1_347_319_1;
  assign _00761_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[379:351] : chn_idata_data_sva_1_379_351_1;
  assign _00762_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[411:383] : chn_idata_data_sva_1_411_383_1;
  assign _00763_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[443:415] : chn_idata_data_sva_1_443_415_1;
  assign _00764_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[475:447] : chn_idata_data_sva_1_475_447_1;
  assign _00765_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) chn_in_rsci_d_mxwt[507:479] : chn_idata_data_sva_1_507_479_1;
  assign _00746_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) cfg_proc_precision_rsci_d : cfg_proc_precision_1_sva_st_64;
  assign _01135_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) cvt_cvt_nand_cse : cvt_unequal_tmp_19;
  assign _00733_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) cfg_mode_eql_rsci_d : cfg_mode_eql_1_sva_4;
  assign _00751_ = chn_idata_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15699" *) cfg_truncate_rsci_d : cfg_truncate_1_sva_2;
  assign _00373_ = _01698_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15673" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2;
  assign _00393_ = _01697_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15664" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7] : FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2;
  assign _01002_ = _01696_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15654" *) cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8] : cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2;
  assign _00757_ = _01695_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15645" *) chn_in_rsci_d_mxwt[27:0] : chn_idata_data_sva_1_27_0_1;
  assign _00372_ = _01694_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15637" *) FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0 : FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2;
  assign _01138_ = _01693_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15629" *) _04743_ : main_stage_v_1;
  assign _01231_ = _01692_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15621" *) _04742_ : reg_chn_out_rsci_ld_core_psct_cse;
  assign _01264_ = and_dcpl_102 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2341_nl : chn_idata_data_sva_3_495_479_1[16];
  assign _01263_ = and_dcpl_102 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2340_nl : chn_idata_data_sva_3_495_479_1[1];
  assign _00853_ = chn_out_and_77_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15610" *) _01263_ : chn_out_rsci_d_240;
  assign _00857_ = chn_out_and_77_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15610" *) _01264_ : chn_out_rsci_d_255;
  assign _01262_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_463_447_1[16] : cvt_mux_2356_nl;
  assign _01261_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2337_nl : cvt_mux_2336_nl;
  assign _01260_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_431_415_1[16] : cvt_mux_2368_nl;
  assign _01259_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2333_nl : cvt_mux_2332_nl;
  assign _01258_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_399_383_1[16] : cvt_mux_2372_nl;
  assign _01257_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2329_nl : cvt_mux_2328_nl;
  assign _01256_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_367_351_1[16] : cvt_mux_2370_nl;
  assign _01255_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2325_nl : cvt_mux_2324_nl;
  assign _01254_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_335_319_1[16] : cvt_mux_2366_nl;
  assign _01253_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2321_nl : cvt_mux_2320_nl;
  assign _01252_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_303_287_1[16] : cvt_mux_2364_nl;
  assign _01251_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2317_nl : cvt_mux_2316_nl;
  assign _01250_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_271_255_1[16] : cvt_mux_2362_nl;
  assign _01249_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2313_nl : cvt_mux_2312_nl;
  assign _01248_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_239_223_1[16] : cvt_mux_2360_nl;
  assign _01247_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2309_nl : cvt_mux_2308_nl;
  assign _01246_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_207_191_1[16] : cvt_mux_2358_nl;
  assign _01245_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2305_nl : cvt_mux_2304_nl;
  assign _01244_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_175_159_1[16] : cvt_mux_2354_nl;
  assign _01243_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2301_nl : cvt_mux_2300_nl;
  assign _01242_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_143_127_1[16] : cvt_mux_2352_nl;
  assign _01241_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2297_nl : cvt_mux_2296_nl;
  assign _01240_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_111_95_1[16] : cvt_mux_2350_nl;
  assign _01239_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2293_nl : cvt_mux_2292_nl;
  assign _01238_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_79_63_1[16] : cvt_mux_2348_nl;
  assign _01237_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2289_nl : cvt_mux_2288_nl;
  assign _01236_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) chn_idata_data_sva_3_47_31_1[16] : cvt_mux_2346_nl;
  assign _01235_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2285_nl : cvt_mux_2284_nl;
  assign _01234_ = cfg_mode_eql_1_sva_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) reg_chn_idata_data_sva_3_15_0_reg : cvt_mux_2373_nl;
  assign _01233_ = and_dcpl_98 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24439|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:24438" *) cvt_mux_2281_nl : cvt_mux_2280_nl;
  assign _00826_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01234_ : chn_out_rsci_d_15;
  assign _00829_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01235_ : chn_out_rsci_d_16;
  assign _00882_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01238_ : chn_out_rsci_d_47;
  assign _00883_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01239_ : chn_out_rsci_d_48;
  assign _00892_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01242_ : chn_out_rsci_d_79;
  assign _00893_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01243_ : chn_out_rsci_d_80;
  assign _00808_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01246_ : chn_out_rsci_d_111;
  assign _00809_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01247_ : chn_out_rsci_d_112;
  assign _00814_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01249_ : chn_out_rsci_d_128;
  assign _00819_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01250_ : chn_out_rsci_d_143;
  assign _00820_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01251_ : chn_out_rsci_d_144;
  assign _00825_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01252_ : chn_out_rsci_d_159;
  assign _00827_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01253_ : chn_out_rsci_d_160;
  assign _00832_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01254_ : chn_out_rsci_d_175;
  assign _00833_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01255_ : chn_out_rsci_d_176;
  assign _00837_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01256_ : chn_out_rsci_d_191;
  assign _00838_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01257_ : chn_out_rsci_d_192;
  assign _00842_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01258_ : chn_out_rsci_d_207;
  assign _00843_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01259_ : chn_out_rsci_d_208;
  assign _00847_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01260_ : chn_out_rsci_d_223;
  assign _00848_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01261_ : chn_out_rsci_d_224;
  assign _00852_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01262_ : chn_out_rsci_d_239;
  assign _00804_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01233_ : chn_out_rsci_d_0;
  assign _00877_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01236_ : chn_out_rsci_d_31;
  assign _00878_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01237_ : chn_out_rsci_d_32;
  assign _00887_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01240_ : chn_out_rsci_d_63;
  assign _00888_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01241_ : chn_out_rsci_d_64;
  assign _00897_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01244_ : chn_out_rsci_d_95;
  assign _00898_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01245_ : chn_out_rsci_d_96;
  assign _00813_ = chn_out_and_32_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15557" *) _01248_ : chn_out_rsci_d_127;
  assign _00850_ = _01691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15515" *) _09357_ : chn_out_rsci_d_237_234;
  assign _00845_ = and_3063_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15495" *) _09355_ : chn_out_rsci_d_221_218;
  assign _00855_ = and_3063_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15495" *) _09356_ : chn_out_rsci_d_253_250;
  assign _00840_ = _01689_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15481" *) _09354_ : chn_out_rsci_d_205_202;
  assign _00835_ = _01687_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15467" *) _09353_ : chn_out_rsci_d_189_186;
  assign _00830_ = _01685_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15453" *) _09352_ : chn_out_rsci_d_173_170;
  assign _00823_ = _01683_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15439" *) _09351_ : chn_out_rsci_d_157_154;
  assign _00811_ = _01681_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15425" *) _09350_ : chn_out_rsci_d_125_122;
  assign _00806_ = _01679_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15411" *) _09349_ : chn_out_rsci_d_109_106;
  assign _00895_ = _01677_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15397" *) _09348_ : chn_out_rsci_d_93_90;
  assign _00885_ = _01675_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15384" *) _09347_ : chn_out_rsci_d_61_58;
  assign _00875_ = _01673_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15370" *) _09346_ : chn_out_rsci_d_29_26;
  assign _00821_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09107_ : chn_out_rsci_d_14;
  assign _00876_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09108_ : chn_out_rsci_d_30;
  assign _00881_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09109_ : chn_out_rsci_d_46;
  assign _00886_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09110_ : chn_out_rsci_d_62;
  assign _00891_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09111_ : chn_out_rsci_d_78;
  assign _00896_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09112_ : chn_out_rsci_d_94;
  assign _00807_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09113_ : chn_out_rsci_d_110;
  assign _00812_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09114_ : chn_out_rsci_d_126;
  assign _00818_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09115_ : chn_out_rsci_d_142;
  assign _00824_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09116_ : chn_out_rsci_d_158;
  assign _00831_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09117_ : chn_out_rsci_d_174;
  assign _00836_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09118_ : chn_out_rsci_d_190;
  assign _00841_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09119_ : chn_out_rsci_d_206;
  assign _00846_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09120_ : chn_out_rsci_d_222;
  assign _00851_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09121_ : chn_out_rsci_d_238;
  assign _00856_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09122_ : chn_out_rsci_d_254;
  assign _00862_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09437_ : chn_out_rsci_d_25_17;
  assign _00884_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09439_ : chn_out_rsci_d_57_49;
  assign _00894_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09441_ : chn_out_rsci_d_89_81;
  assign _00810_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09443_ : chn_out_rsci_d_121_113;
  assign _00815_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09444_ : chn_out_rsci_d_137_129;
  assign _00822_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09445_ : chn_out_rsci_d_153_145;
  assign _00828_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09446_ : chn_out_rsci_d_169_161;
  assign _00834_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09447_ : chn_out_rsci_d_185_177;
  assign _00839_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09448_ : chn_out_rsci_d_201_193;
  assign _00844_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09449_ : chn_out_rsci_d_217_209;
  assign _00849_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09450_ : chn_out_rsci_d_233_225;
  assign _00854_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09451_ : chn_out_rsci_d_249_241;
  assign _00858_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01656_ : chn_out_rsci_d_256;
  assign _00859_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01657_ : chn_out_rsci_d_257;
  assign _00860_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01658_ : chn_out_rsci_d_258;
  assign _00861_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01659_ : chn_out_rsci_d_259;
  assign _00863_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01660_ : chn_out_rsci_d_260;
  assign _00864_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01661_ : chn_out_rsci_d_261;
  assign _00865_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01662_ : chn_out_rsci_d_262;
  assign _00866_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01663_ : chn_out_rsci_d_263;
  assign _00867_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01664_ : chn_out_rsci_d_264;
  assign _00868_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01665_ : chn_out_rsci_d_265;
  assign _00869_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01666_ : chn_out_rsci_d_266;
  assign _00870_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01667_ : chn_out_rsci_d_267;
  assign _00871_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01668_ : chn_out_rsci_d_268;
  assign _00872_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01669_ : chn_out_rsci_d_269;
  assign _00873_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01670_ : chn_out_rsci_d_270;
  assign _00874_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _01671_ : chn_out_rsci_d_271;
  assign _00899_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09391_ : chn_out_rsci_d_9_1;
  assign _00879_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09438_ : chn_out_rsci_d_41_33;
  assign _00889_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09440_ : chn_out_rsci_d_73_65;
  assign _00805_ = chn_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15187" *) _09442_ : chn_out_rsci_d_105_97;
  assign _00816_ = and_3024_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15113" *) _09342_ : chn_out_rsci_d_13_10;
  assign _00880_ = and_3024_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15113" *) _09343_ : chn_out_rsci_d_45_42;
  assign _00890_ = and_3024_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15113" *) _09344_ : chn_out_rsci_d_77_74;
  assign _00817_ = and_3024_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15113" *) _09345_ : chn_out_rsci_d_141_138;
  assign _00802_ = _01655_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15102" *) chn_in_rsci_ld_core_psct_mx0c0 : chn_in_rsci_ld_core_psct;
  assign _00801_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15093" *) _04732_ : chn_in_rsci_iswt0;
  assign _00900_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:15093" *) and_dcpl_103 : chn_out_rsci_iswt0;
  assign cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl = { chn_in_rsci_d_mxwt[63], chn_in_rsci_d_mxwt[63:32] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22409" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl = { chn_in_rsci_d_mxwt[95], chn_in_rsci_d_mxwt[95:64] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22412" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl = { chn_in_rsci_d_mxwt[287], chn_in_rsci_d_mxwt[287:256] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22415" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl = { chn_in_rsci_d_mxwt[127], chn_in_rsci_d_mxwt[127:96] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22418" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl = { chn_in_rsci_d_mxwt[191], chn_in_rsci_d_mxwt[191:160] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22423" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl = { chn_in_rsci_d_mxwt[255], chn_in_rsci_d_mxwt[255:224] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22428" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl = { chn_in_rsci_d_mxwt[223], chn_in_rsci_d_mxwt[223:192] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22433" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl = { chn_in_rsci_d_mxwt[319], chn_in_rsci_d_mxwt[319:288] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22438" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl = { chn_in_rsci_d_mxwt[383], chn_in_rsci_d_mxwt[383:352] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22443" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl = { chn_in_rsci_d_mxwt[351], chn_in_rsci_d_mxwt[351:320] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22448" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl = { chn_in_rsci_d_mxwt[447], chn_in_rsci_d_mxwt[447:416] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22453" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl = { chn_in_rsci_d_mxwt[511], chn_in_rsci_d_mxwt[511:480] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22458" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl = { chn_in_rsci_d_mxwt[479], chn_in_rsci_d_mxwt[479:448] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22463" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl = { chn_in_rsci_d_mxwt[415], chn_in_rsci_d_mxwt[415:384] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22468" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl = { chn_in_rsci_d_mxwt[159], chn_in_rsci_d_mxwt[159:128] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22473" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  assign cvt_1_IntSubExt_32U_32U_33U_o_acc_nl = { chn_in_rsci_d_mxwt[31], chn_in_rsci_d_mxwt[31:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:22480" *) { cfg_offset_rsci_d[31], cfg_offset_rsci_d };
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8322" *)
  NV_NVDLA_SDP_CORE_c_core_chn_in_rsci NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_inst (
    .chn_in_rsc_lz(chn_in_rsc_lz),
    .chn_in_rsc_vz(chn_in_rsc_vz),
    .chn_in_rsc_z(chn_in_rsc_z),
    .chn_in_rsci_bawt(chn_in_rsci_bawt),
    .chn_in_rsci_d_mxwt(chn_in_rsci_d_mxwt),
    .chn_in_rsci_iswt0(chn_in_rsci_iswt0),
    .chn_in_rsci_ld_core_psct(chn_in_rsci_ld_core_psct),
    .chn_in_rsci_oswt(chn_in_rsci_oswt),
    .chn_in_rsci_wen_comp(chn_in_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8338" *)
  NV_NVDLA_SDP_CORE_c_core_chn_out_rsci NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_inst (
    .chn_out_rsc_lz(chn_out_rsc_lz),
    .chn_out_rsc_vz(chn_out_rsc_vz),
    .chn_out_rsc_z(chn_out_rsc_z),
    .chn_out_rsci_bawt(chn_out_rsci_bawt),
    .chn_out_rsci_d({ chn_out_rsci_d_271, chn_out_rsci_d_270, chn_out_rsci_d_269, chn_out_rsci_d_268, chn_out_rsci_d_267, chn_out_rsci_d_266, chn_out_rsci_d_265, chn_out_rsci_d_264, chn_out_rsci_d_263, chn_out_rsci_d_262, chn_out_rsci_d_261, chn_out_rsci_d_260, chn_out_rsci_d_259, chn_out_rsci_d_258, chn_out_rsci_d_257, chn_out_rsci_d_256, chn_out_rsci_d_255, chn_out_rsci_d_254, chn_out_rsci_d_253_250, chn_out_rsci_d_249_241, chn_out_rsci_d_240, chn_out_rsci_d_239, chn_out_rsci_d_238, chn_out_rsci_d_237_234, chn_out_rsci_d_233_225, chn_out_rsci_d_224, chn_out_rsci_d_223, chn_out_rsci_d_222, chn_out_rsci_d_221_218, chn_out_rsci_d_217_209, chn_out_rsci_d_208, chn_out_rsci_d_207, chn_out_rsci_d_206, chn_out_rsci_d_205_202, chn_out_rsci_d_201_193, chn_out_rsci_d_192, chn_out_rsci_d_191, chn_out_rsci_d_190, chn_out_rsci_d_189_186, chn_out_rsci_d_185_177, chn_out_rsci_d_176, chn_out_rsci_d_175, chn_out_rsci_d_174, chn_out_rsci_d_173_170, chn_out_rsci_d_169_161, chn_out_rsci_d_160, chn_out_rsci_d_159, chn_out_rsci_d_158, chn_out_rsci_d_157_154, chn_out_rsci_d_153_145, chn_out_rsci_d_144, chn_out_rsci_d_143, chn_out_rsci_d_142, chn_out_rsci_d_141_138, chn_out_rsci_d_137_129, chn_out_rsci_d_128, chn_out_rsci_d_127, chn_out_rsci_d_126, chn_out_rsci_d_125_122, chn_out_rsci_d_121_113, chn_out_rsci_d_112, chn_out_rsci_d_111, chn_out_rsci_d_110, chn_out_rsci_d_109_106, chn_out_rsci_d_105_97, chn_out_rsci_d_96, chn_out_rsci_d_95, chn_out_rsci_d_94, chn_out_rsci_d_93_90, chn_out_rsci_d_89_81, chn_out_rsci_d_80, chn_out_rsci_d_79, chn_out_rsci_d_78, chn_out_rsci_d_77_74, chn_out_rsci_d_73_65, chn_out_rsci_d_64, chn_out_rsci_d_63, chn_out_rsci_d_62, chn_out_rsci_d_61_58, chn_out_rsci_d_57_49, chn_out_rsci_d_48, chn_out_rsci_d_47, chn_out_rsci_d_46, chn_out_rsci_d_45_42, chn_out_rsci_d_41_33, chn_out_rsci_d_32, chn_out_rsci_d_31, chn_out_rsci_d_30, chn_out_rsci_d_29_26, chn_out_rsci_d_25_17, chn_out_rsci_d_16, chn_out_rsci_d_15, chn_out_rsci_d_14, chn_out_rsci_d_13_10, chn_out_rsci_d_9_1, chn_out_rsci_d_0 }),
    .chn_out_rsci_iswt0(chn_out_rsci_iswt0),
    .chn_out_rsci_ld_core_psct(reg_chn_out_rsci_ld_core_psct_cse),
    .chn_out_rsci_oswt(chn_out_rsci_oswt),
    .chn_out_rsci_wen_comp(chn_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8362" *)
  NV_NVDLA_SDP_CORE_c_core_core_fsm NV_NVDLA_SDP_CORE_c_core_core_fsm_inst (
    .core_wen(core_wen),
    .fsm_output(fsm_output),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8354" *)
  NV_NVDLA_SDP_CORE_c_core_staller NV_NVDLA_SDP_CORE_c_core_staller_inst (
    .chn_in_rsci_wen_comp(chn_in_rsci_wen_comp),
    .chn_out_rsci_wen_comp(chn_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7312" *)
  \$paramod\SDP_C_mgc_in_wire_v1\rscid=7\width=1  cfg_mode_eql_rsci (
    .d(cfg_mode_eql_rsci_d),
    .z(cfg_mode_eql_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7287" *)
  \$paramod\SDP_C_mgc_in_wire_v1\rscid=2\width=32  cfg_offset_rsci (
    .d(cfg_offset_rsci_d),
    .z(cfg_offset_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7307" *)
  \$paramod\SDP_C_mgc_in_wire_v1\rscid=6\width=2  cfg_out_precision_rsci (
    .d(cfg_out_precision_rsci_d),
    .z(cfg_out_precision_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7302" *)
  \$paramod\SDP_C_mgc_in_wire_v1\rscid=5\width=2  cfg_proc_precision_rsci (
    .d(cfg_proc_precision_rsci_d),
    .z(cfg_proc_precision_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7292" *)
  \$paramod\SDP_C_mgc_in_wire_v1\rscid=3\width=16  cfg_scale_rsci (
    .d(cfg_scale_rsci_d),
    .z(cfg_scale_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7297" *)
  \$paramod\SDP_C_mgc_in_wire_v1\rscid=4\width=6  cfg_truncate_rsci (
    .d(cfg_truncate_rsci_d),
    .z(cfg_truncate_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7824" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
    .a({ cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25),
    .z(cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8148" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg (
    .a(1'b1),
    .s(nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8140" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
    .a({ 1'b1, chn_idata_data_sva_1_315_287_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2, nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] }),
    .z(cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8157" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_10_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7349" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_10_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
    .a(IntMulExt_33U_16U_49U_return_10_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7501" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_10_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
    .a({ IntMulExt_33U_16U_49U_return_10_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7653" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2, nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7832" *)
  SDP_C_leading_sign_17_0 cvt_10_leading_sign_17_0_2_rg (
    .mantissa({ cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7836" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
    .a({ cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26),
    .z(cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8174" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg (
    .a(1'b1),
    .s(nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8166" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
    .a({ 1'b1, chn_idata_data_sva_1_347_319_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2, nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] }),
    .z(cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8183" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_11_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7365" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_11_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
    .a(IntMulExt_33U_16U_49U_return_11_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7517" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_11_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
    .a({ IntMulExt_33U_16U_49U_return_11_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7662" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2, nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7844" *)
  SDP_C_leading_sign_17_0 cvt_11_leading_sign_17_0_2_rg (
    .mantissa({ cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7848" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
    .a({ cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27),
    .z(cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8200" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg (
    .a(1'b1),
    .s(nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8192" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
    .a({ 1'b1, chn_idata_data_sva_1_379_351_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2, nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] }),
    .z(cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8209" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_12_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7357" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_12_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
    .a(IntMulExt_33U_16U_49U_return_12_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7509" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_12_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
    .a({ IntMulExt_33U_16U_49U_return_12_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7671" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2, nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7856" *)
  SDP_C_leading_sign_17_0 cvt_12_leading_sign_17_0_3_rg (
    .mantissa({ cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7860" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
    .a({ cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28),
    .z(cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8226" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg (
    .a(1'b1),
    .s(nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8218" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
    .a({ 1'b1, chn_idata_data_sva_1_411_383_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2, nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] }),
    .z(cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8235" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_13_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7397" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_13_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
    .a(IntMulExt_33U_16U_49U_return_13_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7549" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_13_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
    .a({ IntMulExt_33U_16U_49U_return_13_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7680" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2, nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7868" *)
  SDP_C_leading_sign_17_0 cvt_13_leading_sign_17_0_2_rg (
    .mantissa({ cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7872" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
    .a({ cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29),
    .z(cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8252" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg (
    .a(1'b1),
    .s(nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8244" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
    .a({ 1'b1, chn_idata_data_sva_1_443_415_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2, nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] }),
    .z(cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8261" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_14_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7373" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_14_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
    .a(IntMulExt_33U_16U_49U_return_14_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7525" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_14_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
    .a({ IntMulExt_33U_16U_49U_return_14_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7689" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2, nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7880" *)
  SDP_C_leading_sign_17_0 cvt_14_leading_sign_17_0_3_rg (
    .mantissa({ cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7884" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
    .a({ cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30),
    .z(cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8278" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg (
    .a(1'b1),
    .s(nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8270" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
    .a({ 1'b1, chn_idata_data_sva_1_475_447_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2, nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] }),
    .z(cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8287" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_15_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7389" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_15_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
    .a(IntMulExt_33U_16U_49U_return_15_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7541" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_15_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
    .a({ IntMulExt_33U_16U_49U_return_15_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7698" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2, nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7892" *)
  SDP_C_leading_sign_17_0 cvt_15_leading_sign_17_0_3_rg (
    .mantissa({ cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7896" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_rg (
    .a({ cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31),
    .z(cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8304" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg (
    .a(1'b1),
    .s(nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8296" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg (
    .a({ 1'b1, chn_idata_data_sva_1_507_479_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2, nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_s[0] }),
    .z(cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8313" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_16_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_4_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7381" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_16_IntShiftRightSat_49U_6U_17U_i_rshift_4_rg (
    .a(IntMulExt_33U_16U_49U_return_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7533" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_16_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_4_rg (
    .a({ IntMulExt_33U_16U_49U_return_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7707" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9, 31'b0000000000000000000000000000000 }),
    .s({ cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2, nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7904" *)
  SDP_C_leading_sign_17_0 cvt_16_leading_sign_17_0_4_rg (
    .mantissa({ cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7716" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_1_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_rg (
    .a({ cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5, FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16),
    .z(FpIntToFloat_17U_5U_10U_else_int_mant_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7916" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg (
    .a(1'b1),
    .s(nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7908" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg (
    .a({ 1'b1, chn_idata_data_sva_1_27_0_1[22:0] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2, nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[0] }),
    .z(cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7924" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_1_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7405" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_1_IntShiftRightSat_49U_6U_17U_i_rshift_rg (
    .a(IntMulExt_33U_16U_49U_return_1_sva_2),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7565" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_1_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_rg (
    .a({ IntMulExt_33U_16U_49U_return_1_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7573" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2, nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7724" *)
  SDP_C_leading_sign_17_0 cvt_1_leading_sign_17_0_rg (
    .mantissa({ cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5, FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7728" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_2_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
    .a({ cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17),
    .z(FpIntToFloat_17U_5U_10U_else_int_mant_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7940" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg (
    .a(1'b1),
    .s(nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7932" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
    .a({ 1'b1, chn_idata_data_sva_1_59_31_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2, nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] }),
    .z(cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7949" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_2_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7413" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_2_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
    .a(IntMulExt_33U_16U_49U_return_2_sva_2),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7445" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_2_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
    .a({ IntMulExt_33U_16U_49U_return_2_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7581" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2, nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7736" *)
  SDP_C_leading_sign_17_0 cvt_2_leading_sign_17_0_1_rg (
    .mantissa({ cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7740" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
    .a({ cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18),
    .z(cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7966" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg (
    .a(1'b1),
    .s(nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7958" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
    .a({ 1'b1, chn_idata_data_sva_1_91_63_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2, nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] }),
    .z(cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7975" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_3_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7421" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_3_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
    .a(IntMulExt_33U_16U_49U_return_3_sva_2),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7461" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_3_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
    .a({ IntMulExt_33U_16U_49U_return_3_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7590" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2, nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7748" *)
  SDP_C_leading_sign_17_0 cvt_3_leading_sign_17_0_1_rg (
    .mantissa({ cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7752" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
    .a({ cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19),
    .z(cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7992" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg (
    .a(1'b1),
    .s(nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7984" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
    .a({ 1'b1, chn_idata_data_sva_1_123_95_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2, nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] }),
    .z(cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8001" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_4_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7317" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_4_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
    .a(IntMulExt_33U_16U_49U_return_4_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7453" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_4_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
    .a({ IntMulExt_33U_16U_49U_return_4_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7599" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2, nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7760" *)
  SDP_C_leading_sign_17_0 cvt_4_leading_sign_17_0_2_rg (
    .mantissa({ cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7764" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
    .a({ cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20),
    .z(cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8018" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg (
    .a(1'b1),
    .s(nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8010" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
    .a({ 1'b1, chn_idata_data_sva_1_155_127_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2, nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] }),
    .z(cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8027" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_5_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7429" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_5_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
    .a(IntMulExt_33U_16U_49U_return_5_sva_2),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7493" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_5_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
    .a({ IntMulExt_33U_16U_49U_return_5_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7608" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2, nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7772" *)
  SDP_C_leading_sign_17_0 cvt_5_leading_sign_17_0_1_rg (
    .mantissa({ cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7776" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
    .a({ cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21),
    .z(cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8044" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg (
    .a(1'b1),
    .s(nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8036" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
    .a({ 1'b1, chn_idata_data_sva_1_187_159_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2, nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] }),
    .z(cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8053" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_6_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7325" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_6_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
    .a(IntMulExt_33U_16U_49U_return_6_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7469" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_6_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
    .a({ IntMulExt_33U_16U_49U_return_6_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7617" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2, nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7784" *)
  SDP_C_leading_sign_17_0 cvt_6_leading_sign_17_0_2_rg (
    .mantissa({ cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7788" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
    .a({ cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22),
    .z(cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8070" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg (
    .a(1'b1),
    .s(nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8062" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
    .a({ 1'b1, chn_idata_data_sva_1_219_191_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2, nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[0] }),
    .z(cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8079" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_7_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7341" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_7_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
    .a(IntMulExt_33U_16U_49U_return_7_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7485" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_7_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
    .a({ IntMulExt_33U_16U_49U_return_7_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7626" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2, nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7796" *)
  SDP_C_leading_sign_17_0 cvt_7_leading_sign_17_0_2_rg (
    .mantissa({ cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7800" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
    .a({ cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23),
    .z(cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8096" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg (
    .a(1'b1),
    .s(nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8088" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
    .a({ 1'b1, chn_idata_data_sva_1_251_223_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2, nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[0] }),
    .z(cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8105" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_8_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7333" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_8_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
    .a(IntMulExt_33U_16U_49U_return_8_sva_1),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7477" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_8_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
    .a({ IntMulExt_33U_16U_49U_return_8_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7635" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2, nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7808" *)
  SDP_C_leading_sign_17_0 cvt_8_leading_sign_17_0_3_rg (
    .mantissa({ cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7812" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=17\signd_a=0\width_s=5\width_z=17  cvt_9_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
    .a({ cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 }),
    .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24),
    .z(FpIntToFloat_17U_5U_10U_else_int_mant_9_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8122" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg (
    .a(1'b1),
    .s(nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
    .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8114" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=24\signd_a=0\width_s=4\width_z=24  cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
    .a({ 1'b1, chn_idata_data_sva_1_283_255_1[23:1] }),
    .s({ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2, nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[0] }),
    .z(cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:8131" *)
  \$paramod\SDP_C_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=5\width_z=24  cvt_9_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg (
    .a(1'b1),
    .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2),
    .z(FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7437" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=49\signd_a=1\width_s=6\width_z=49  cvt_9_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
    .a(IntMulExt_33U_16U_49U_return_9_sva_2),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7557" *)
  \$paramod\SDP_C_mgc_shift_r_v4\width_a=112\signd_a=1\width_s=6\width_z=112  cvt_9_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
    .a({ IntMulExt_33U_16U_49U_return_9_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_2),
    .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7644" *)
  \$paramod\SDP_C_mgc_shift_br_v4\width_a=42\signd_a=0\width_s=6\width_z=75  cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg (
    .a({ 1'b1, FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8, 31'b0000000000000000000000000000000 }),
    .s({ cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2, nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[0] }),
    .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:7820" *)
  SDP_C_leading_sign_17_0 cvt_9_leading_sign_17_0_1_rg (
    .mantissa({ cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 }),
    .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24)
  );
  assign _00000_[2] = and_1179_nl;
  assign _00002_[2:1] = { FpIntToFloat_17U_5U_10U_o_expo_or_15_nl, FpIntToFloat_17U_5U_10U_o_expo_and_31_nl };
  assign _00171_[9] = _00171_[10];
  assign _00172_[9] = _00172_[10];
  assign _00173_[9] = _00173_[10];
  assign _00174_[9] = _00174_[10];
  assign _00175_[9] = _00175_[10];
  assign _00176_[9] = _00176_[10];
  assign _00177_[9] = _00177_[10];
  assign _00178_[9] = _00178_[10];
  assign _00179_[9] = _00179_[10];
  assign _00180_[9] = _00180_[10];
  assign _00181_[9] = _00181_[10];
  assign _00182_[9] = _00182_[10];
  assign _00183_[9] = _00183_[10];
  assign _00184_[9] = _00184_[10];
  assign _00185_[9] = _00185_[10];
  assign _00186_[9] = _00186_[10];
  assign _00187_[1] = _00187_[2];
  assign _00188_[1] = _00188_[2];
  assign _00189_[1] = _00189_[2];
  assign _00190_[2:1] = { or_dcpl_109, or_dcpl_109 };
  assign _00191_[2:1] = { or_dcpl_111, or_dcpl_111 };
  assign _00192_[2:1] = { or_dcpl_114, or_dcpl_114 };
  assign _00193_[2:1] = { or_dcpl_116, or_dcpl_116 };
  assign _00194_[2:1] = { or_dcpl_120, or_dcpl_120 };
  assign _00195_[1] = _00195_[2];
  assign _00196_[2:1] = { or_dcpl_125, or_dcpl_125 };
  assign _00197_[2:1] = { or_dcpl_127, or_dcpl_127 };
  assign _00198_[2:1] = { or_dcpl_131, or_dcpl_131 };
  assign _00199_[2:1] = { or_dcpl_133, or_dcpl_133 };
  assign _00200_[2:1] = { or_dcpl_137, or_dcpl_137 };
  assign _00201_[2:1] = { or_dcpl_140, or_dcpl_140 };
  assign _00202_[2:1] = { or_dcpl_144, or_dcpl_144 };
  assign _00235_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  assign _00236_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  assign _00237_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  assign _00238_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0;
  assign _00239_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0;
  assign _00240_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0;
  assign _00241_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0;
  assign _00242_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0;
  assign _00243_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0;
  assign _00244_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0;
  assign _00245_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0;
  assign _00246_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0;
  assign _00247_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0;
  assign _00248_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0;
  assign _00249_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0;
  assign _00250_[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  assign _03846_[1:0] = _03521_;
  assign _03864_[8:0] = cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  assign FpFloatToInt_16U_5U_10U_shift_and_8_cse = FpFloatToInt_16U_5U_10U_shift_and_5_cse;
  assign and_1038_cse = and_1023_nl;
  assign and_976_cse = and_1013_nl;
  assign chn_in_rsci_oswt_unreg = or_tmp_3487;
  assign chn_out_rsci_oswt_unreg = and_dcpl_73;
  assign cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign cvt_10_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1 = cvt_10_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign cvt_10_IntSaturation_17U_8U_else_if_acc_2_itm_10 = cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign cvt_11_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1 = cvt_11_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign cvt_11_IntSaturation_17U_8U_else_if_acc_2_itm_10 = cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign cvt_12_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1 = cvt_12_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign cvt_12_IntSaturation_17U_8U_else_if_acc_3_itm_10 = cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign cvt_13_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1 = cvt_13_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign cvt_13_IntSaturation_17U_8U_else_if_acc_2_itm_10 = cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign cvt_14_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1 = cvt_14_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign cvt_14_IntSaturation_17U_8U_else_if_acc_3_itm_10 = cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign cvt_15_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1 = cvt_15_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign cvt_15_IntSaturation_17U_8U_else_if_acc_3_itm_10 = cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1 = cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11];
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4 = cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl[4];
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1 = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl[8];
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1 = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8];
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1 = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7];
  assign cvt_16_IntSaturation_17U_16U_else_if_acc_4_itm_2_1 = cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl[2];
  assign cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1 = cvt_16_IntSaturation_17U_16U_if_acc_4_nl[2];
  assign cvt_16_IntSaturation_17U_8U_else_if_acc_4_itm_10 = cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl[10];
  assign cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1 = cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl[11];
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4 = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl[4];
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1 = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8];
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1 = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8];
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7];
  assign cvt_1_IntSaturation_17U_16U_else_if_acc_itm_2_1 = cvt_1_IntSaturation_17U_16U_else_if_acc_nl[2];
  assign cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1 = cvt_1_IntSaturation_17U_16U_if_acc_nl[2];
  assign cvt_1_IntSaturation_17U_8U_else_if_acc_itm_10 = cvt_1_IntSaturation_17U_8U_else_if_acc_nl[10];
  assign cvt_1_IntSaturation_17U_8U_if_acc_itm_10_1 = cvt_1_IntSaturation_17U_8U_if_acc_nl[10];
  assign cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign cvt_2_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1 = cvt_2_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign cvt_2_IntSaturation_17U_8U_else_if_acc_1_itm_10 = cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1 = and_550_cse;
  assign cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign cvt_3_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1 = cvt_3_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign cvt_3_IntSaturation_17U_8U_else_if_acc_1_itm_10 = cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign cvt_3_IntSaturation_17U_8U_if_acc_1_itm_10_1 = cvt_3_IntSaturation_17U_8U_if_acc_1_nl[10];
  assign cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign cvt_4_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1 = cvt_4_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign cvt_4_IntSaturation_17U_8U_else_if_acc_2_itm_10 = cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign cvt_5_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1 = cvt_5_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign cvt_5_IntSaturation_17U_8U_else_if_acc_1_itm_10 = cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign cvt_5_IntSaturation_17U_8U_if_acc_1_itm_10_1 = cvt_5_IntSaturation_17U_8U_if_acc_1_nl[10];
  assign cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign cvt_6_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1 = cvt_6_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign cvt_6_IntSaturation_17U_8U_else_if_acc_2_itm_10 = cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11];
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4];
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8];
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8];
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7];
  assign cvt_7_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl[2];
  assign cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1 = cvt_7_IntSaturation_17U_16U_if_acc_2_nl[2];
  assign cvt_7_IntSaturation_17U_8U_else_if_acc_2_itm_10 = cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl[10];
  assign cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11];
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4];
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8];
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8];
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7];
  assign cvt_8_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl[2];
  assign cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1 = cvt_8_IntSaturation_17U_16U_if_acc_3_nl[2];
  assign cvt_8_IntSaturation_17U_8U_else_if_acc_3_itm_10 = cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl[10];
  assign cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11];
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4];
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8];
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8];
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7];
  assign cvt_9_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl[2];
  assign cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1 = cvt_9_IntSaturation_17U_16U_if_acc_1_nl[2];
  assign cvt_9_IntSaturation_17U_8U_else_if_acc_1_itm_10 = cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl[10];
  assign cvt_9_IntSaturation_17U_8U_if_acc_1_itm_10_1 = cvt_9_IntSaturation_17U_8U_if_acc_1_nl[10];
  assign cvt_else_equal_tmp_45_mx1 = cvt_else_equal_tmp_39_mx1;
  assign cvt_else_equal_tmp_46_mx1 = cvt_else_equal_tmp_40_mx1;
  assign cvt_else_nor_dfs_15_mx1 = cvt_else_nor_dfs_13_mx1;
  assign mux_1046_nl = mux_tmp_1047;
  assign mux_1108_nl = mux_tmp_1109;
  assign mux_1281_nl = mux_tmp_1280;
  assign mux_1338_nl = mux_tmp_1337;
  assign mux_1340_nl = mux_tmp_1337;
  assign mux_175_nl = mux_169_nl;
  assign mux_1772_nl = mux_1762_cse;
  assign mux_1785_nl = mux_1780_nl;
  assign mux_2172_nl = mux_2183_nl;
  assign mux_2173_nl = mux_2185_nl;
  assign mux_2174_nl = mux_2186_nl;
  assign mux_2216_nl = mux_2215_nl;
  assign mux_2221_nl = mux_2219_nl;
  assign mux_919_nl = mux_1832_nl;
  assign mux_tmp_1282 = mux_tmp_1280;
  assign mux_tmp_1339 = mux_tmp_1337;
  assign mux_tmp_1341 = mux_tmp_1337;
  assign mux_tmp_2206 = mux_2208_nl;
  assign nand_tmp_30 = mux_tmp_1047;
  assign nand_tmp_36 = mux_tmp_1109;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva;
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva[15:0] = FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva;
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[16:0] = FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva;
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10:0] = FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0;
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0[2:0] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva;
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[44:0] = IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva;
  assign nl_NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_inst_chn_out_rsci_d = { chn_out_rsci_d_271, chn_out_rsci_d_270, chn_out_rsci_d_269, chn_out_rsci_d_268, chn_out_rsci_d_267, chn_out_rsci_d_266, chn_out_rsci_d_265, chn_out_rsci_d_264, chn_out_rsci_d_263, chn_out_rsci_d_262, chn_out_rsci_d_261, chn_out_rsci_d_260, chn_out_rsci_d_259, chn_out_rsci_d_258, chn_out_rsci_d_257, chn_out_rsci_d_256, chn_out_rsci_d_255, chn_out_rsci_d_254, chn_out_rsci_d_253_250, chn_out_rsci_d_249_241, chn_out_rsci_d_240, chn_out_rsci_d_239, chn_out_rsci_d_238, chn_out_rsci_d_237_234, chn_out_rsci_d_233_225, chn_out_rsci_d_224, chn_out_rsci_d_223, chn_out_rsci_d_222, chn_out_rsci_d_221_218, chn_out_rsci_d_217_209, chn_out_rsci_d_208, chn_out_rsci_d_207, chn_out_rsci_d_206, chn_out_rsci_d_205_202, chn_out_rsci_d_201_193, chn_out_rsci_d_192, chn_out_rsci_d_191, chn_out_rsci_d_190, chn_out_rsci_d_189_186, chn_out_rsci_d_185_177, chn_out_rsci_d_176, chn_out_rsci_d_175, chn_out_rsci_d_174, chn_out_rsci_d_173_170, chn_out_rsci_d_169_161, chn_out_rsci_d_160, chn_out_rsci_d_159, chn_out_rsci_d_158, chn_out_rsci_d_157_154, chn_out_rsci_d_153_145, chn_out_rsci_d_144, chn_out_rsci_d_143, chn_out_rsci_d_142, chn_out_rsci_d_141_138, chn_out_rsci_d_137_129, chn_out_rsci_d_128, chn_out_rsci_d_127, chn_out_rsci_d_126, chn_out_rsci_d_125_122, chn_out_rsci_d_121_113, chn_out_rsci_d_112, chn_out_rsci_d_111, chn_out_rsci_d_110, chn_out_rsci_d_109_106, chn_out_rsci_d_105_97, chn_out_rsci_d_96, chn_out_rsci_d_95, chn_out_rsci_d_94, chn_out_rsci_d_93_90, chn_out_rsci_d_89_81, chn_out_rsci_d_80, chn_out_rsci_d_79, chn_out_rsci_d_78, chn_out_rsci_d_77_74, chn_out_rsci_d_73_65, chn_out_rsci_d_64, chn_out_rsci_d_63, chn_out_rsci_d_62, chn_out_rsci_d_61_58, chn_out_rsci_d_57_49, chn_out_rsci_d_48, chn_out_rsci_d_47, chn_out_rsci_d_46, chn_out_rsci_d_45_42, chn_out_rsci_d_41_33, chn_out_rsci_d_32, chn_out_rsci_d_31, chn_out_rsci_d_30, chn_out_rsci_d_29_26, chn_out_rsci_d_25_17, chn_out_rsci_d_16, chn_out_rsci_d_15, chn_out_rsci_d_14, chn_out_rsci_d_13_10, chn_out_rsci_d_9_1, chn_out_rsci_d_0 };
  assign nl_cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0] = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  assign nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0] = cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  assign nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0] = cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  assign nl_cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = { cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 };
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = chn_idata_data_sva_1_315_287_1[23:1];
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2;
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0] = cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign nl_cvt_10_FpMantRNE_17U_11U_else_acc_2_nl[9:0] = cvt_10_FpMantRNE_17U_11U_else_acc_2_nl;
  assign nl_cvt_10_FpMantRNE_24U_11U_else_acc_2_nl[9:0] = cvt_10_FpMantRNE_24U_11U_else_acc_2_nl;
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0] = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0] = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0] = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0] = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  assign nl_cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl[2:0] = cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl;
  assign nl_cvt_10_IntSaturation_17U_16U_if_acc_2_nl[2:0] = cvt_10_IntSaturation_17U_16U_if_acc_2_nl;
  assign nl_cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl[10:0] = cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl;
  assign nl_cvt_10_IntSaturation_17U_8U_if_acc_2_nl[10:0] = cvt_10_IntSaturation_17U_8U_if_acc_2_nl;
  assign nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0] = cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  assign nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0] = cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  assign nl_cvt_10_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = { IntMulExt_33U_16U_49U_return_10_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0] = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  assign nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:1] = cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign nl_cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0] = cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl;
  assign nl_cvt_10_leading_sign_17_0_2_rg_mantissa = { cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 };
  assign nl_cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0] = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  assign nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0] = cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  assign nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0] = cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  assign nl_cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = { cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 };
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = chn_idata_data_sva_1_347_319_1[23:1];
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2;
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0] = cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign nl_cvt_11_FpMantRNE_17U_11U_else_acc_2_nl[9:0] = cvt_11_FpMantRNE_17U_11U_else_acc_2_nl;
  assign nl_cvt_11_FpMantRNE_24U_11U_else_acc_2_nl[9:0] = cvt_11_FpMantRNE_24U_11U_else_acc_2_nl;
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0] = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0] = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0] = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0] = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  assign nl_cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl[2:0] = cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl;
  assign nl_cvt_11_IntSaturation_17U_16U_if_acc_2_nl[2:0] = cvt_11_IntSaturation_17U_16U_if_acc_2_nl;
  assign nl_cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl[10:0] = cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl;
  assign nl_cvt_11_IntSaturation_17U_8U_if_acc_2_nl[10:0] = cvt_11_IntSaturation_17U_8U_if_acc_2_nl;
  assign nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0] = cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  assign nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0] = cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  assign nl_cvt_11_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = { IntMulExt_33U_16U_49U_return_11_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0] = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  assign nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:1] = cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign nl_cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0] = cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl;
  assign nl_cvt_11_leading_sign_17_0_2_rg_mantissa = { cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 };
  assign nl_cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0] = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  assign nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0] = cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  assign nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0] = cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  assign nl_cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = { cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 };
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = chn_idata_data_sva_1_379_351_1[23:1];
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2;
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0] = cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign nl_cvt_12_FpMantRNE_17U_11U_else_acc_3_nl[9:0] = cvt_12_FpMantRNE_17U_11U_else_acc_3_nl;
  assign nl_cvt_12_FpMantRNE_24U_11U_else_acc_3_nl[9:0] = cvt_12_FpMantRNE_24U_11U_else_acc_3_nl;
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0] = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0] = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0] = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0] = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  assign nl_cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl[2:0] = cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl;
  assign nl_cvt_12_IntSaturation_17U_16U_if_acc_3_nl[2:0] = cvt_12_IntSaturation_17U_16U_if_acc_3_nl;
  assign nl_cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl[10:0] = cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl;
  assign nl_cvt_12_IntSaturation_17U_8U_if_acc_3_nl[10:0] = cvt_12_IntSaturation_17U_8U_if_acc_3_nl;
  assign nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0] = cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  assign nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17:0] = cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  assign nl_cvt_12_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = { IntMulExt_33U_16U_49U_return_12_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0] = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  assign nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:1] = cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign nl_cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0] = cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl;
  assign nl_cvt_12_leading_sign_17_0_3_rg_mantissa = { cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 };
  assign nl_cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0] = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  assign nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0] = cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  assign nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0] = cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  assign nl_cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = { cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 };
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = chn_idata_data_sva_1_411_383_1[23:1];
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2;
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0] = cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign nl_cvt_13_FpMantRNE_17U_11U_else_acc_2_nl[9:0] = cvt_13_FpMantRNE_17U_11U_else_acc_2_nl;
  assign nl_cvt_13_FpMantRNE_24U_11U_else_acc_2_nl[9:0] = cvt_13_FpMantRNE_24U_11U_else_acc_2_nl;
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0] = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0] = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0] = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0] = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  assign nl_cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl[2:0] = cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl;
  assign nl_cvt_13_IntSaturation_17U_16U_if_acc_2_nl[2:0] = cvt_13_IntSaturation_17U_16U_if_acc_2_nl;
  assign nl_cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl[10:0] = cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl;
  assign nl_cvt_13_IntSaturation_17U_8U_if_acc_2_nl[10:0] = cvt_13_IntSaturation_17U_8U_if_acc_2_nl;
  assign nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0] = cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  assign nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0] = cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  assign nl_cvt_13_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = { IntMulExt_33U_16U_49U_return_13_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0] = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  assign nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:1] = cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign nl_cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0] = cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl;
  assign nl_cvt_13_leading_sign_17_0_2_rg_mantissa = { cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 };
  assign nl_cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0] = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  assign nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0] = cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  assign nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0] = cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  assign nl_cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = { cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 };
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = chn_idata_data_sva_1_443_415_1[23:1];
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2;
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0] = cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign nl_cvt_14_FpMantRNE_17U_11U_else_acc_3_nl[9:0] = cvt_14_FpMantRNE_17U_11U_else_acc_3_nl;
  assign nl_cvt_14_FpMantRNE_24U_11U_else_acc_3_nl[9:0] = cvt_14_FpMantRNE_24U_11U_else_acc_3_nl;
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0] = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0] = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0] = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0] = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  assign nl_cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl[2:0] = cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl;
  assign nl_cvt_14_IntSaturation_17U_16U_if_acc_3_nl[2:0] = cvt_14_IntSaturation_17U_16U_if_acc_3_nl;
  assign nl_cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl[10:0] = cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl;
  assign nl_cvt_14_IntSaturation_17U_8U_if_acc_3_nl[10:0] = cvt_14_IntSaturation_17U_8U_if_acc_3_nl;
  assign nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0] = cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  assign nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[0];
  assign nl_cvt_14_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = { IntMulExt_33U_16U_49U_return_14_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0] = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  assign nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:1] = cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign nl_cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0] = cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl;
  assign nl_cvt_14_leading_sign_17_0_3_rg_mantissa = { cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 };
  assign nl_cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0] = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  assign nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0] = cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  assign nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0] = cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  assign nl_cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = { cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 };
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = chn_idata_data_sva_1_475_447_1[23:1];
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2;
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0] = cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign nl_cvt_15_FpMantRNE_17U_11U_else_acc_3_nl[9:0] = cvt_15_FpMantRNE_17U_11U_else_acc_3_nl;
  assign nl_cvt_15_FpMantRNE_24U_11U_else_acc_3_nl[9:0] = cvt_15_FpMantRNE_24U_11U_else_acc_3_nl;
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0] = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0] = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0] = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0] = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  assign nl_cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl[2:0] = cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl;
  assign nl_cvt_15_IntSaturation_17U_16U_if_acc_3_nl[2:0] = cvt_15_IntSaturation_17U_16U_if_acc_3_nl;
  assign nl_cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl[10:0] = cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl;
  assign nl_cvt_15_IntSaturation_17U_8U_if_acc_3_nl[10:0] = cvt_15_IntSaturation_17U_8U_if_acc_3_nl;
  assign nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0] = cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  assign nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17:0] = cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  assign nl_cvt_15_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = { IntMulExt_33U_16U_49U_return_15_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0] = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  assign nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:1] = cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign nl_cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0] = cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl;
  assign nl_cvt_15_leading_sign_17_0_3_rg_mantissa = { cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 };
  assign nl_cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11:0] = cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl;
  assign nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl[4:0] = cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl;
  assign nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl[4:0] = cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl;
  assign nl_cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_rg_a = { cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 };
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_a = chn_idata_data_sva_1_507_479_1[23:1];
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2;
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl[22:0] = cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl;
  assign nl_cvt_16_FpMantRNE_17U_11U_else_acc_4_nl[9:0] = cvt_16_FpMantRNE_17U_11U_else_acc_4_nl;
  assign nl_cvt_16_FpMantRNE_24U_11U_else_acc_4_nl[9:0] = cvt_16_FpMantRNE_24U_11U_else_acc_4_nl;
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl[8:0] = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl;
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8:0] = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl;
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp[4:0] = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp;
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7:0] = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl;
  assign nl_cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl[2:0] = cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl;
  assign nl_cvt_16_IntSaturation_17U_16U_if_acc_4_nl[2:0] = cvt_16_IntSaturation_17U_16U_if_acc_4_nl;
  assign nl_cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl[10:0] = cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl;
  assign nl_cvt_16_IntSaturation_17U_8U_if_acc_4_nl[10:0] = cvt_16_IntSaturation_17U_8U_if_acc_4_nl;
  assign nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17:0] = cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl;
  assign nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17:0] = cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl;
  assign nl_cvt_16_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_4_rg_a = { IntMulExt_33U_16U_49U_return_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[49:0] = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp;
  assign nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9, 31'b0000000000000000000000000000000 };
  assign nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_s[2:1] = cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2[1:0];
  assign nl_cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl[32:0] = cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl;
  assign nl_cvt_16_leading_sign_17_0_4_rg_mantissa = { cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 };
  assign nl_cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl[11:0] = cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl;
  assign nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl[4:0] = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl;
  assign nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl[4:0] = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl;
  assign nl_cvt_1_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_rg_a = { cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5, FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 };
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a = chn_idata_data_sva_1_27_0_1[22:0];
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2;
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl[22:0] = cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  assign nl_cvt_1_FpMantRNE_17U_11U_else_acc_nl[9:0] = cvt_1_FpMantRNE_17U_11U_else_acc_nl;
  assign nl_cvt_1_FpMantRNE_24U_11U_else_acc_nl[9:0] = cvt_1_FpMantRNE_24U_11U_else_acc_nl;
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8:0] = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl;
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8:0] = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl;
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp[4:0] = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp;
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7:0] = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl;
  assign nl_cvt_1_IntSaturation_17U_16U_else_if_acc_nl[2:0] = cvt_1_IntSaturation_17U_16U_else_if_acc_nl;
  assign nl_cvt_1_IntSaturation_17U_16U_if_acc_nl[2:0] = cvt_1_IntSaturation_17U_16U_if_acc_nl;
  assign nl_cvt_1_IntSaturation_17U_8U_else_if_acc_nl[10:0] = cvt_1_IntSaturation_17U_8U_else_if_acc_nl;
  assign nl_cvt_1_IntSaturation_17U_8U_if_acc_nl[10:0] = cvt_1_IntSaturation_17U_8U_if_acc_nl;
  assign nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17:0] = cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl;
  assign nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17:0] = cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl;
  assign nl_cvt_1_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_rg_a = { IntMulExt_33U_16U_49U_return_1_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[49:0] = cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp;
  assign nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_s[5:1] = cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2;
  assign nl_cvt_1_IntSubExt_32U_32U_33U_o_acc_nl[32:0] = cvt_1_IntSubExt_32U_32U_33U_o_acc_nl;
  assign nl_cvt_1_leading_sign_17_0_rg_mantissa = { cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5, FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 };
  assign nl_cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0] = cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  assign nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0] = cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  assign nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0] = cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  assign nl_cvt_2_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = { cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 };
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = chn_idata_data_sva_1_59_31_1[23:1];
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2;
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0] = cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign nl_cvt_2_FpMantRNE_17U_11U_else_acc_1_nl[9:0] = cvt_2_FpMantRNE_17U_11U_else_acc_1_nl;
  assign nl_cvt_2_FpMantRNE_24U_11U_else_acc_1_nl[9:0] = cvt_2_FpMantRNE_24U_11U_else_acc_1_nl;
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0] = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0] = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0] = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0] = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  assign nl_cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl[2:0] = cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl;
  assign nl_cvt_2_IntSaturation_17U_16U_if_acc_1_nl[2:0] = cvt_2_IntSaturation_17U_16U_if_acc_1_nl;
  assign nl_cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl[10:0] = cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl;
  assign nl_cvt_2_IntSaturation_17U_8U_if_acc_1_nl[10:0] = cvt_2_IntSaturation_17U_8U_if_acc_1_nl;
  assign nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0] = cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  assign nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0] = cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  assign nl_cvt_2_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = { IntMulExt_33U_16U_49U_return_2_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0] = cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  assign nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:1] = cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign nl_cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0] = cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl;
  assign nl_cvt_2_leading_sign_17_0_1_rg_mantissa = { cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 };
  assign nl_cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0] = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  assign nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0] = cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  assign nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0] = cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  assign nl_cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = { cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 };
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = chn_idata_data_sva_1_91_63_1[23:1];
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2;
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0] = cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign nl_cvt_3_FpMantRNE_17U_11U_else_acc_1_nl[9:0] = cvt_3_FpMantRNE_17U_11U_else_acc_1_nl;
  assign nl_cvt_3_FpMantRNE_24U_11U_else_acc_1_nl[9:0] = cvt_3_FpMantRNE_24U_11U_else_acc_1_nl;
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0] = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0] = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0] = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0] = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  assign nl_cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl[2:0] = cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl;
  assign nl_cvt_3_IntSaturation_17U_16U_if_acc_1_nl[2:0] = cvt_3_IntSaturation_17U_16U_if_acc_1_nl;
  assign nl_cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl[10:0] = cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl;
  assign nl_cvt_3_IntSaturation_17U_8U_if_acc_1_nl[10:0] = cvt_3_IntSaturation_17U_8U_if_acc_1_nl;
  assign nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0] = cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  assign nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0] = cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  assign nl_cvt_3_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = { IntMulExt_33U_16U_49U_return_3_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0] = cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  assign nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:1] = cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign nl_cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0] = cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl;
  assign nl_cvt_3_leading_sign_17_0_1_rg_mantissa = { cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 };
  assign nl_cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0] = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  assign nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0] = cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  assign nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0] = cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  assign nl_cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = { cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 };
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = chn_idata_data_sva_1_123_95_1[23:1];
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2;
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0] = cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign nl_cvt_4_FpMantRNE_17U_11U_else_acc_2_nl[9:0] = cvt_4_FpMantRNE_17U_11U_else_acc_2_nl;
  assign nl_cvt_4_FpMantRNE_24U_11U_else_acc_2_nl[9:0] = cvt_4_FpMantRNE_24U_11U_else_acc_2_nl;
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0] = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0] = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0] = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0] = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  assign nl_cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl[2:0] = cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl;
  assign nl_cvt_4_IntSaturation_17U_16U_if_acc_2_nl[2:0] = cvt_4_IntSaturation_17U_16U_if_acc_2_nl;
  assign nl_cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl[10:0] = cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl;
  assign nl_cvt_4_IntSaturation_17U_8U_if_acc_2_nl[10:0] = cvt_4_IntSaturation_17U_8U_if_acc_2_nl;
  assign nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0] = cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  assign nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0] = cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  assign nl_cvt_4_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = { IntMulExt_33U_16U_49U_return_4_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0] = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  assign nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[4:1] = cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[3:0];
  assign nl_cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0] = cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl;
  assign nl_cvt_4_leading_sign_17_0_2_rg_mantissa = { cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 };
  assign nl_cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0] = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  assign nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0] = cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  assign nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0] = cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  assign nl_cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = { cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 };
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = chn_idata_data_sva_1_155_127_1[23:1];
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2;
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0] = cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign nl_cvt_5_FpMantRNE_17U_11U_else_acc_1_nl[9:0] = cvt_5_FpMantRNE_17U_11U_else_acc_1_nl;
  assign nl_cvt_5_FpMantRNE_24U_11U_else_acc_1_nl[9:0] = cvt_5_FpMantRNE_24U_11U_else_acc_1_nl;
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0] = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0] = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0] = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0] = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  assign nl_cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl[2:0] = cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl;
  assign nl_cvt_5_IntSaturation_17U_16U_if_acc_1_nl[2:0] = cvt_5_IntSaturation_17U_16U_if_acc_1_nl;
  assign nl_cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl[10:0] = cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl;
  assign nl_cvt_5_IntSaturation_17U_8U_if_acc_1_nl[10:0] = cvt_5_IntSaturation_17U_8U_if_acc_1_nl;
  assign nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0] = cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  assign nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0] = cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  assign nl_cvt_5_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = { IntMulExt_33U_16U_49U_return_5_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0] = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  assign nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:1] = cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign nl_cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0] = cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl;
  assign nl_cvt_5_leading_sign_17_0_1_rg_mantissa = { cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 };
  assign nl_cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0] = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  assign nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0] = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  assign nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0] = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  assign nl_cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = { cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 };
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = chn_idata_data_sva_1_187_159_1[23:1];
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2;
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0] = cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign nl_cvt_6_FpMantRNE_17U_11U_else_acc_2_nl[9:0] = cvt_6_FpMantRNE_17U_11U_else_acc_2_nl;
  assign nl_cvt_6_FpMantRNE_24U_11U_else_acc_2_nl[9:0] = cvt_6_FpMantRNE_24U_11U_else_acc_2_nl;
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0] = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0] = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0] = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0] = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  assign nl_cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl[2:0] = cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl;
  assign nl_cvt_6_IntSaturation_17U_16U_if_acc_2_nl[2:0] = cvt_6_IntSaturation_17U_16U_if_acc_2_nl;
  assign nl_cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl[10:0] = cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl;
  assign nl_cvt_6_IntSaturation_17U_8U_if_acc_2_nl[10:0] = cvt_6_IntSaturation_17U_8U_if_acc_2_nl;
  assign nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0] = cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  assign nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0] = cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  assign nl_cvt_6_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = { IntMulExt_33U_16U_49U_return_6_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0] = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  assign nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:1] = cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign nl_cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0] = cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl;
  assign nl_cvt_6_leading_sign_17_0_2_rg_mantissa = { cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 };
  assign nl_cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0] = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  assign nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0] = cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  assign nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0] = cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  assign nl_cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = { cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 };
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = chn_idata_data_sva_1_219_191_1[23:1];
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2;
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0] = cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  assign nl_cvt_7_FpMantRNE_17U_11U_else_acc_2_nl[9:0] = cvt_7_FpMantRNE_17U_11U_else_acc_2_nl;
  assign nl_cvt_7_FpMantRNE_24U_11U_else_acc_2_nl[9:0] = cvt_7_FpMantRNE_24U_11U_else_acc_2_nl;
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0] = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0] = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0] = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0] = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  assign nl_cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl[2:0] = cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl;
  assign nl_cvt_7_IntSaturation_17U_16U_if_acc_2_nl[2:0] = cvt_7_IntSaturation_17U_16U_if_acc_2_nl;
  assign nl_cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl[10:0] = cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl;
  assign nl_cvt_7_IntSaturation_17U_8U_if_acc_2_nl[10:0] = cvt_7_IntSaturation_17U_8U_if_acc_2_nl;
  assign nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0] = cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  assign nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0] = cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  assign nl_cvt_7_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = { IntMulExt_33U_16U_49U_return_7_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0] = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  assign nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:1] = cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  assign nl_cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0] = cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl;
  assign nl_cvt_7_leading_sign_17_0_2_rg_mantissa = { cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 };
  assign nl_cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0] = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  assign nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0] = cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  assign nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0] = cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  assign nl_cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = { cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 };
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = chn_idata_data_sva_1_251_223_1[23:1];
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2;
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0] = cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  assign nl_cvt_8_FpMantRNE_17U_11U_else_acc_3_nl[9:0] = cvt_8_FpMantRNE_17U_11U_else_acc_3_nl;
  assign nl_cvt_8_FpMantRNE_24U_11U_else_acc_3_nl[9:0] = cvt_8_FpMantRNE_24U_11U_else_acc_3_nl;
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0] = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0] = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0] = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0] = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  assign nl_cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl[2:0] = cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl;
  assign nl_cvt_8_IntSaturation_17U_16U_if_acc_3_nl[2:0] = cvt_8_IntSaturation_17U_16U_if_acc_3_nl;
  assign nl_cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl[10:0] = cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl;
  assign nl_cvt_8_IntSaturation_17U_8U_if_acc_3_nl[10:0] = cvt_8_IntSaturation_17U_8U_if_acc_3_nl;
  assign nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0] = cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  assign nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17:0] = cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  assign nl_cvt_8_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = { IntMulExt_33U_16U_49U_return_8_sva_1, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0] = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  assign nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:1] = cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  assign nl_cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0] = cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl;
  assign nl_cvt_8_leading_sign_17_0_3_rg_mantissa = { cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg, reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg, FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 };
  assign nl_cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0] = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  assign nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0] = cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  assign nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0] = cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  assign nl_cvt_9_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = { cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 };
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = chn_idata_data_sva_1_283_255_1[23:1];
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:1] = FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2;
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0] = cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  assign nl_cvt_9_FpMantRNE_17U_11U_else_acc_1_nl[9:0] = cvt_9_FpMantRNE_17U_11U_else_acc_1_nl;
  assign nl_cvt_9_FpMantRNE_24U_11U_else_acc_1_nl[9:0] = cvt_9_FpMantRNE_24U_11U_else_acc_1_nl;
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0] = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0] = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0] = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0] = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  assign nl_cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl[2:0] = cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl;
  assign nl_cvt_9_IntSaturation_17U_16U_if_acc_1_nl[2:0] = cvt_9_IntSaturation_17U_16U_if_acc_1_nl;
  assign nl_cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl[10:0] = cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl;
  assign nl_cvt_9_IntSaturation_17U_8U_if_acc_1_nl[10:0] = cvt_9_IntSaturation_17U_8U_if_acc_1_nl;
  assign nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0] = cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  assign nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0] = cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  assign nl_cvt_9_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = { IntMulExt_33U_16U_49U_return_9_sva_2, 63'b000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0] = cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  assign nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = { FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8, 31'b0000000000000000000000000000000 };
  assign nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:1] = cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  assign nl_cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0] = cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl;
  assign nl_cvt_9_leading_sign_17_0_1_rg_mantissa = { cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16, FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6, FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 };
  assign oWidth_aWidth_bWidth_prb = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_1 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_10 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_11 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_12 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_13 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_14 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_15 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_2 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_3 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_4 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_5 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_6 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_7 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_8 = and_550_cse;
  assign oWidth_aWidth_bWidth_prb_9 = and_550_cse;
  assign oWidth_mWidth_prb = and_550_cse;
  assign oWidth_mWidth_prb_1 = and_550_cse;
  assign oWidth_mWidth_prb_10 = and_550_cse;
  assign oWidth_mWidth_prb_11 = and_550_cse;
  assign oWidth_mWidth_prb_12 = and_550_cse;
  assign oWidth_mWidth_prb_13 = and_550_cse;
  assign oWidth_mWidth_prb_14 = and_550_cse;
  assign oWidth_mWidth_prb_15 = and_550_cse;
  assign oWidth_mWidth_prb_2 = and_550_cse;
  assign oWidth_mWidth_prb_3 = and_550_cse;
  assign oWidth_mWidth_prb_4 = and_550_cse;
  assign oWidth_mWidth_prb_5 = and_550_cse;
  assign oWidth_mWidth_prb_6 = and_550_cse;
  assign oWidth_mWidth_prb_7 = and_550_cse;
  assign oWidth_mWidth_prb_8 = and_550_cse;
  assign oWidth_mWidth_prb_9 = and_550_cse;
  assign or_dcpl_210 = or_dcpl_197;
endmodule
